* circuit generated from ALSIM
rrea n2_18380_8346 _X_n2_18380_8346 2.500000e-01
rr1cc n3_11630_7221 _X_n3_11630_7221 2.500000e-01
vb9 _X_n2_12755_4971 0 0
rr16 n2_16130_15096 _X_n2_16130_15096 2.500000e-01
rrec n2_17255_8346 _X_n2_17255_8346 2.500000e-01
vc1 _X_n2_15005_1596 0 0
rr1ce n3_13880_471 _X_n3_13880_471 2.500000e-01
rr100 n2_15005_10596 _X_n2_15005_10596 2.500000e-01
rr18 n2_20630_17346 _X_n2_20630_17346 2.500000e-01
rree n2_16130_8346 _X_n2_16130_8346 2.500000e-01
vc3 _X_n2_15005_2721 0 0
rr20 n2_19505_20721 _X_n2_19505_20721 2.500000e-01
rr102 n2_13880_10596 _X_n2_13880_10596 2.500000e-01
vc5 _X_n2_15005_3846 0 0
rr22 n2_17255_20721 _X_n2_17255_20721 2.500000e-01
rr104 n2_12755_10596 _X_n2_12755_10596 2.500000e-01
rr1da n3_20630_471 _X_n3_20630_471 2.500000e-01
vc7 _X_n2_15005_4971 0 0
rr24 n2_17255_19596 _X_n2_17255_19596 2.500000e-01
rr106 n2_11630_10596 _X_n2_11630_10596 2.500000e-01
rrfa n2_18380_10596 _X_n2_18380_10596 2.500000e-01
rr1dc n3_20630_2721 _X_n3_20630_2721 2.500000e-01
vc9 _X_n2_17255_471 0 0
rr26 n2_17255_18471 _X_n2_17255_18471 2.500000e-01
rr108 n2_1505_471 _X_n2_1505_471 2.500000e-01
rrfc n2_17255_10596 _X_n2_17255_10596 2.500000e-01
vd1 _X_n2_20630_1596 0 0
rr1de n3_18380_2721 _X_n3_18380_2721 2.500000e-01
rr110 n2_3755_3846 _X_n2_3755_3846 2.500000e-01
rr28 n2_17255_17346 _X_n2_17255_17346 2.500000e-01
rrfe n2_16130_10596 _X_n2_16130_10596 2.500000e-01
vd3 _X_n2_20630_3846 0 0
rr30 n2_15005_17346 _X_n2_15005_17346 2.500000e-01
rr112 n2_6005_471 _X_n2_6005_471 2.500000e-01
vd5 _X_n2_19505_3846 0 0
rr32 n2_15005_16221 _X_n2_15005_16221 2.500000e-01
rr114 n2_6005_1596 _X_n2_6005_1596 2.500000e-01
rr1ea n3_16130_7221 _X_n3_16130_7221 2.500000e-01
vd7 _X_n2_18380_3846 0 0
rr34 n2_15005_15096 _X_n2_15005_15096 2.500000e-01
rr116 n2_6005_2721 _X_n2_6005_2721 2.500000e-01
rr1ec n3_13880_7221 _X_n3_13880_7221 2.500000e-01
vd9 _X_n2_17255_3846 0 0
rr36 n2_12755_20721 _X_n2_12755_20721 2.500000e-01
rr118 n2_6005_3846 _X_n2_6005_3846 2.500000e-01
ve1 _X_n2_17255_6096 0 0
rr1ee n3_20630_9471 _X_n3_20630_9471 2.500000e-01
rr120 n2_8255_1596 _X_n2_8255_1596 2.500000e-01
rr38 n2_12755_19596 _X_n2_12755_19596 2.500000e-01
ve3 _X_n2_16130_6096 0 0
rr40 n2_12755_15096 _X_n2_12755_15096 2.500000e-01
rr122 n2_8255_2721 _X_n2_8255_2721 2.500000e-01
ve5 _X_n2_15005_6096 0 0
rr42 n2_12755_13971 _X_n2_12755_13971 2.500000e-01
rr124 n2_8255_3846 _X_n2_8255_3846 2.500000e-01
rr1fa n3_18380_11721 _X_n3_18380_11721 2.500000e-01
ve7 _X_n2_20630_8346 0 0
rr44 n2_12755_12846 _X_n2_12755_12846 2.500000e-01
rr126 n2_8255_4971 _X_n2_8255_4971 2.500000e-01
rr1fc n3_16130_11721 _X_n3_16130_11721 2.500000e-01
ve9 _X_n2_19505_8346 0 0
rr46 n2_10505_20721 _X_n2_10505_20721 2.500000e-01
rr128 n2_8255_6096 _X_n2_8255_6096 2.500000e-01
vf1 _X_n2_15005_8346 0 0
rr1fe n3_13880_11721 _X_n3_13880_11721 2.500000e-01
rr130 n2_10505_1596 _X_n2_10505_1596 2.500000e-01
rr48 n2_10505_19596 _X_n2_10505_19596 2.500000e-01
vf3 _X_n2_13880_8346 0 0
rr50 n2_10505_15096 _X_n2_10505_15096 2.500000e-01
rr132 n2_10505_2721 _X_n2_10505_2721 2.500000e-01
v1a1 _X_n3_7130_471 0 1.8
vf5 _X_n2_12755_8346 0 0
rr52 n2_10505_13971 _X_n2_10505_13971 2.500000e-01
vab _X_n2_7130_10596 0 0
rr134 n2_10505_3846 _X_n2_10505_3846 2.500000e-01
v1a3 _X_n3_7130_2721 0 1.8
vf7 _X_n2_20630_10596 0 0
rr54 n2_10505_12846 _X_n2_10505_12846 2.500000e-01
vad _X_n2_8255_10596 0 0
rr136 n2_10505_4971 _X_n2_10505_4971 2.500000e-01
v1a5 _X_n3_7130_4971 0 1.8
vf9 _X_n2_19505_10596 0 0
rr56 n2_10505_11721 _X_n2_10505_11721 2.500000e-01
vaf _X_n2_9380_10596 0 0
rr138 n2_10505_6096 _X_n2_10505_6096 2.500000e-01
v1a7 _X_n3_7130_7221 0 1.8
rr140 n2_10505_10596 _X_n2_10505_10596 2.500000e-01
rr58 n2_8255_20721 _X_n2_8255_20721 2.500000e-01
rr60 n2_8255_16221 _X_n2_8255_16221 2.500000e-01
v1a9 _X_n3_9380_471 0 1.8
rr142 n2_380_8346 _X_n2_380_8346 2.500000e-01
v1b1 _X_n3_9380_9471 0 1.8
vbb _X_n2_12755_6096 0 0
rr62 n2_8255_15096 _X_n2_8255_15096 2.500000e-01
rr144 n2_1505_8346 _X_n2_1505_8346 2.500000e-01
v1b3 _X_n3_380_9471 0 1.8
vbd _X_n2_12755_7221 0 0
rr1a n2_19505_17346 _X_n2_19505_17346 2.500000e-01
rr64 n2_8255_13971 _X_n2_8255_13971 2.500000e-01
rr146 n2_2630_8346 _X_n2_2630_8346 2.500000e-01
v1b5 _X_n3_2630_9471 0 1.8
vbf _X_n2_15005_471 0 0
rr1c n2_18380_17346 _X_n2_18380_17346 2.500000e-01
rr66 n2_6005_20721 _X_n2_6005_20721 2.500000e-01
rr148 n2_3755_8346 _X_n2_3755_8346 2.500000e-01
v1b7 _X_n3_4880_9471 0 1.8
rr150 n2_380_6096 _X_n2_380_6096 2.500000e-01
rr1e n2_20630_19596 _X_n2_20630_19596 2.500000e-01
rr68 n2_6005_19596 _X_n2_6005_19596 2.500000e-01
rr70 n2_3755_20721 _X_n2_3755_20721 2.500000e-01
v1b9 _X_n3_7130_9471 0 1.8
rr152 n2_1505_6096 _X_n2_1505_6096 2.500000e-01
rr0 n2_20630_12846 _X_n2_20630_12846 2.500000e-01
v1c1 _X_n3_380_4971 0 1.8
vcb _X_n2_17255_1596 0 0
rr72 n2_3755_19596 _X_n2_3755_19596 2.500000e-01
rr154 n2_2630_6096 _X_n2_2630_6096 2.500000e-01
rr10a n2_3755_471 _X_n2_3755_471 2.500000e-01
rr2 n2_19505_12846 _X_n2_19505_12846 2.500000e-01
v1c3 _X_n3_2630_4971 0 1.8
vcd _X_n2_17255_2721 0 0
rr2a n2_15005_20721 _X_n2_15005_20721 2.500000e-01
rr74 n2_3755_18471 _X_n2_3755_18471 2.500000e-01
rr156 n2_3755_6096 _X_n2_3755_6096 2.500000e-01
rr10c n2_3755_1596 _X_n2_3755_1596 2.500000e-01
rr4 n2_18380_12846 _X_n2_18380_12846 2.500000e-01
v1c5 _X_n3_380_2721 0 1.8
vcf _X_n2_19505_471 0 0
rr2c n2_15005_19596 _X_n2_15005_19596 2.500000e-01
rr76 n2_1505_20721 _X_n2_1505_20721 2.500000e-01
rr158 n2_4880_6096 _X_n2_4880_6096 2.500000e-01
rr10e n2_3755_2721 _X_n2_3755_2721 2.500000e-01
rr6 n2_17255_12846 _X_n2_17255_12846 2.500000e-01
v1c7 _X_n3_11630_471 0 1.8
rr160 n2_380_1596 _X_n2_380_1596 2.500000e-01
rr2e n2_15005_18471 _X_n2_15005_18471 2.500000e-01
rr78 n2_380_19596 _X_n2_380_19596 2.500000e-01
rr8 n2_16130_12846 _X_n2_16130_12846 2.500000e-01
rr80 n2_3755_17346 _X_n2_3755_17346 2.500000e-01
v1c9 _X_n3_11630_2721 0 1.8
rr162 n3_9380_20721 _X_n3_9380_20721 2.500000e-01
v1d1 _X_n3_13880_2721 0 1.8
vdb _X_n2_20630_6096 0 0
rr82 n2_380_15096 _X_n2_380_15096 2.500000e-01
rr164 n3_9380_18471 _X_n3_9380_18471 2.500000e-01
rr11a n2_6005_4971 _X_n2_6005_4971 2.500000e-01
v1d3 _X_n3_13880_4971 0 1.8
vdd _X_n2_19505_6096 0 0
rr3a n2_12755_18471 _X_n2_12755_18471 2.500000e-01
rr84 n2_1505_15096 _X_n2_1505_15096 2.500000e-01
rr166 n3_9380_16221 _X_n3_9380_16221 2.500000e-01
rr11c n2_6005_6096 _X_n2_6005_6096 2.500000e-01
v1d5 _X_n3_16130_471 0 1.8
vdf _X_n2_18380_6096 0 0
v11 _X_n2_19505_15096 0 0
rr3c n2_12755_17346 _X_n2_12755_17346 2.500000e-01
rr86 n2_2630_15096 _X_n2_2630_15096 2.500000e-01
rr168 n3_9380_13971 _X_n3_9380_13971 2.500000e-01
rr11e n2_8255_471 _X_n2_8255_471 2.500000e-01
v1d7 _X_n3_16130_2721 0 1.8
rr170 n3_4880_20721 _X_n3_4880_20721 2.500000e-01
v13 _X_n2_18380_15096 0 0
rr3e n2_12755_16221 _X_n2_12755_16221 2.500000e-01
rr88 n2_3755_15096 _X_n2_3755_15096 2.500000e-01
rr90 n2_1505_12846 _X_n2_1505_12846 2.500000e-01
v1d9 _X_n3_18380_471 0 1.8
rr172 n3_4880_18471 _X_n3_4880_18471 2.500000e-01
v15 _X_n2_17255_15096 0 0
v1e1 _X_n3_20630_4971 0 1.8
veb _X_n2_18380_8346 0 0
rr92 n2_2630_12846 _X_n2_2630_12846 2.500000e-01
rr174 n3_2630_20721 _X_n3_2630_20721 2.500000e-01
rr12a n2_8255_7221 _X_n2_8255_7221 2.500000e-01
v17 _X_n2_16130_15096 0 0
v1e3 _X_n3_18380_4971 0 1.8
ved _X_n2_17255_8346 0 0
rr4a n2_10505_18471 _X_n2_10505_18471 2.500000e-01
rr94 n2_3755_12846 _X_n2_3755_12846 2.500000e-01
rr176 n3_380_20721 _X_n3_380_20721 2.500000e-01
rr12c n2_8255_8346 _X_n2_8255_8346 2.500000e-01
v19 _X_n2_20630_17346 0 0
v1e5 _X_n3_16130_4971 0 1.8
vef _X_n2_16130_8346 0 0
v21 _X_n2_19505_20721 0 0
rr4c n2_10505_17346 _X_n2_10505_17346 2.500000e-01
rr96 n2_4880_12846 _X_n2_4880_12846 2.500000e-01
rr178 n3_380_18471 _X_n3_380_18471 2.500000e-01
rr12e n2_10505_471 _X_n2_10505_471 2.500000e-01
v1e7 _X_n3_20630_7221 0 1.8
rr180 n3_4880_16221 _X_n3_4880_16221 2.500000e-01
v23 _X_n2_17255_20721 0 0
rr4e n2_10505_16221 _X_n2_10505_16221 2.500000e-01
rr98 n2_6005_12846 _X_n2_6005_12846 2.500000e-01
v1e9 _X_n3_18380_7221 0 1.8
rr182 n3_380_13971 _X_n3_380_13971 2.500000e-01
v25 _X_n2_17255_19596 0 0
v1f1 _X_n3_18380_9471 0 1.8
vfb _X_n2_18380_10596 0 0
rr184 n3_2630_13971 _X_n3_2630_13971 2.500000e-01
rr13a n2_10505_7221 _X_n2_10505_7221 2.500000e-01
v27 _X_n2_17255_18471 0 0
v1f3 _X_n3_16130_9471 0 1.8
vfd _X_n2_17255_10596 0 0
rr5a n2_8255_19596 _X_n2_8255_19596 2.500000e-01
rr186 n3_4880_13971 _X_n3_4880_13971 2.500000e-01
rr13c n2_10505_8346 _X_n2_10505_8346 2.500000e-01
v29 _X_n2_17255_17346 0 0
v1f5 _X_n3_13880_9471 0 1.8
v1ab _X_n3_9380_2721 0 1.8
vff _X_n2_16130_10596 0 0
v31 _X_n2_15005_17346 0 0
rr5c n2_8255_18471 _X_n2_8255_18471 2.500000e-01
rr188 n3_7130_13971 _X_n3_7130_13971 2.500000e-01
rr13e n2_10505_9471 _X_n2_10505_9471 2.500000e-01
rr200 n3_20630_13971 _X_n3_20630_13971 2.500000e-01
v1f7 _X_n3_11630_9471 0 1.8
v1ad _X_n3_9380_4971 0 1.8
rr190 n3_7130_11721 _X_n3_7130_11721 2.500000e-01
* layer: M5,VDD net: 1
R554 n1_333_383 n1_521_383 1.342857e-01
R555 n1_521_383 n1_2400_383 1.342143e+00
R556 n1_2400_383 n1_2583_383 1.307143e-01
R557 n1_2583_383 n1_2771_383 1.342857e-01
R558 n1_2771_383 n1_2864_383 6.642857e-02
R559 n1_333_2543 n1_521_2543 1.342857e-01
R560 n1_521_2543 n1_2400_2543 1.342143e+00
R561 n1_2400_2543 n1_2583_2543 1.307143e-01
R562 n1_2583_2543 n1_2771_2543 1.342857e-01
R563 n1_2771_2543 n1_2864_2543 6.642857e-02
R564 n1_2864_2543 n1_4650_2543 1.275714e+00
R565 n1_4650_2543 n1_4833_2543 1.307143e-01
R566 n1_4833_2543 n1_5021_2543 1.342857e-01
R567 n1_5021_2543 n1_5114_2543 6.642857e-02
R568 n1_5114_2543 n1_6900_2543 1.275714e+00
R569 n1_6900_2543 n1_7083_2543 1.307143e-01
R570 n1_7083_2543 n1_7271_2543 1.342857e-01
R571 n1_7271_2543 n1_7364_2543 6.642857e-02
R572 n1_7364_2543 n1_9150_2543 1.275714e+00
R573 n1_9150_2543 n1_9333_2543 1.307143e-01
R574 n1_9333_2543 n1_9521_2543 1.342857e-01
R575 n1_9521_2543 n1_9614_2543 6.642857e-02
R576 n1_333_18527 n1_380_18527 3.357143e-02
R577 n1_380_18527 n1_521_18527 1.007143e-01
R578 n1_521_18527 n1_2400_18527 1.342143e+00
R579 n1_2400_18527 n1_2583_18527 1.307143e-01
R580 n1_2583_18527 n1_2630_18527 3.357143e-02
R581 n1_2630_18527 n1_2771_18527 1.007143e-01
R582 n1_2771_18527 n1_2864_18527 6.642857e-02
R583 n1_2864_18527 n1_4650_18527 1.275714e+00
R584 n1_4650_18527 n1_4833_18527 1.307143e-01
R585 n1_4833_18527 n1_4880_18527 3.357143e-02
R586 n1_4880_18527 n1_5021_18527 1.007143e-01
R587 n1_5021_18527 n1_5114_18527 6.642857e-02
R588 n1_5114_18527 n1_6900_18527 1.275714e+00
R589 n1_6900_18527 n1_7083_18527 1.307143e-01
R590 n1_7083_18527 n1_7130_18527 3.357143e-02
R591 n1_7130_18527 n1_7271_18527 1.007143e-01
R592 n1_7271_18527 n1_7364_18527 6.642857e-02
R593 n1_7364_18527 n1_9150_18527 1.275714e+00
R594 n1_9150_18527 n1_9333_18527 1.307143e-01
R595 n1_9333_18527 n1_9380_18527 3.357143e-02
R596 n1_9380_18527 n1_9521_18527 1.007143e-01
R597 n1_9521_18527 n1_9614_18527 6.642857e-02
R598 n1_333_20687 n1_380_20687 3.357143e-02
R599 n1_380_20687 n1_521_20687 1.007143e-01
R600 n1_521_20687 n1_2400_20687 1.342143e+00
R601 n1_2400_20687 n1_2583_20687 1.307143e-01
R602 n1_2583_20687 n1_2630_20687 3.357143e-02
R603 n1_2630_20687 n1_2771_20687 1.007143e-01
R604 n1_2771_20687 n1_2864_20687 6.642857e-02
R605 n1_2864_20687 n1_4650_20687 1.275714e+00
R606 n1_4650_20687 n1_4833_20687 1.307143e-01
R607 n1_4833_20687 n1_4880_20687 3.357143e-02
R608 n1_4880_20687 n1_5021_20687 1.007143e-01
R609 n1_5021_20687 n1_5114_20687 6.642857e-02
R610 n1_5114_20687 n1_6900_20687 1.275714e+00
R611 n1_6900_20687 n1_7083_20687 1.307143e-01
R612 n1_7083_20687 n1_7130_20687 3.357143e-02
R613 n1_7130_20687 n1_7271_20687 1.007143e-01
R614 n1_7271_20687 n1_7364_20687 6.642857e-02
R615 n1_7364_20687 n1_9150_20687 1.275714e+00
R616 n1_9150_20687 n1_9333_20687 1.307143e-01
R617 n1_9333_20687 n1_9380_20687 3.357143e-02
R618 n1_9380_20687 n1_9521_20687 1.007143e-01
R619 n1_9521_20687 n1_9614_20687 6.642857e-02
R620 n1_333_1079 n1_521_1079 1.074286e+00
R621 n1_521_1079 n1_2400_1079 1.073714e+01
R622 n1_2400_1079 n1_2583_1079 1.045714e+00
R623 n1_2583_1079 n1_2771_1079 1.074286e+00
R624 n1_2771_1079 n1_2864_1079 5.314286e-01
R625 n1_2864_1079 n1_4650_1079 1.020571e+01
R626 n1_4650_1079 n1_4833_1079 1.045714e+00
R627 n1_4833_1079 n1_5021_1079 1.074286e+00
R628 n1_5021_1079 n1_5114_1079 5.314286e-01
R629 n1_5114_1079 n1_6900_1079 1.020571e+01
R630 n1_6900_1079 n1_7083_1079 1.045714e+00
R631 n1_7083_1079 n1_7271_1079 1.074286e+00
R632 n1_7271_1079 n1_7364_1079 5.314286e-01
R633 n1_7364_1079 n1_9150_1079 1.020571e+01
R634 n1_9150_1079 n1_9333_1079 1.045714e+00
R635 n1_9333_1079 n1_9521_1079 1.074286e+00
R636 n1_9521_1079 n1_9614_1079 5.314286e-01
R637 n1_333_431 n1_380_431 2.685714e-01
R638 n1_380_431 n1_521_431 8.057143e-01
R639 n1_521_431 n1_2400_431 1.073714e+01
R640 n1_2400_431 n1_2583_431 1.045714e+00
R641 n1_2583_431 n1_2630_431 2.685714e-01
R642 n1_2630_431 n1_2771_431 8.057143e-01
R643 n1_2771_431 n1_2864_431 5.314286e-01
R644 n1_2864_431 n1_4650_431 1.020571e+01
R645 n1_4650_431 n1_4833_431 1.045714e+00
R646 n1_4833_431 n1_4880_431 2.685714e-01
R647 n1_4880_431 n1_5021_431 8.057143e-01
R648 n1_5021_431 n1_5114_431 5.314286e-01
R649 n1_5114_431 n1_6900_431 1.020571e+01
R650 n1_6900_431 n1_7083_431 1.045714e+00
R651 n1_7083_431 n1_7130_431 2.685714e-01
R652 n1_7130_431 n1_7271_431 8.057143e-01
R653 n1_7271_431 n1_7364_431 5.314286e-01
R654 n1_7364_431 n1_9150_431 1.020571e+01
R655 n1_9150_431 n1_9333_431 1.045714e+00
R656 n1_9333_431 n1_9380_431 2.685714e-01
R657 n1_9380_431 n1_9521_431 8.057143e-01
R658 n1_9521_431 n1_9614_431 5.314286e-01
R659 n1_333_464 n1_380_464 2.685714e-01
R660 n1_380_464 n1_2400_464 1.154286e+01
R661 n1_2400_464 n1_2583_464 1.045714e+00
R662 n1_2583_464 n1_2630_464 2.685714e-01
R663 n1_2630_464 n1_2864_464 1.337143e+00
R664 n1_2864_464 n1_4650_464 1.020571e+01
R665 n1_4650_464 n1_4833_464 1.045714e+00
R666 n1_4833_464 n1_4880_464 2.685714e-01
R667 n1_4880_464 n1_5114_464 1.337143e+00
R668 n1_5114_464 n1_6900_464 1.020571e+01
R669 n1_6900_464 n1_7083_464 1.045714e+00
R670 n1_7083_464 n1_7130_464 2.685714e-01
R671 n1_7130_464 n1_7364_464 1.337143e+00
R672 n1_7364_464 n1_9150_464 1.020571e+01
R673 n1_9150_464 n1_9333_464 1.045714e+00
R674 n1_9333_464 n1_9380_464 2.685714e-01
R675 n1_9380_464 n1_9614_464 1.337143e+00
R676 n1_333_647 n1_521_647 1.074286e+00
R677 n1_521_647 n1_2400_647 1.073714e+01
R678 n1_2400_647 n1_2583_647 1.045714e+00
R679 n1_2583_647 n1_2771_647 1.074286e+00
R680 n1_2771_647 n1_2864_647 5.314286e-01
R681 n1_2864_647 n1_4650_647 1.020571e+01
R682 n1_4650_647 n1_4833_647 1.045714e+00
R683 n1_4833_647 n1_5021_647 1.074286e+00
R684 n1_5021_647 n1_5114_647 5.314286e-01
R685 n1_5114_647 n1_6900_647 1.020571e+01
R686 n1_6900_647 n1_7083_647 1.045714e+00
R687 n1_7083_647 n1_7271_647 1.074286e+00
R688 n1_7271_647 n1_7364_647 5.314286e-01
R689 n1_7364_647 n1_9150_647 1.020571e+01
R690 n1_9150_647 n1_9333_647 1.045714e+00
R691 n1_9333_647 n1_9521_647 1.074286e+00
R692 n1_9521_647 n1_9614_647 5.314286e-01
R693 n1_333_680 n1_521_680 1.074286e+00
R694 n1_521_680 n1_2400_680 1.073714e+01
R695 n1_2400_680 n1_2583_680 1.045714e+00
R696 n1_2583_680 n1_2771_680 1.074286e+00
R697 n1_2771_680 n1_2864_680 5.314286e-01
R698 n1_2864_680 n1_4650_680 1.020571e+01
R699 n1_4650_680 n1_4833_680 1.045714e+00
R700 n1_4833_680 n1_5021_680 1.074286e+00
R701 n1_5021_680 n1_5114_680 5.314286e-01
R702 n1_5114_680 n1_6900_680 1.020571e+01
R703 n1_6900_680 n1_7083_680 1.045714e+00
R704 n1_7083_680 n1_7271_680 1.074286e+00
R705 n1_7271_680 n1_7364_680 5.314286e-01
R706 n1_7364_680 n1_9150_680 1.020571e+01
R707 n1_9150_680 n1_9333_680 1.045714e+00
R708 n1_9333_680 n1_9521_680 1.074286e+00
R709 n1_9521_680 n1_9614_680 5.314286e-01
R710 n1_333_863 n1_521_863 1.074286e+00
R711 n1_521_863 n1_2400_863 1.073714e+01
R712 n1_2400_863 n1_2583_863 1.045714e+00
R713 n1_2583_863 n1_2771_863 1.074286e+00
R714 n1_2771_863 n1_2864_863 5.314286e-01
R715 n1_2864_863 n1_4650_863 1.020571e+01
R716 n1_4650_863 n1_4833_863 1.045714e+00
R717 n1_4833_863 n1_5021_863 1.074286e+00
R718 n1_5021_863 n1_5114_863 5.314286e-01
R719 n1_5114_863 n1_6900_863 1.020571e+01
R720 n1_6900_863 n1_7083_863 1.045714e+00
R721 n1_7083_863 n1_7271_863 1.074286e+00
R722 n1_7271_863 n1_7364_863 5.314286e-01
R723 n1_7364_863 n1_9150_863 1.020571e+01
R724 n1_9150_863 n1_9333_863 1.045714e+00
R725 n1_9333_863 n1_9521_863 1.074286e+00
R726 n1_9521_863 n1_9614_863 5.314286e-01
R727 n1_333_896 n1_521_896 1.074286e+00
R728 n1_521_896 n1_2400_896 1.073714e+01
R729 n1_2400_896 n1_2583_896 1.045714e+00
R730 n1_2583_896 n1_2771_896 1.074286e+00
R731 n1_2771_896 n1_2864_896 5.314286e-01
R732 n1_2864_896 n1_4650_896 1.020571e+01
R733 n1_4650_896 n1_4833_896 1.045714e+00
R734 n1_4833_896 n1_5021_896 1.074286e+00
R735 n1_5021_896 n1_5114_896 5.314286e-01
R736 n1_5114_896 n1_6900_896 1.020571e+01
R737 n1_6900_896 n1_7083_896 1.045714e+00
R738 n1_7083_896 n1_7271_896 1.074286e+00
R739 n1_7271_896 n1_7364_896 5.314286e-01
R740 n1_7364_896 n1_9150_896 1.020571e+01
R741 n1_9150_896 n1_9333_896 1.045714e+00
R742 n1_9333_896 n1_9521_896 1.074286e+00
R743 n1_9521_896 n1_9614_896 5.314286e-01
R744 n1_333_9287 n1_521_9287 1.074286e+00
R745 n1_521_9287 n1_2583_9287 1.178286e+01
R746 n1_2583_9287 n1_2771_9287 1.074286e+00
R747 n1_2771_9287 n1_4833_9287 1.178286e+01
R748 n1_4833_9287 n1_5021_9287 1.074286e+00
R749 n1_5021_9287 n1_7083_9287 1.178286e+01
R750 n1_7083_9287 n1_7271_9287 1.074286e+00
R751 n1_7271_9287 n1_9333_9287 1.178286e+01
R752 n1_9333_9287 n1_9521_9287 1.074286e+00
R753 n1_11583_9287 n1_11771_9287 1.074286e+00
R754 n1_11771_9287 n1_13833_9287 1.178286e+01
R755 n1_13833_9287 n1_14021_9287 1.074286e+00
R756 n1_14021_9287 n1_16083_9287 1.178286e+01
R757 n1_16083_9287 n1_16271_9287 1.074286e+00
R758 n1_16271_9287 n1_18333_9287 1.178286e+01
R759 n1_18333_9287 n1_18521_9287 1.074286e+00
R760 n1_18521_9287 n1_20583_9287 1.178286e+01
R761 n1_20583_9287 n1_20771_9287 1.074286e+00
R762 n1_333_9320 n1_521_9320 1.074286e+00
R763 n1_521_9320 n1_2583_9320 1.178286e+01
R764 n1_2583_9320 n1_2771_9320 1.074286e+00
R765 n1_2771_9320 n1_4833_9320 1.178286e+01
R766 n1_4833_9320 n1_5021_9320 1.074286e+00
R767 n1_5021_9320 n1_7083_9320 1.178286e+01
R768 n1_7083_9320 n1_7271_9320 1.074286e+00
R769 n1_7271_9320 n1_9333_9320 1.178286e+01
R770 n1_9333_9320 n1_9521_9320 1.074286e+00
R771 n1_11583_9320 n1_11771_9320 1.074286e+00
R772 n1_11771_9320 n1_13833_9320 1.178286e+01
R773 n1_13833_9320 n1_14021_9320 1.074286e+00
R774 n1_14021_9320 n1_16083_9320 1.178286e+01
R775 n1_16083_9320 n1_16271_9320 1.074286e+00
R776 n1_16271_9320 n1_18333_9320 1.178286e+01
R777 n1_18333_9320 n1_18521_9320 1.074286e+00
R778 n1_18521_9320 n1_20583_9320 1.178286e+01
R779 n1_20583_9320 n1_20771_9320 1.074286e+00
R780 n1_333_9503 n1_380_9503 2.685714e-01
R781 n1_380_9503 n1_521_9503 8.057143e-01
R782 n1_521_9503 n1_2583_9503 1.178286e+01
R783 n1_2583_9503 n1_2630_9503 2.685714e-01
R784 n1_2630_9503 n1_2771_9503 8.057143e-01
R785 n1_2771_9503 n1_4833_9503 1.178286e+01
R786 n1_4833_9503 n1_4880_9503 2.685714e-01
R787 n1_4880_9503 n1_5021_9503 8.057143e-01
R788 n1_5021_9503 n1_7083_9503 1.178286e+01
R789 n1_7083_9503 n1_7130_9503 2.685714e-01
R790 n1_7130_9503 n1_7271_9503 8.057143e-01
R791 n1_7271_9503 n1_9333_9503 1.178286e+01
R792 n1_9333_9503 n1_9380_9503 2.685714e-01
R793 n1_9380_9503 n1_9521_9503 8.057143e-01
R794 n1_11583_9503 n1_11630_9503 2.685714e-01
R795 n1_11630_9503 n1_11771_9503 8.057143e-01
R796 n1_11771_9503 n1_13833_9503 1.178286e+01
R797 n1_13833_9503 n1_13880_9503 2.685714e-01
R798 n1_13880_9503 n1_14021_9503 8.057143e-01
R799 n1_14021_9503 n1_16083_9503 1.178286e+01
R800 n1_16083_9503 n1_16130_9503 2.685714e-01
R801 n1_16130_9503 n1_16271_9503 8.057143e-01
R802 n1_16271_9503 n1_18333_9503 1.178286e+01
R803 n1_18333_9503 n1_18380_9503 2.685714e-01
R804 n1_18380_9503 n1_18521_9503 8.057143e-01
R805 n1_18521_9503 n1_20583_9503 1.178286e+01
R806 n1_20583_9503 n1_20630_9503 2.685714e-01
R807 n1_20630_9503 n1_20771_9503 8.057143e-01
R808 n1_333_9536 n1_380_9536 2.685714e-01
R809 n1_380_9536 n1_521_9536 8.057143e-01
R810 n1_521_9536 n1_2583_9536 1.178286e+01
R811 n1_2583_9536 n1_2630_9536 2.685714e-01
R812 n1_2630_9536 n1_2771_9536 8.057143e-01
R813 n1_2771_9536 n1_4833_9536 1.178286e+01
R814 n1_4833_9536 n1_4880_9536 2.685714e-01
R815 n1_4880_9536 n1_5021_9536 8.057143e-01
R816 n1_5021_9536 n1_7083_9536 1.178286e+01
R817 n1_7083_9536 n1_7130_9536 2.685714e-01
R818 n1_7130_9536 n1_7271_9536 8.057143e-01
R819 n1_7271_9536 n1_9333_9536 1.178286e+01
R820 n1_9333_9536 n1_9380_9536 2.685714e-01
R821 n1_9380_9536 n1_9521_9536 8.057143e-01
R822 n1_11583_9536 n1_11630_9536 2.685714e-01
R823 n1_11630_9536 n1_11771_9536 8.057143e-01
R824 n1_11771_9536 n1_13833_9536 1.178286e+01
R825 n1_13833_9536 n1_13880_9536 2.685714e-01
R826 n1_13880_9536 n1_14021_9536 8.057143e-01
R827 n1_14021_9536 n1_16083_9536 1.178286e+01
R828 n1_16083_9536 n1_16130_9536 2.685714e-01
R829 n1_16130_9536 n1_16271_9536 8.057143e-01
R830 n1_16271_9536 n1_18333_9536 1.178286e+01
R831 n1_18333_9536 n1_18380_9536 2.685714e-01
R832 n1_18380_9536 n1_18521_9536 8.057143e-01
R833 n1_18521_9536 n1_20583_9536 1.178286e+01
R834 n1_20583_9536 n1_20630_9536 2.685714e-01
R835 n1_20630_9536 n1_20771_9536 8.057143e-01
R836 n1_333_9719 n1_521_9719 1.074286e+00
R837 n1_521_9719 n1_2583_9719 1.178286e+01
R838 n1_2583_9719 n1_2771_9719 1.074286e+00
R839 n1_2771_9719 n1_4833_9719 1.178286e+01
R840 n1_4833_9719 n1_5021_9719 1.074286e+00
R841 n1_5021_9719 n1_7083_9719 1.178286e+01
R842 n1_7083_9719 n1_7271_9719 1.074286e+00
R843 n1_7271_9719 n1_9333_9719 1.178286e+01
R844 n1_9333_9719 n1_9521_9719 1.074286e+00
R845 n1_11583_9719 n1_11771_9719 1.074286e+00
R846 n1_11771_9719 n1_13833_9719 1.178286e+01
R847 n1_13833_9719 n1_14021_9719 1.074286e+00
R848 n1_14021_9719 n1_16083_9719 1.178286e+01
R849 n1_16083_9719 n1_16271_9719 1.074286e+00
R850 n1_16271_9719 n1_18333_9719 1.178286e+01
R851 n1_18333_9719 n1_18521_9719 1.074286e+00
R852 n1_18521_9719 n1_20583_9719 1.178286e+01
R853 n1_20583_9719 n1_20771_9719 1.074286e+00
R854 n1_333_9752 n1_521_9752 1.074286e+00
R855 n1_521_9752 n1_2583_9752 1.178286e+01
R856 n1_2583_9752 n1_2771_9752 1.074286e+00
R857 n1_2771_9752 n1_4833_9752 1.178286e+01
R858 n1_4833_9752 n1_5021_9752 1.074286e+00
R859 n1_5021_9752 n1_7083_9752 1.178286e+01
R860 n1_7083_9752 n1_7271_9752 1.074286e+00
R861 n1_7271_9752 n1_9333_9752 1.178286e+01
R862 n1_9333_9752 n1_9521_9752 1.074286e+00
R863 n1_11583_9752 n1_11771_9752 1.074286e+00
R864 n1_11771_9752 n1_13833_9752 1.178286e+01
R865 n1_13833_9752 n1_14021_9752 1.074286e+00
R866 n1_14021_9752 n1_16083_9752 1.178286e+01
R867 n1_16083_9752 n1_16271_9752 1.074286e+00
R868 n1_16271_9752 n1_18333_9752 1.178286e+01
R869 n1_18333_9752 n1_18521_9752 1.074286e+00
R870 n1_18521_9752 n1_20583_9752 1.178286e+01
R871 n1_20583_9752 n1_20771_9752 1.074286e+00
R872 n1_333_9935 n1_521_9935 1.074286e+00
R873 n1_521_9935 n1_2583_9935 1.178286e+01
R874 n1_2583_9935 n1_2771_9935 1.074286e+00
R875 n1_2771_9935 n1_4833_9935 1.178286e+01
R876 n1_4833_9935 n1_5021_9935 1.074286e+00
R877 n1_5021_9935 n1_7083_9935 1.178286e+01
R878 n1_7083_9935 n1_7271_9935 1.074286e+00
R879 n1_7271_9935 n1_9333_9935 1.178286e+01
R880 n1_9333_9935 n1_9521_9935 1.074286e+00
R881 n1_11583_9935 n1_11771_9935 1.074286e+00
R882 n1_11771_9935 n1_13833_9935 1.178286e+01
R883 n1_13833_9935 n1_14021_9935 1.074286e+00
R884 n1_14021_9935 n1_16083_9935 1.178286e+01
R885 n1_16083_9935 n1_16271_9935 1.074286e+00
R886 n1_16271_9935 n1_18333_9935 1.178286e+01
R887 n1_18333_9935 n1_18521_9935 1.074286e+00
R888 n1_18521_9935 n1_20583_9935 1.178286e+01
R889 n1_20583_9935 n1_20771_9935 1.074286e+00
R890 n1_333_9968 n1_521_9968 1.074286e+00
R891 n1_521_9968 n1_2583_9968 1.178286e+01
R892 n1_2583_9968 n1_2771_9968 1.074286e+00
R893 n1_2771_9968 n1_4833_9968 1.178286e+01
R894 n1_4833_9968 n1_5021_9968 1.074286e+00
R895 n1_5021_9968 n1_7083_9968 1.178286e+01
R896 n1_7083_9968 n1_7271_9968 1.074286e+00
R897 n1_7271_9968 n1_9333_9968 1.178286e+01
R898 n1_9333_9968 n1_9521_9968 1.074286e+00
R899 n1_11583_9968 n1_11771_9968 1.074286e+00
R900 n1_11771_9968 n1_13833_9968 1.178286e+01
R901 n1_13833_9968 n1_14021_9968 1.074286e+00
R902 n1_14021_9968 n1_16083_9968 1.178286e+01
R903 n1_16083_9968 n1_16271_9968 1.074286e+00
R904 n1_16271_9968 n1_18333_9968 1.178286e+01
R905 n1_18333_9968 n1_18521_9968 1.074286e+00
R906 n1_18521_9968 n1_20583_9968 1.178286e+01
R907 n1_20583_9968 n1_20771_9968 1.074286e+00
R908 n1_333_10151 n1_521_10151 1.074286e+00
R909 n1_521_10151 n1_2583_10151 1.178286e+01
R910 n1_2583_10151 n1_2771_10151 1.074286e+00
R911 n1_2771_10151 n1_4833_10151 1.178286e+01
R912 n1_4833_10151 n1_5021_10151 1.074286e+00
R913 n1_5021_10151 n1_7083_10151 1.178286e+01
R914 n1_7083_10151 n1_7271_10151 1.074286e+00
R915 n1_7271_10151 n1_9333_10151 1.178286e+01
R916 n1_9333_10151 n1_9521_10151 1.074286e+00
R917 n1_11583_10151 n1_11771_10151 1.074286e+00
R918 n1_11771_10151 n1_13833_10151 1.178286e+01
R919 n1_13833_10151 n1_14021_10151 1.074286e+00
R920 n1_14021_10151 n1_16083_10151 1.178286e+01
R921 n1_16083_10151 n1_16271_10151 1.074286e+00
R922 n1_16271_10151 n1_18333_10151 1.178286e+01
R923 n1_18333_10151 n1_18521_10151 1.074286e+00
R924 n1_18521_10151 n1_20583_10151 1.178286e+01
R925 n1_20583_10151 n1_20771_10151 1.074286e+00
R926 n1_333_10184 n1_521_10184 1.074286e+00
R927 n1_521_10184 n1_2583_10184 1.178286e+01
R928 n1_2583_10184 n1_2771_10184 1.074286e+00
R929 n1_2771_10184 n1_4833_10184 1.178286e+01
R930 n1_4833_10184 n1_5021_10184 1.074286e+00
R931 n1_5021_10184 n1_7083_10184 1.178286e+01
R932 n1_7083_10184 n1_7271_10184 1.074286e+00
R933 n1_7271_10184 n1_9333_10184 1.178286e+01
R934 n1_9333_10184 n1_9521_10184 1.074286e+00
R935 n1_11583_10184 n1_11771_10184 1.074286e+00
R936 n1_11771_10184 n1_13833_10184 1.178286e+01
R937 n1_13833_10184 n1_14021_10184 1.074286e+00
R938 n1_14021_10184 n1_16083_10184 1.178286e+01
R939 n1_16083_10184 n1_16271_10184 1.074286e+00
R940 n1_16271_10184 n1_18333_10184 1.178286e+01
R941 n1_18333_10184 n1_18521_10184 1.074286e+00
R942 n1_18521_10184 n1_20583_10184 1.178286e+01
R943 n1_20583_10184 n1_20771_10184 1.074286e+00
R944 n1_333_10367 n1_521_10367 1.074286e+00
R945 n1_521_10367 n1_2583_10367 1.178286e+01
R946 n1_2583_10367 n1_2771_10367 1.074286e+00
R947 n1_2771_10367 n1_4833_10367 1.178286e+01
R948 n1_4833_10367 n1_5021_10367 1.074286e+00
R949 n1_5021_10367 n1_7083_10367 1.178286e+01
R950 n1_7083_10367 n1_7271_10367 1.074286e+00
R951 n1_7271_10367 n1_9333_10367 1.178286e+01
R952 n1_9333_10367 n1_9521_10367 1.074286e+00
R953 n1_11583_10367 n1_11771_10367 1.074286e+00
R954 n1_11771_10367 n1_13833_10367 1.178286e+01
R955 n1_13833_10367 n1_14021_10367 1.074286e+00
R956 n1_14021_10367 n1_16083_10367 1.178286e+01
R957 n1_16083_10367 n1_16271_10367 1.074286e+00
R958 n1_16271_10367 n1_18333_10367 1.178286e+01
R959 n1_18333_10367 n1_18521_10367 1.074286e+00
R960 n1_18521_10367 n1_20583_10367 1.178286e+01
R961 n1_20583_10367 n1_20771_10367 1.074286e+00
R962 n1_333_10400 n1_521_10400 1.074286e+00
R963 n1_521_10400 n1_2583_10400 1.178286e+01
R964 n1_2583_10400 n1_2771_10400 1.074286e+00
R965 n1_2771_10400 n1_4833_10400 1.178286e+01
R966 n1_4833_10400 n1_5021_10400 1.074286e+00
R967 n1_5021_10400 n1_7083_10400 1.178286e+01
R968 n1_7083_10400 n1_7271_10400 1.074286e+00
R969 n1_7271_10400 n1_9333_10400 1.178286e+01
R970 n1_9333_10400 n1_9521_10400 1.074286e+00
R971 n1_11583_10400 n1_11771_10400 1.074286e+00
R972 n1_11771_10400 n1_13833_10400 1.178286e+01
R973 n1_13833_10400 n1_14021_10400 1.074286e+00
R974 n1_14021_10400 n1_16083_10400 1.178286e+01
R975 n1_16083_10400 n1_16271_10400 1.074286e+00
R976 n1_16271_10400 n1_18333_10400 1.178286e+01
R977 n1_18333_10400 n1_18521_10400 1.074286e+00
R978 n1_18521_10400 n1_20583_10400 1.178286e+01
R979 n1_20583_10400 n1_20771_10400 1.074286e+00
R980 n1_521_10616 n1_2771_10616 1.285714e+01
R981 n1_2771_10616 n1_5021_10616 1.285714e+01
R982 n1_5021_10616 n1_7271_10616 1.285714e+01
R983 n1_7271_10616 n1_9521_10616 1.285714e+01
R984 n1_11771_10616 n1_14021_10616 1.285714e+01
R985 n1_14021_10616 n1_16271_10616 1.285714e+01
R986 n1_16271_10616 n1_18521_10616 1.285714e+01
R987 n1_18521_10616 n1_20771_10616 1.285714e+01
R988 n1_333_10799 n1_521_10799 1.074286e+00
R989 n1_521_10799 n1_2583_10799 1.178286e+01
R990 n1_2583_10799 n1_2771_10799 1.074286e+00
R991 n1_2771_10799 n1_4833_10799 1.178286e+01
R992 n1_4833_10799 n1_5021_10799 1.074286e+00
R993 n1_5021_10799 n1_7083_10799 1.178286e+01
R994 n1_7083_10799 n1_7271_10799 1.074286e+00
R995 n1_7271_10799 n1_9333_10799 1.178286e+01
R996 n1_9333_10799 n1_9521_10799 1.074286e+00
R997 n1_11583_10799 n1_11771_10799 1.074286e+00
R998 n1_11771_10799 n1_13833_10799 1.178286e+01
R999 n1_13833_10799 n1_14021_10799 1.074286e+00
R1000 n1_14021_10799 n1_16083_10799 1.178286e+01
R1001 n1_16083_10799 n1_16271_10799 1.074286e+00
R1002 n1_16271_10799 n1_18333_10799 1.178286e+01
R1003 n1_18333_10799 n1_18521_10799 1.074286e+00
R1004 n1_18521_10799 n1_20583_10799 1.178286e+01
R1005 n1_20583_10799 n1_20771_10799 1.074286e+00
R1006 n1_333_10832 n1_521_10832 1.074286e+00
R1007 n1_521_10832 n1_2583_10832 1.178286e+01
R1008 n1_2583_10832 n1_2771_10832 1.074286e+00
R1009 n1_2771_10832 n1_4833_10832 1.178286e+01
R1010 n1_4833_10832 n1_5021_10832 1.074286e+00
R1011 n1_5021_10832 n1_7083_10832 1.178286e+01
R1012 n1_7083_10832 n1_7271_10832 1.074286e+00
R1013 n1_7271_10832 n1_9333_10832 1.178286e+01
R1014 n1_9333_10832 n1_9521_10832 1.074286e+00
R1015 n1_11583_10832 n1_11771_10832 1.074286e+00
R1016 n1_11771_10832 n1_13833_10832 1.178286e+01
R1017 n1_13833_10832 n1_14021_10832 1.074286e+00
R1018 n1_14021_10832 n1_16083_10832 1.178286e+01
R1019 n1_16083_10832 n1_16271_10832 1.074286e+00
R1020 n1_16271_10832 n1_18333_10832 1.178286e+01
R1021 n1_18333_10832 n1_18521_10832 1.074286e+00
R1022 n1_18521_10832 n1_20583_10832 1.178286e+01
R1023 n1_20583_10832 n1_20771_10832 1.074286e+00
R1024 n1_333_11015 n1_521_11015 1.074286e+00
R1025 n1_521_11015 n1_2583_11015 1.178286e+01
R1026 n1_2583_11015 n1_2771_11015 1.074286e+00
R1027 n1_2771_11015 n1_4833_11015 1.178286e+01
R1028 n1_4833_11015 n1_5021_11015 1.074286e+00
R1029 n1_5021_11015 n1_7083_11015 1.178286e+01
R1030 n1_7083_11015 n1_7271_11015 1.074286e+00
R1031 n1_7271_11015 n1_9333_11015 1.178286e+01
R1032 n1_9333_11015 n1_9521_11015 1.074286e+00
R1033 n1_11583_11015 n1_11771_11015 1.074286e+00
R1034 n1_11771_11015 n1_13833_11015 1.178286e+01
R1035 n1_13833_11015 n1_14021_11015 1.074286e+00
R1036 n1_14021_11015 n1_16083_11015 1.178286e+01
R1037 n1_16083_11015 n1_16271_11015 1.074286e+00
R1038 n1_16271_11015 n1_18333_11015 1.178286e+01
R1039 n1_18333_11015 n1_18521_11015 1.074286e+00
R1040 n1_18521_11015 n1_20583_11015 1.178286e+01
R1041 n1_20583_11015 n1_20771_11015 1.074286e+00
R1042 n1_333_11048 n1_521_11048 1.074286e+00
R1043 n1_521_11048 n1_2583_11048 1.178286e+01
R1044 n1_2583_11048 n1_2771_11048 1.074286e+00
R1045 n1_2771_11048 n1_4833_11048 1.178286e+01
R1046 n1_4833_11048 n1_5021_11048 1.074286e+00
R1047 n1_5021_11048 n1_7083_11048 1.178286e+01
R1048 n1_7083_11048 n1_7271_11048 1.074286e+00
R1049 n1_7271_11048 n1_9333_11048 1.178286e+01
R1050 n1_9333_11048 n1_9521_11048 1.074286e+00
R1051 n1_11583_11048 n1_11771_11048 1.074286e+00
R1052 n1_11771_11048 n1_13833_11048 1.178286e+01
R1053 n1_13833_11048 n1_14021_11048 1.074286e+00
R1054 n1_14021_11048 n1_16083_11048 1.178286e+01
R1055 n1_16083_11048 n1_16271_11048 1.074286e+00
R1056 n1_16271_11048 n1_18333_11048 1.178286e+01
R1057 n1_18333_11048 n1_18521_11048 1.074286e+00
R1058 n1_18521_11048 n1_20583_11048 1.178286e+01
R1059 n1_20583_11048 n1_20771_11048 1.074286e+00
R1060 n1_333_11231 n1_521_11231 1.074286e+00
R1061 n1_521_11231 n1_2583_11231 1.178286e+01
R1062 n1_2583_11231 n1_2771_11231 1.074286e+00
R1063 n1_2771_11231 n1_4833_11231 1.178286e+01
R1064 n1_4833_11231 n1_5021_11231 1.074286e+00
R1065 n1_5021_11231 n1_7083_11231 1.178286e+01
R1066 n1_7083_11231 n1_7271_11231 1.074286e+00
R1067 n1_7271_11231 n1_9333_11231 1.178286e+01
R1068 n1_9333_11231 n1_9521_11231 1.074286e+00
R1069 n1_11583_11231 n1_11771_11231 1.074286e+00
R1070 n1_11771_11231 n1_13833_11231 1.178286e+01
R1071 n1_13833_11231 n1_14021_11231 1.074286e+00
R1072 n1_14021_11231 n1_16083_11231 1.178286e+01
R1073 n1_16083_11231 n1_16271_11231 1.074286e+00
R1074 n1_16271_11231 n1_18333_11231 1.178286e+01
R1075 n1_18333_11231 n1_18521_11231 1.074286e+00
R1076 n1_18521_11231 n1_20583_11231 1.178286e+01
R1077 n1_20583_11231 n1_20771_11231 1.074286e+00
R1078 n1_333_11264 n1_521_11264 1.074286e+00
R1079 n1_521_11264 n1_2583_11264 1.178286e+01
R1080 n1_2583_11264 n1_2771_11264 1.074286e+00
R1081 n1_2771_11264 n1_4833_11264 1.178286e+01
R1082 n1_4833_11264 n1_5021_11264 1.074286e+00
R1083 n1_5021_11264 n1_7083_11264 1.178286e+01
R1084 n1_7083_11264 n1_7271_11264 1.074286e+00
R1085 n1_7271_11264 n1_9333_11264 1.178286e+01
R1086 n1_9333_11264 n1_9521_11264 1.074286e+00
R1087 n1_11583_11264 n1_11771_11264 1.074286e+00
R1088 n1_11771_11264 n1_13833_11264 1.178286e+01
R1089 n1_13833_11264 n1_14021_11264 1.074286e+00
R1090 n1_14021_11264 n1_16083_11264 1.178286e+01
R1091 n1_16083_11264 n1_16271_11264 1.074286e+00
R1092 n1_16271_11264 n1_18333_11264 1.178286e+01
R1093 n1_18333_11264 n1_18521_11264 1.074286e+00
R1094 n1_18521_11264 n1_20583_11264 1.178286e+01
R1095 n1_20583_11264 n1_20771_11264 1.074286e+00
R1096 n1_333_11447 n1_521_11447 1.074286e+00
R1097 n1_521_11447 n1_2583_11447 1.178286e+01
R1098 n1_2583_11447 n1_2771_11447 1.074286e+00
R1099 n1_2771_11447 n1_4833_11447 1.178286e+01
R1100 n1_4833_11447 n1_5021_11447 1.074286e+00
R1101 n1_5021_11447 n1_7083_11447 1.178286e+01
R1102 n1_7083_11447 n1_7271_11447 1.074286e+00
R1103 n1_7271_11447 n1_9333_11447 1.178286e+01
R1104 n1_9333_11447 n1_9521_11447 1.074286e+00
R1105 n1_11583_11447 n1_11771_11447 1.074286e+00
R1106 n1_11771_11447 n1_13833_11447 1.178286e+01
R1107 n1_13833_11447 n1_14021_11447 1.074286e+00
R1108 n1_14021_11447 n1_16083_11447 1.178286e+01
R1109 n1_16083_11447 n1_16271_11447 1.074286e+00
R1110 n1_16271_11447 n1_18333_11447 1.178286e+01
R1111 n1_18333_11447 n1_18521_11447 1.074286e+00
R1112 n1_18521_11447 n1_20583_11447 1.178286e+01
R1113 n1_20583_11447 n1_20771_11447 1.074286e+00
R1114 n1_333_11480 n1_521_11480 1.074286e+00
R1115 n1_521_11480 n1_2583_11480 1.178286e+01
R1116 n1_2583_11480 n1_2771_11480 1.074286e+00
R1117 n1_2771_11480 n1_4833_11480 1.178286e+01
R1118 n1_4833_11480 n1_5021_11480 1.074286e+00
R1119 n1_5021_11480 n1_7083_11480 1.178286e+01
R1120 n1_7083_11480 n1_7271_11480 1.074286e+00
R1121 n1_7271_11480 n1_9333_11480 1.178286e+01
R1122 n1_9333_11480 n1_9521_11480 1.074286e+00
R1123 n1_11583_11480 n1_11771_11480 1.074286e+00
R1124 n1_11771_11480 n1_13833_11480 1.178286e+01
R1125 n1_13833_11480 n1_14021_11480 1.074286e+00
R1126 n1_14021_11480 n1_16083_11480 1.178286e+01
R1127 n1_16083_11480 n1_16271_11480 1.074286e+00
R1128 n1_16271_11480 n1_18333_11480 1.178286e+01
R1129 n1_18333_11480 n1_18521_11480 1.074286e+00
R1130 n1_18521_11480 n1_20583_11480 1.178286e+01
R1131 n1_20583_11480 n1_20771_11480 1.074286e+00
R1132 n1_333_11663 n1_380_11663 2.685714e-01
R1133 n1_380_11663 n1_521_11663 8.057143e-01
R1134 n1_521_11663 n1_2583_11663 1.178286e+01
R1135 n1_2583_11663 n1_2630_11663 2.685714e-01
R1136 n1_2630_11663 n1_2771_11663 8.057143e-01
R1137 n1_2771_11663 n1_4833_11663 1.178286e+01
R1138 n1_4833_11663 n1_4880_11663 2.685714e-01
R1139 n1_4880_11663 n1_5021_11663 8.057143e-01
R1140 n1_5021_11663 n1_7083_11663 1.178286e+01
R1141 n1_7083_11663 n1_7130_11663 2.685714e-01
R1142 n1_7130_11663 n1_7271_11663 8.057143e-01
R1143 n1_7271_11663 n1_9333_11663 1.178286e+01
R1144 n1_9333_11663 n1_9380_11663 2.685714e-01
R1145 n1_9380_11663 n1_9521_11663 8.057143e-01
R1146 n1_11583_11663 n1_11630_11663 2.685714e-01
R1147 n1_11630_11663 n1_11771_11663 8.057143e-01
R1148 n1_11771_11663 n1_13833_11663 1.178286e+01
R1149 n1_13833_11663 n1_13880_11663 2.685714e-01
R1150 n1_13880_11663 n1_14021_11663 8.057143e-01
R1151 n1_14021_11663 n1_16083_11663 1.178286e+01
R1152 n1_16083_11663 n1_16130_11663 2.685714e-01
R1153 n1_16130_11663 n1_16271_11663 8.057143e-01
R1154 n1_16271_11663 n1_18333_11663 1.178286e+01
R1155 n1_18333_11663 n1_18380_11663 2.685714e-01
R1156 n1_18380_11663 n1_18521_11663 8.057143e-01
R1157 n1_18521_11663 n1_20583_11663 1.178286e+01
R1158 n1_20583_11663 n1_20630_11663 2.685714e-01
R1159 n1_20630_11663 n1_20771_11663 8.057143e-01
R1160 n1_333_11696 n1_380_11696 2.685714e-01
R1161 n1_380_11696 n1_521_11696 8.057143e-01
R1162 n1_521_11696 n1_2583_11696 1.178286e+01
R1163 n1_2583_11696 n1_2630_11696 2.685714e-01
R1164 n1_2630_11696 n1_2771_11696 8.057143e-01
R1165 n1_2771_11696 n1_4833_11696 1.178286e+01
R1166 n1_4833_11696 n1_4880_11696 2.685714e-01
R1167 n1_4880_11696 n1_5021_11696 8.057143e-01
R1168 n1_5021_11696 n1_7083_11696 1.178286e+01
R1169 n1_7083_11696 n1_7130_11696 2.685714e-01
R1170 n1_7130_11696 n1_7271_11696 8.057143e-01
R1171 n1_7271_11696 n1_9333_11696 1.178286e+01
R1172 n1_9333_11696 n1_9380_11696 2.685714e-01
R1173 n1_9380_11696 n1_9521_11696 8.057143e-01
R1174 n1_11583_11696 n1_11630_11696 2.685714e-01
R1175 n1_11630_11696 n1_11771_11696 8.057143e-01
R1176 n1_11771_11696 n1_13833_11696 1.178286e+01
R1177 n1_13833_11696 n1_13880_11696 2.685714e-01
R1178 n1_13880_11696 n1_14021_11696 8.057143e-01
R1179 n1_14021_11696 n1_16083_11696 1.178286e+01
R1180 n1_16083_11696 n1_16130_11696 2.685714e-01
R1181 n1_16130_11696 n1_16271_11696 8.057143e-01
R1182 n1_16271_11696 n1_18333_11696 1.178286e+01
R1183 n1_18333_11696 n1_18380_11696 2.685714e-01
R1184 n1_18380_11696 n1_18521_11696 8.057143e-01
R1185 n1_18521_11696 n1_20583_11696 1.178286e+01
R1186 n1_20583_11696 n1_20630_11696 2.685714e-01
R1187 n1_20630_11696 n1_20771_11696 8.057143e-01
R1188 n1_333_11879 n1_521_11879 1.074286e+00
R1189 n1_521_11879 n1_2583_11879 1.178286e+01
R1190 n1_2583_11879 n1_2771_11879 1.074286e+00
R1191 n1_2771_11879 n1_4833_11879 1.178286e+01
R1192 n1_4833_11879 n1_5021_11879 1.074286e+00
R1193 n1_5021_11879 n1_7083_11879 1.178286e+01
R1194 n1_7083_11879 n1_7271_11879 1.074286e+00
R1195 n1_7271_11879 n1_9333_11879 1.178286e+01
R1196 n1_9333_11879 n1_9521_11879 1.074286e+00
R1197 n1_11583_11879 n1_11771_11879 1.074286e+00
R1198 n1_11771_11879 n1_13833_11879 1.178286e+01
R1199 n1_13833_11879 n1_14021_11879 1.074286e+00
R1200 n1_14021_11879 n1_16083_11879 1.178286e+01
R1201 n1_16083_11879 n1_16271_11879 1.074286e+00
R1202 n1_16271_11879 n1_18333_11879 1.178286e+01
R1203 n1_18333_11879 n1_18521_11879 1.074286e+00
R1204 n1_18521_11879 n1_20583_11879 1.178286e+01
R1205 n1_20583_11879 n1_20771_11879 1.074286e+00
R1206 n1_333_11912 n1_521_11912 1.074286e+00
R1207 n1_521_11912 n1_2583_11912 1.178286e+01
R1208 n1_2583_11912 n1_2771_11912 1.074286e+00
R1209 n1_2771_11912 n1_4833_11912 1.178286e+01
R1210 n1_4833_11912 n1_5021_11912 1.074286e+00
R1211 n1_5021_11912 n1_7083_11912 1.178286e+01
R1212 n1_7083_11912 n1_7271_11912 1.074286e+00
R1213 n1_7271_11912 n1_9333_11912 1.178286e+01
R1214 n1_9333_11912 n1_9521_11912 1.074286e+00
R1215 n1_11583_11912 n1_11771_11912 1.074286e+00
R1216 n1_11771_11912 n1_13833_11912 1.178286e+01
R1217 n1_13833_11912 n1_14021_11912 1.074286e+00
R1218 n1_14021_11912 n1_16083_11912 1.178286e+01
R1219 n1_16083_11912 n1_16271_11912 1.074286e+00
R1220 n1_16271_11912 n1_18333_11912 1.178286e+01
R1221 n1_18333_11912 n1_18521_11912 1.074286e+00
R1222 n1_18521_11912 n1_20583_11912 1.178286e+01
R1223 n1_20583_11912 n1_20771_11912 1.074286e+00
R1224 n1_333_1112 n1_521_1112 1.074286e+00
R1225 n1_521_1112 n1_2400_1112 1.073714e+01
R1226 n1_2400_1112 n1_2583_1112 1.045714e+00
R1227 n1_2583_1112 n1_2771_1112 1.074286e+00
R1228 n1_2771_1112 n1_2864_1112 5.314286e-01
R1229 n1_2864_1112 n1_4650_1112 1.020571e+01
R1230 n1_4650_1112 n1_4833_1112 1.045714e+00
R1231 n1_4833_1112 n1_5021_1112 1.074286e+00
R1232 n1_5021_1112 n1_5114_1112 5.314286e-01
R1233 n1_5114_1112 n1_6900_1112 1.020571e+01
R1234 n1_6900_1112 n1_7083_1112 1.045714e+00
R1235 n1_7083_1112 n1_7271_1112 1.074286e+00
R1236 n1_7271_1112 n1_7364_1112 5.314286e-01
R1237 n1_7364_1112 n1_9150_1112 1.020571e+01
R1238 n1_9150_1112 n1_9333_1112 1.045714e+00
R1239 n1_9333_1112 n1_9521_1112 1.074286e+00
R1240 n1_9521_1112 n1_9614_1112 5.314286e-01
R1241 n1_11400_1112 n1_11583_1112 1.045714e+00
R1242 n1_11583_1112 n1_11771_1112 1.074286e+00
R1243 n1_11771_1112 n1_11864_1112 5.314286e-01
R1244 n1_11864_1112 n1_13650_1112 1.020571e+01
R1245 n1_13650_1112 n1_13833_1112 1.045714e+00
R1246 n1_13833_1112 n1_14021_1112 1.074286e+00
R1247 n1_14021_1112 n1_14114_1112 5.314286e-01
R1248 n1_14114_1112 n1_15900_1112 1.020571e+01
R1249 n1_15900_1112 n1_16083_1112 1.045714e+00
R1250 n1_16083_1112 n1_16271_1112 1.074286e+00
R1251 n1_16271_1112 n1_16364_1112 5.314286e-01
R1252 n1_16364_1112 n1_18150_1112 1.020571e+01
R1253 n1_18150_1112 n1_18333_1112 1.045714e+00
R1254 n1_18333_1112 n1_18521_1112 1.074286e+00
R1255 n1_18521_1112 n1_18614_1112 5.314286e-01
R1256 n1_18614_1112 n1_20583_1112 1.125143e+01
R1257 n1_20583_1112 n1_20771_1112 1.074286e+00
R1258 n1_333_1295 n1_521_1295 1.074286e+00
R1259 n1_521_1295 n1_2400_1295 1.073714e+01
R1260 n1_2400_1295 n1_2583_1295 1.045714e+00
R1261 n1_2583_1295 n1_2771_1295 1.074286e+00
R1262 n1_2771_1295 n1_2864_1295 5.314286e-01
R1263 n1_2864_1295 n1_4650_1295 1.020571e+01
R1264 n1_4650_1295 n1_4833_1295 1.045714e+00
R1265 n1_4833_1295 n1_5021_1295 1.074286e+00
R1266 n1_5021_1295 n1_5114_1295 5.314286e-01
R1267 n1_5114_1295 n1_6900_1295 1.020571e+01
R1268 n1_6900_1295 n1_7083_1295 1.045714e+00
R1269 n1_7083_1295 n1_7271_1295 1.074286e+00
R1270 n1_7271_1295 n1_7364_1295 5.314286e-01
R1271 n1_7364_1295 n1_9150_1295 1.020571e+01
R1272 n1_9150_1295 n1_9333_1295 1.045714e+00
R1273 n1_9333_1295 n1_9521_1295 1.074286e+00
R1274 n1_9521_1295 n1_9614_1295 5.314286e-01
R1275 n1_11400_1295 n1_11583_1295 1.045714e+00
R1276 n1_11583_1295 n1_11771_1295 1.074286e+00
R1277 n1_11771_1295 n1_11864_1295 5.314286e-01
R1278 n1_11864_1295 n1_13650_1295 1.020571e+01
R1279 n1_13650_1295 n1_13833_1295 1.045714e+00
R1280 n1_13833_1295 n1_14021_1295 1.074286e+00
R1281 n1_14021_1295 n1_14114_1295 5.314286e-01
R1282 n1_14114_1295 n1_15900_1295 1.020571e+01
R1283 n1_15900_1295 n1_16083_1295 1.045714e+00
R1284 n1_16083_1295 n1_16271_1295 1.074286e+00
R1285 n1_16271_1295 n1_16364_1295 5.314286e-01
R1286 n1_16364_1295 n1_18150_1295 1.020571e+01
R1287 n1_18150_1295 n1_18333_1295 1.045714e+00
R1288 n1_18333_1295 n1_18521_1295 1.074286e+00
R1289 n1_18521_1295 n1_18614_1295 5.314286e-01
R1290 n1_18614_1295 n1_20583_1295 1.125143e+01
R1291 n1_20583_1295 n1_20771_1295 1.074286e+00
R1292 n1_333_1328 n1_521_1328 1.074286e+00
R1293 n1_521_1328 n1_2400_1328 1.073714e+01
R1294 n1_2400_1328 n1_2583_1328 1.045714e+00
R1295 n1_2583_1328 n1_2771_1328 1.074286e+00
R1296 n1_2771_1328 n1_2864_1328 5.314286e-01
R1297 n1_2864_1328 n1_4650_1328 1.020571e+01
R1298 n1_4650_1328 n1_4833_1328 1.045714e+00
R1299 n1_4833_1328 n1_5021_1328 1.074286e+00
R1300 n1_5021_1328 n1_5114_1328 5.314286e-01
R1301 n1_5114_1328 n1_6900_1328 1.020571e+01
R1302 n1_6900_1328 n1_7083_1328 1.045714e+00
R1303 n1_7083_1328 n1_7271_1328 1.074286e+00
R1304 n1_7271_1328 n1_7364_1328 5.314286e-01
R1305 n1_7364_1328 n1_9150_1328 1.020571e+01
R1306 n1_9150_1328 n1_9333_1328 1.045714e+00
R1307 n1_9333_1328 n1_9521_1328 1.074286e+00
R1308 n1_9521_1328 n1_9614_1328 5.314286e-01
R1309 n1_11400_1328 n1_11583_1328 1.045714e+00
R1310 n1_11583_1328 n1_11771_1328 1.074286e+00
R1311 n1_11771_1328 n1_11864_1328 5.314286e-01
R1312 n1_11864_1328 n1_13650_1328 1.020571e+01
R1313 n1_13650_1328 n1_13833_1328 1.045714e+00
R1314 n1_13833_1328 n1_14021_1328 1.074286e+00
R1315 n1_14021_1328 n1_14114_1328 5.314286e-01
R1316 n1_14114_1328 n1_15900_1328 1.020571e+01
R1317 n1_15900_1328 n1_16083_1328 1.045714e+00
R1318 n1_16083_1328 n1_16271_1328 1.074286e+00
R1319 n1_16271_1328 n1_16364_1328 5.314286e-01
R1320 n1_16364_1328 n1_18150_1328 1.020571e+01
R1321 n1_18150_1328 n1_18333_1328 1.045714e+00
R1322 n1_18333_1328 n1_18521_1328 1.074286e+00
R1323 n1_18521_1328 n1_18614_1328 5.314286e-01
R1324 n1_18614_1328 n1_20583_1328 1.125143e+01
R1325 n1_20583_1328 n1_20771_1328 1.074286e+00
R1326 n1_521_1511 n1_2400_1511 1.073714e+01
R1327 n1_2400_1511 n1_2771_1511 2.120000e+00
R1328 n1_2771_1511 n1_2864_1511 5.314286e-01
R1329 n1_2864_1511 n1_4650_1511 1.020571e+01
R1330 n1_4650_1511 n1_5021_1511 2.120000e+00
R1331 n1_5021_1511 n1_5114_1511 5.314286e-01
R1332 n1_5114_1511 n1_6900_1511 1.020571e+01
R1333 n1_6900_1511 n1_7271_1511 2.120000e+00
R1334 n1_7271_1511 n1_7364_1511 5.314286e-01
R1335 n1_7364_1511 n1_9150_1511 1.020571e+01
R1336 n1_9150_1511 n1_9521_1511 2.120000e+00
R1337 n1_9521_1511 n1_9614_1511 5.314286e-01
R1338 n1_11400_1511 n1_11771_1511 2.120000e+00
R1339 n1_11771_1511 n1_11864_1511 5.314286e-01
R1340 n1_11864_1511 n1_13650_1511 1.020571e+01
R1341 n1_13650_1511 n1_14021_1511 2.120000e+00
R1342 n1_14021_1511 n1_14114_1511 5.314286e-01
R1343 n1_14114_1511 n1_15900_1511 1.020571e+01
R1344 n1_15900_1511 n1_16271_1511 2.120000e+00
R1345 n1_16271_1511 n1_16364_1511 5.314286e-01
R1346 n1_16364_1511 n1_18150_1511 1.020571e+01
R1347 n1_18150_1511 n1_18521_1511 2.120000e+00
R1348 n1_18521_1511 n1_18614_1511 5.314286e-01
R1349 n1_18614_1511 n1_20771_1511 1.232571e+01
R1350 n1_521_1544 n1_2400_1544 1.073714e+01
R1351 n1_2400_1544 n1_2771_1544 2.120000e+00
R1352 n1_2771_1544 n1_2864_1544 5.314286e-01
R1353 n1_2864_1544 n1_4650_1544 1.020571e+01
R1354 n1_4650_1544 n1_5021_1544 2.120000e+00
R1355 n1_5021_1544 n1_5114_1544 5.314286e-01
R1356 n1_5114_1544 n1_6900_1544 1.020571e+01
R1357 n1_6900_1544 n1_7271_1544 2.120000e+00
R1358 n1_7271_1544 n1_7364_1544 5.314286e-01
R1359 n1_7364_1544 n1_9150_1544 1.020571e+01
R1360 n1_9150_1544 n1_9521_1544 2.120000e+00
R1361 n1_9521_1544 n1_9614_1544 5.314286e-01
R1362 n1_11400_1544 n1_11771_1544 2.120000e+00
R1363 n1_11771_1544 n1_11864_1544 5.314286e-01
R1364 n1_11864_1544 n1_13650_1544 1.020571e+01
R1365 n1_13650_1544 n1_14021_1544 2.120000e+00
R1366 n1_14021_1544 n1_14114_1544 5.314286e-01
R1367 n1_14114_1544 n1_15900_1544 1.020571e+01
R1368 n1_15900_1544 n1_16271_1544 2.120000e+00
R1369 n1_16271_1544 n1_16364_1544 5.314286e-01
R1370 n1_16364_1544 n1_18150_1544 1.020571e+01
R1371 n1_18150_1544 n1_18521_1544 2.120000e+00
R1372 n1_18521_1544 n1_18614_1544 5.314286e-01
R1373 n1_18614_1544 n1_20771_1544 1.232571e+01
R1374 n1_333_1727 n1_521_1727 1.074286e+00
R1375 n1_521_1727 n1_2400_1727 1.073714e+01
R1376 n1_2400_1727 n1_2583_1727 1.045714e+00
R1377 n1_2583_1727 n1_2771_1727 1.074286e+00
R1378 n1_2771_1727 n1_2864_1727 5.314286e-01
R1379 n1_2864_1727 n1_4650_1727 1.020571e+01
R1380 n1_4650_1727 n1_4833_1727 1.045714e+00
R1381 n1_4833_1727 n1_5021_1727 1.074286e+00
R1382 n1_5021_1727 n1_5114_1727 5.314286e-01
R1383 n1_5114_1727 n1_6900_1727 1.020571e+01
R1384 n1_6900_1727 n1_7083_1727 1.045714e+00
R1385 n1_7083_1727 n1_7271_1727 1.074286e+00
R1386 n1_7271_1727 n1_7364_1727 5.314286e-01
R1387 n1_7364_1727 n1_9150_1727 1.020571e+01
R1388 n1_9150_1727 n1_9333_1727 1.045714e+00
R1389 n1_9333_1727 n1_9521_1727 1.074286e+00
R1390 n1_9521_1727 n1_9614_1727 5.314286e-01
R1391 n1_11400_1727 n1_11583_1727 1.045714e+00
R1392 n1_11583_1727 n1_11771_1727 1.074286e+00
R1393 n1_11771_1727 n1_11864_1727 5.314286e-01
R1394 n1_11864_1727 n1_13650_1727 1.020571e+01
R1395 n1_13650_1727 n1_13833_1727 1.045714e+00
R1396 n1_13833_1727 n1_14021_1727 1.074286e+00
R1397 n1_14021_1727 n1_14114_1727 5.314286e-01
R1398 n1_14114_1727 n1_15900_1727 1.020571e+01
R1399 n1_15900_1727 n1_16083_1727 1.045714e+00
R1400 n1_16083_1727 n1_16271_1727 1.074286e+00
R1401 n1_16271_1727 n1_16364_1727 5.314286e-01
R1402 n1_16364_1727 n1_18150_1727 1.020571e+01
R1403 n1_18150_1727 n1_18333_1727 1.045714e+00
R1404 n1_18333_1727 n1_18521_1727 1.074286e+00
R1405 n1_18521_1727 n1_18614_1727 5.314286e-01
R1406 n1_18614_1727 n1_20583_1727 1.125143e+01
R1407 n1_20583_1727 n1_20771_1727 1.074286e+00
R1408 n1_333_1760 n1_521_1760 1.074286e+00
R1409 n1_521_1760 n1_2400_1760 1.073714e+01
R1410 n1_2400_1760 n1_2583_1760 1.045714e+00
R1411 n1_2583_1760 n1_2771_1760 1.074286e+00
R1412 n1_2771_1760 n1_2864_1760 5.314286e-01
R1413 n1_2864_1760 n1_4650_1760 1.020571e+01
R1414 n1_4650_1760 n1_4833_1760 1.045714e+00
R1415 n1_4833_1760 n1_5021_1760 1.074286e+00
R1416 n1_5021_1760 n1_5114_1760 5.314286e-01
R1417 n1_5114_1760 n1_6900_1760 1.020571e+01
R1418 n1_6900_1760 n1_7083_1760 1.045714e+00
R1419 n1_7083_1760 n1_7271_1760 1.074286e+00
R1420 n1_7271_1760 n1_7364_1760 5.314286e-01
R1421 n1_7364_1760 n1_9150_1760 1.020571e+01
R1422 n1_9150_1760 n1_9333_1760 1.045714e+00
R1423 n1_9333_1760 n1_9521_1760 1.074286e+00
R1424 n1_9521_1760 n1_9614_1760 5.314286e-01
R1425 n1_11400_1760 n1_11583_1760 1.045714e+00
R1426 n1_11583_1760 n1_11771_1760 1.074286e+00
R1427 n1_11771_1760 n1_11864_1760 5.314286e-01
R1428 n1_11864_1760 n1_13650_1760 1.020571e+01
R1429 n1_13650_1760 n1_13833_1760 1.045714e+00
R1430 n1_13833_1760 n1_14021_1760 1.074286e+00
R1431 n1_14021_1760 n1_14114_1760 5.314286e-01
R1432 n1_14114_1760 n1_15900_1760 1.020571e+01
R1433 n1_15900_1760 n1_16083_1760 1.045714e+00
R1434 n1_16083_1760 n1_16271_1760 1.074286e+00
R1435 n1_16271_1760 n1_16364_1760 5.314286e-01
R1436 n1_16364_1760 n1_18150_1760 1.020571e+01
R1437 n1_18150_1760 n1_18333_1760 1.045714e+00
R1438 n1_18333_1760 n1_18521_1760 1.074286e+00
R1439 n1_18521_1760 n1_18614_1760 5.314286e-01
R1440 n1_18614_1760 n1_20583_1760 1.125143e+01
R1441 n1_20583_1760 n1_20771_1760 1.074286e+00
R1442 n1_333_1943 n1_521_1943 1.074286e+00
R1443 n1_521_1943 n1_2400_1943 1.073714e+01
R1444 n1_2400_1943 n1_2583_1943 1.045714e+00
R1445 n1_2583_1943 n1_2771_1943 1.074286e+00
R1446 n1_2771_1943 n1_2864_1943 5.314286e-01
R1447 n1_2864_1943 n1_4650_1943 1.020571e+01
R1448 n1_4650_1943 n1_4833_1943 1.045714e+00
R1449 n1_4833_1943 n1_5021_1943 1.074286e+00
R1450 n1_5021_1943 n1_5114_1943 5.314286e-01
R1451 n1_5114_1943 n1_6900_1943 1.020571e+01
R1452 n1_6900_1943 n1_7083_1943 1.045714e+00
R1453 n1_7083_1943 n1_7271_1943 1.074286e+00
R1454 n1_7271_1943 n1_7364_1943 5.314286e-01
R1455 n1_7364_1943 n1_9150_1943 1.020571e+01
R1456 n1_9150_1943 n1_9333_1943 1.045714e+00
R1457 n1_9333_1943 n1_9521_1943 1.074286e+00
R1458 n1_9521_1943 n1_9614_1943 5.314286e-01
R1459 n1_11400_1943 n1_11583_1943 1.045714e+00
R1460 n1_11583_1943 n1_11771_1943 1.074286e+00
R1461 n1_11771_1943 n1_11864_1943 5.314286e-01
R1462 n1_11864_1943 n1_13650_1943 1.020571e+01
R1463 n1_13650_1943 n1_13833_1943 1.045714e+00
R1464 n1_13833_1943 n1_14021_1943 1.074286e+00
R1465 n1_14021_1943 n1_14114_1943 5.314286e-01
R1466 n1_14114_1943 n1_15900_1943 1.020571e+01
R1467 n1_15900_1943 n1_16083_1943 1.045714e+00
R1468 n1_16083_1943 n1_16271_1943 1.074286e+00
R1469 n1_16271_1943 n1_16364_1943 5.314286e-01
R1470 n1_16364_1943 n1_18150_1943 1.020571e+01
R1471 n1_18150_1943 n1_18333_1943 1.045714e+00
R1472 n1_18333_1943 n1_18521_1943 1.074286e+00
R1473 n1_18521_1943 n1_18614_1943 5.314286e-01
R1474 n1_18614_1943 n1_20583_1943 1.125143e+01
R1475 n1_20583_1943 n1_20771_1943 1.074286e+00
R1476 n1_333_1976 n1_521_1976 1.074286e+00
R1477 n1_521_1976 n1_2400_1976 1.073714e+01
R1478 n1_2400_1976 n1_2583_1976 1.045714e+00
R1479 n1_2583_1976 n1_2771_1976 1.074286e+00
R1480 n1_2771_1976 n1_2864_1976 5.314286e-01
R1481 n1_2864_1976 n1_4650_1976 1.020571e+01
R1482 n1_4650_1976 n1_4833_1976 1.045714e+00
R1483 n1_4833_1976 n1_5021_1976 1.074286e+00
R1484 n1_5021_1976 n1_5114_1976 5.314286e-01
R1485 n1_5114_1976 n1_6900_1976 1.020571e+01
R1486 n1_6900_1976 n1_7083_1976 1.045714e+00
R1487 n1_7083_1976 n1_7271_1976 1.074286e+00
R1488 n1_7271_1976 n1_7364_1976 5.314286e-01
R1489 n1_7364_1976 n1_9150_1976 1.020571e+01
R1490 n1_9150_1976 n1_9333_1976 1.045714e+00
R1491 n1_9333_1976 n1_9521_1976 1.074286e+00
R1492 n1_9521_1976 n1_9614_1976 5.314286e-01
R1493 n1_11400_1976 n1_11583_1976 1.045714e+00
R1494 n1_11583_1976 n1_11771_1976 1.074286e+00
R1495 n1_11771_1976 n1_11864_1976 5.314286e-01
R1496 n1_11864_1976 n1_13650_1976 1.020571e+01
R1497 n1_13650_1976 n1_13833_1976 1.045714e+00
R1498 n1_13833_1976 n1_14021_1976 1.074286e+00
R1499 n1_14021_1976 n1_14114_1976 5.314286e-01
R1500 n1_14114_1976 n1_15900_1976 1.020571e+01
R1501 n1_15900_1976 n1_16083_1976 1.045714e+00
R1502 n1_16083_1976 n1_16271_1976 1.074286e+00
R1503 n1_16271_1976 n1_16364_1976 5.314286e-01
R1504 n1_16364_1976 n1_18150_1976 1.020571e+01
R1505 n1_18150_1976 n1_18333_1976 1.045714e+00
R1506 n1_18333_1976 n1_18521_1976 1.074286e+00
R1507 n1_18521_1976 n1_18614_1976 5.314286e-01
R1508 n1_18614_1976 n1_20583_1976 1.125143e+01
R1509 n1_20583_1976 n1_20771_1976 1.074286e+00
R1510 n1_333_2159 n1_521_2159 1.074286e+00
R1511 n1_521_2159 n1_2400_2159 1.073714e+01
R1512 n1_2400_2159 n1_2583_2159 1.045714e+00
R1513 n1_2583_2159 n1_2771_2159 1.074286e+00
R1514 n1_2771_2159 n1_2864_2159 5.314286e-01
R1515 n1_2864_2159 n1_4650_2159 1.020571e+01
R1516 n1_4650_2159 n1_4833_2159 1.045714e+00
R1517 n1_4833_2159 n1_5021_2159 1.074286e+00
R1518 n1_5021_2159 n1_5114_2159 5.314286e-01
R1519 n1_5114_2159 n1_6900_2159 1.020571e+01
R1520 n1_6900_2159 n1_7083_2159 1.045714e+00
R1521 n1_7083_2159 n1_7271_2159 1.074286e+00
R1522 n1_7271_2159 n1_7364_2159 5.314286e-01
R1523 n1_7364_2159 n1_9150_2159 1.020571e+01
R1524 n1_9150_2159 n1_9333_2159 1.045714e+00
R1525 n1_9333_2159 n1_9521_2159 1.074286e+00
R1526 n1_9521_2159 n1_9614_2159 5.314286e-01
R1527 n1_11400_2159 n1_11583_2159 1.045714e+00
R1528 n1_11583_2159 n1_11771_2159 1.074286e+00
R1529 n1_11771_2159 n1_11864_2159 5.314286e-01
R1530 n1_11864_2159 n1_13650_2159 1.020571e+01
R1531 n1_13650_2159 n1_13833_2159 1.045714e+00
R1532 n1_13833_2159 n1_14021_2159 1.074286e+00
R1533 n1_14021_2159 n1_14114_2159 5.314286e-01
R1534 n1_14114_2159 n1_15900_2159 1.020571e+01
R1535 n1_15900_2159 n1_16083_2159 1.045714e+00
R1536 n1_16083_2159 n1_16271_2159 1.074286e+00
R1537 n1_16271_2159 n1_16364_2159 5.314286e-01
R1538 n1_16364_2159 n1_18150_2159 1.020571e+01
R1539 n1_18150_2159 n1_18333_2159 1.045714e+00
R1540 n1_18333_2159 n1_18521_2159 1.074286e+00
R1541 n1_18521_2159 n1_18614_2159 5.314286e-01
R1542 n1_18614_2159 n1_20583_2159 1.125143e+01
R1543 n1_20583_2159 n1_20771_2159 1.074286e+00
R1544 n1_333_2192 n1_521_2192 1.074286e+00
R1545 n1_521_2192 n1_2400_2192 1.073714e+01
R1546 n1_2400_2192 n1_2583_2192 1.045714e+00
R1547 n1_2583_2192 n1_2771_2192 1.074286e+00
R1548 n1_2771_2192 n1_2864_2192 5.314286e-01
R1549 n1_2864_2192 n1_4650_2192 1.020571e+01
R1550 n1_4650_2192 n1_4833_2192 1.045714e+00
R1551 n1_4833_2192 n1_5021_2192 1.074286e+00
R1552 n1_5021_2192 n1_5114_2192 5.314286e-01
R1553 n1_5114_2192 n1_6900_2192 1.020571e+01
R1554 n1_6900_2192 n1_7083_2192 1.045714e+00
R1555 n1_7083_2192 n1_7271_2192 1.074286e+00
R1556 n1_7271_2192 n1_7364_2192 5.314286e-01
R1557 n1_7364_2192 n1_9150_2192 1.020571e+01
R1558 n1_9150_2192 n1_9333_2192 1.045714e+00
R1559 n1_9333_2192 n1_9521_2192 1.074286e+00
R1560 n1_9521_2192 n1_9614_2192 5.314286e-01
R1561 n1_11400_2192 n1_11583_2192 1.045714e+00
R1562 n1_11583_2192 n1_11771_2192 1.074286e+00
R1563 n1_11771_2192 n1_11864_2192 5.314286e-01
R1564 n1_11864_2192 n1_13650_2192 1.020571e+01
R1565 n1_13650_2192 n1_13833_2192 1.045714e+00
R1566 n1_13833_2192 n1_14021_2192 1.074286e+00
R1567 n1_14021_2192 n1_14114_2192 5.314286e-01
R1568 n1_14114_2192 n1_15900_2192 1.020571e+01
R1569 n1_15900_2192 n1_16083_2192 1.045714e+00
R1570 n1_16083_2192 n1_16271_2192 1.074286e+00
R1571 n1_16271_2192 n1_16364_2192 5.314286e-01
R1572 n1_16364_2192 n1_18150_2192 1.020571e+01
R1573 n1_18150_2192 n1_18333_2192 1.045714e+00
R1574 n1_18333_2192 n1_18521_2192 1.074286e+00
R1575 n1_18521_2192 n1_18614_2192 5.314286e-01
R1576 n1_18614_2192 n1_20583_2192 1.125143e+01
R1577 n1_20583_2192 n1_20771_2192 1.074286e+00
R1578 n1_333_2375 n1_521_2375 1.074286e+00
R1579 n1_521_2375 n1_2400_2375 1.073714e+01
R1580 n1_2400_2375 n1_2583_2375 1.045714e+00
R1581 n1_2583_2375 n1_2771_2375 1.074286e+00
R1582 n1_2771_2375 n1_2864_2375 5.314286e-01
R1583 n1_2864_2375 n1_4650_2375 1.020571e+01
R1584 n1_4650_2375 n1_4833_2375 1.045714e+00
R1585 n1_4833_2375 n1_5021_2375 1.074286e+00
R1586 n1_5021_2375 n1_5114_2375 5.314286e-01
R1587 n1_5114_2375 n1_6900_2375 1.020571e+01
R1588 n1_6900_2375 n1_7083_2375 1.045714e+00
R1589 n1_7083_2375 n1_7271_2375 1.074286e+00
R1590 n1_7271_2375 n1_7364_2375 5.314286e-01
R1591 n1_7364_2375 n1_9150_2375 1.020571e+01
R1592 n1_9150_2375 n1_9333_2375 1.045714e+00
R1593 n1_9333_2375 n1_9521_2375 1.074286e+00
R1594 n1_9521_2375 n1_9614_2375 5.314286e-01
R1595 n1_11400_2375 n1_11583_2375 1.045714e+00
R1596 n1_11583_2375 n1_11771_2375 1.074286e+00
R1597 n1_11771_2375 n1_11864_2375 5.314286e-01
R1598 n1_11864_2375 n1_13650_2375 1.020571e+01
R1599 n1_13650_2375 n1_13833_2375 1.045714e+00
R1600 n1_13833_2375 n1_14021_2375 1.074286e+00
R1601 n1_14021_2375 n1_14114_2375 5.314286e-01
R1602 n1_14114_2375 n1_15900_2375 1.020571e+01
R1603 n1_15900_2375 n1_16083_2375 1.045714e+00
R1604 n1_16083_2375 n1_16271_2375 1.074286e+00
R1605 n1_16271_2375 n1_16364_2375 5.314286e-01
R1606 n1_16364_2375 n1_18150_2375 1.020571e+01
R1607 n1_18150_2375 n1_18333_2375 1.045714e+00
R1608 n1_18333_2375 n1_18521_2375 1.074286e+00
R1609 n1_18521_2375 n1_18614_2375 5.314286e-01
R1610 n1_18614_2375 n1_20583_2375 1.125143e+01
R1611 n1_20583_2375 n1_20771_2375 1.074286e+00
R1612 n1_333_2408 n1_521_2408 1.074286e+00
R1613 n1_521_2408 n1_2400_2408 1.073714e+01
R1614 n1_2400_2408 n1_2583_2408 1.045714e+00
R1615 n1_2583_2408 n1_2771_2408 1.074286e+00
R1616 n1_2771_2408 n1_2864_2408 5.314286e-01
R1617 n1_2864_2408 n1_4650_2408 1.020571e+01
R1618 n1_4650_2408 n1_4833_2408 1.045714e+00
R1619 n1_4833_2408 n1_5021_2408 1.074286e+00
R1620 n1_5021_2408 n1_5114_2408 5.314286e-01
R1621 n1_5114_2408 n1_6900_2408 1.020571e+01
R1622 n1_6900_2408 n1_7083_2408 1.045714e+00
R1623 n1_7083_2408 n1_7271_2408 1.074286e+00
R1624 n1_7271_2408 n1_7364_2408 5.314286e-01
R1625 n1_7364_2408 n1_9150_2408 1.020571e+01
R1626 n1_9150_2408 n1_9333_2408 1.045714e+00
R1627 n1_9333_2408 n1_9521_2408 1.074286e+00
R1628 n1_9521_2408 n1_9614_2408 5.314286e-01
R1629 n1_11400_2408 n1_11583_2408 1.045714e+00
R1630 n1_11583_2408 n1_11771_2408 1.074286e+00
R1631 n1_11771_2408 n1_11864_2408 5.314286e-01
R1632 n1_11864_2408 n1_13650_2408 1.020571e+01
R1633 n1_13650_2408 n1_13833_2408 1.045714e+00
R1634 n1_13833_2408 n1_14021_2408 1.074286e+00
R1635 n1_14021_2408 n1_14114_2408 5.314286e-01
R1636 n1_14114_2408 n1_15900_2408 1.020571e+01
R1637 n1_15900_2408 n1_16083_2408 1.045714e+00
R1638 n1_16083_2408 n1_16271_2408 1.074286e+00
R1639 n1_16271_2408 n1_16364_2408 5.314286e-01
R1640 n1_16364_2408 n1_18150_2408 1.020571e+01
R1641 n1_18150_2408 n1_18333_2408 1.045714e+00
R1642 n1_18333_2408 n1_18521_2408 1.074286e+00
R1643 n1_18521_2408 n1_18614_2408 5.314286e-01
R1644 n1_18614_2408 n1_20583_2408 1.125143e+01
R1645 n1_20583_2408 n1_20771_2408 1.074286e+00
R1646 n1_333_2591 n1_521_2591 1.074286e+00
R1647 n1_521_2591 n1_2400_2591 1.073714e+01
R1648 n1_2400_2591 n1_2583_2591 1.045714e+00
R1649 n1_2583_2591 n1_2771_2591 1.074286e+00
R1650 n1_2771_2591 n1_2864_2591 5.314286e-01
R1651 n1_2864_2591 n1_4650_2591 1.020571e+01
R1652 n1_4650_2591 n1_4833_2591 1.045714e+00
R1653 n1_4833_2591 n1_5021_2591 1.074286e+00
R1654 n1_5021_2591 n1_5114_2591 5.314286e-01
R1655 n1_5114_2591 n1_6900_2591 1.020571e+01
R1656 n1_6900_2591 n1_7083_2591 1.045714e+00
R1657 n1_7083_2591 n1_7271_2591 1.074286e+00
R1658 n1_7271_2591 n1_7364_2591 5.314286e-01
R1659 n1_7364_2591 n1_9150_2591 1.020571e+01
R1660 n1_9150_2591 n1_9333_2591 1.045714e+00
R1661 n1_9333_2591 n1_9521_2591 1.074286e+00
R1662 n1_9521_2591 n1_9614_2591 5.314286e-01
R1663 n1_11400_2591 n1_11583_2591 1.045714e+00
R1664 n1_11583_2591 n1_11771_2591 1.074286e+00
R1665 n1_11771_2591 n1_11864_2591 5.314286e-01
R1666 n1_11864_2591 n1_13650_2591 1.020571e+01
R1667 n1_13650_2591 n1_13833_2591 1.045714e+00
R1668 n1_13833_2591 n1_14021_2591 1.074286e+00
R1669 n1_14021_2591 n1_14114_2591 5.314286e-01
R1670 n1_14114_2591 n1_15900_2591 1.020571e+01
R1671 n1_15900_2591 n1_16083_2591 1.045714e+00
R1672 n1_16083_2591 n1_16271_2591 1.074286e+00
R1673 n1_16271_2591 n1_16364_2591 5.314286e-01
R1674 n1_16364_2591 n1_18150_2591 1.020571e+01
R1675 n1_18150_2591 n1_18333_2591 1.045714e+00
R1676 n1_18333_2591 n1_18521_2591 1.074286e+00
R1677 n1_18521_2591 n1_18614_2591 5.314286e-01
R1678 n1_18614_2591 n1_20583_2591 1.125143e+01
R1679 n1_20583_2591 n1_20771_2591 1.074286e+00
R1680 n1_333_2624 n1_521_2624 1.074286e+00
R1681 n1_521_2624 n1_2400_2624 1.073714e+01
R1682 n1_2400_2624 n1_2583_2624 1.045714e+00
R1683 n1_2583_2624 n1_2771_2624 1.074286e+00
R1684 n1_2771_2624 n1_2864_2624 5.314286e-01
R1685 n1_2864_2624 n1_4650_2624 1.020571e+01
R1686 n1_4650_2624 n1_4833_2624 1.045714e+00
R1687 n1_4833_2624 n1_5021_2624 1.074286e+00
R1688 n1_5021_2624 n1_5114_2624 5.314286e-01
R1689 n1_5114_2624 n1_6900_2624 1.020571e+01
R1690 n1_6900_2624 n1_7083_2624 1.045714e+00
R1691 n1_7083_2624 n1_7271_2624 1.074286e+00
R1692 n1_7271_2624 n1_7364_2624 5.314286e-01
R1693 n1_7364_2624 n1_9150_2624 1.020571e+01
R1694 n1_9150_2624 n1_9333_2624 1.045714e+00
R1695 n1_9333_2624 n1_9521_2624 1.074286e+00
R1696 n1_9521_2624 n1_9614_2624 5.314286e-01
R1697 n1_11400_2624 n1_11583_2624 1.045714e+00
R1698 n1_11583_2624 n1_11771_2624 1.074286e+00
R1699 n1_11771_2624 n1_11864_2624 5.314286e-01
R1700 n1_11864_2624 n1_13650_2624 1.020571e+01
R1701 n1_13650_2624 n1_13833_2624 1.045714e+00
R1702 n1_13833_2624 n1_14021_2624 1.074286e+00
R1703 n1_14021_2624 n1_14114_2624 5.314286e-01
R1704 n1_14114_2624 n1_15900_2624 1.020571e+01
R1705 n1_15900_2624 n1_16083_2624 1.045714e+00
R1706 n1_16083_2624 n1_16271_2624 1.074286e+00
R1707 n1_16271_2624 n1_16364_2624 5.314286e-01
R1708 n1_16364_2624 n1_18150_2624 1.020571e+01
R1709 n1_18150_2624 n1_18333_2624 1.045714e+00
R1710 n1_18333_2624 n1_18521_2624 1.074286e+00
R1711 n1_18521_2624 n1_18614_2624 5.314286e-01
R1712 n1_18614_2624 n1_20583_2624 1.125143e+01
R1713 n1_20583_2624 n1_20771_2624 1.074286e+00
R1714 n1_333_2807 n1_521_2807 1.074286e+00
R1715 n1_521_2807 n1_2583_2807 1.178286e+01
R1716 n1_2583_2807 n1_2771_2807 1.074286e+00
R1717 n1_2771_2807 n1_4833_2807 1.178286e+01
R1718 n1_4833_2807 n1_5021_2807 1.074286e+00
R1719 n1_5021_2807 n1_7083_2807 1.178286e+01
R1720 n1_7083_2807 n1_7271_2807 1.074286e+00
R1721 n1_7271_2807 n1_9333_2807 1.178286e+01
R1722 n1_9333_2807 n1_9521_2807 1.074286e+00
R1723 n1_11583_2807 n1_11771_2807 1.074286e+00
R1724 n1_11771_2807 n1_13833_2807 1.178286e+01
R1725 n1_13833_2807 n1_14021_2807 1.074286e+00
R1726 n1_14021_2807 n1_16083_2807 1.178286e+01
R1727 n1_16083_2807 n1_16271_2807 1.074286e+00
R1728 n1_16271_2807 n1_18333_2807 1.178286e+01
R1729 n1_18333_2807 n1_18521_2807 1.074286e+00
R1730 n1_18521_2807 n1_20583_2807 1.178286e+01
R1731 n1_20583_2807 n1_20771_2807 1.074286e+00
R1732 n1_333_2840 n1_521_2840 1.074286e+00
R1733 n1_521_2840 n1_2583_2840 1.178286e+01
R1734 n1_2583_2840 n1_2771_2840 1.074286e+00
R1735 n1_2771_2840 n1_4833_2840 1.178286e+01
R1736 n1_4833_2840 n1_5021_2840 1.074286e+00
R1737 n1_5021_2840 n1_7083_2840 1.178286e+01
R1738 n1_7083_2840 n1_7271_2840 1.074286e+00
R1739 n1_7271_2840 n1_9333_2840 1.178286e+01
R1740 n1_9333_2840 n1_9521_2840 1.074286e+00
R1741 n1_11583_2840 n1_11771_2840 1.074286e+00
R1742 n1_11771_2840 n1_13833_2840 1.178286e+01
R1743 n1_13833_2840 n1_14021_2840 1.074286e+00
R1744 n1_14021_2840 n1_16083_2840 1.178286e+01
R1745 n1_16083_2840 n1_16271_2840 1.074286e+00
R1746 n1_16271_2840 n1_18333_2840 1.178286e+01
R1747 n1_18333_2840 n1_18521_2840 1.074286e+00
R1748 n1_18521_2840 n1_20583_2840 1.178286e+01
R1749 n1_20583_2840 n1_20771_2840 1.074286e+00
R1750 n1_333_3023 n1_521_3023 1.074286e+00
R1751 n1_521_3023 n1_2583_3023 1.178286e+01
R1752 n1_2583_3023 n1_2771_3023 1.074286e+00
R1753 n1_2771_3023 n1_4833_3023 1.178286e+01
R1754 n1_4833_3023 n1_5021_3023 1.074286e+00
R1755 n1_5021_3023 n1_7083_3023 1.178286e+01
R1756 n1_7083_3023 n1_7271_3023 1.074286e+00
R1757 n1_7271_3023 n1_9333_3023 1.178286e+01
R1758 n1_9333_3023 n1_9521_3023 1.074286e+00
R1759 n1_11583_3023 n1_11771_3023 1.074286e+00
R1760 n1_11771_3023 n1_13833_3023 1.178286e+01
R1761 n1_13833_3023 n1_14021_3023 1.074286e+00
R1762 n1_14021_3023 n1_16083_3023 1.178286e+01
R1763 n1_16083_3023 n1_16271_3023 1.074286e+00
R1764 n1_16271_3023 n1_18333_3023 1.178286e+01
R1765 n1_18333_3023 n1_18521_3023 1.074286e+00
R1766 n1_18521_3023 n1_20583_3023 1.178286e+01
R1767 n1_20583_3023 n1_20771_3023 1.074286e+00
R1768 n1_333_3056 n1_521_3056 1.074286e+00
R1769 n1_521_3056 n1_2583_3056 1.178286e+01
R1770 n1_2583_3056 n1_2771_3056 1.074286e+00
R1771 n1_2771_3056 n1_4833_3056 1.178286e+01
R1772 n1_4833_3056 n1_5021_3056 1.074286e+00
R1773 n1_5021_3056 n1_7083_3056 1.178286e+01
R1774 n1_7083_3056 n1_7271_3056 1.074286e+00
R1775 n1_7271_3056 n1_9333_3056 1.178286e+01
R1776 n1_9333_3056 n1_9521_3056 1.074286e+00
R1777 n1_11583_3056 n1_11771_3056 1.074286e+00
R1778 n1_11771_3056 n1_13833_3056 1.178286e+01
R1779 n1_13833_3056 n1_14021_3056 1.074286e+00
R1780 n1_14021_3056 n1_16083_3056 1.178286e+01
R1781 n1_16083_3056 n1_16271_3056 1.074286e+00
R1782 n1_16271_3056 n1_18333_3056 1.178286e+01
R1783 n1_18333_3056 n1_18521_3056 1.074286e+00
R1784 n1_18521_3056 n1_20583_3056 1.178286e+01
R1785 n1_20583_3056 n1_20771_3056 1.074286e+00
R1786 n1_333_3239 n1_521_3239 1.074286e+00
R1787 n1_521_3239 n1_2583_3239 1.178286e+01
R1788 n1_2583_3239 n1_2771_3239 1.074286e+00
R1789 n1_2771_3239 n1_4833_3239 1.178286e+01
R1790 n1_4833_3239 n1_5021_3239 1.074286e+00
R1791 n1_5021_3239 n1_7083_3239 1.178286e+01
R1792 n1_7083_3239 n1_7271_3239 1.074286e+00
R1793 n1_7271_3239 n1_9333_3239 1.178286e+01
R1794 n1_9333_3239 n1_9521_3239 1.074286e+00
R1795 n1_11583_3239 n1_11771_3239 1.074286e+00
R1796 n1_11771_3239 n1_13833_3239 1.178286e+01
R1797 n1_13833_3239 n1_14021_3239 1.074286e+00
R1798 n1_14021_3239 n1_16083_3239 1.178286e+01
R1799 n1_16083_3239 n1_16271_3239 1.074286e+00
R1800 n1_16271_3239 n1_18333_3239 1.178286e+01
R1801 n1_18333_3239 n1_18521_3239 1.074286e+00
R1802 n1_18521_3239 n1_20583_3239 1.178286e+01
R1803 n1_20583_3239 n1_20771_3239 1.074286e+00
R1804 n1_333_3272 n1_521_3272 1.074286e+00
R1805 n1_521_3272 n1_2583_3272 1.178286e+01
R1806 n1_2583_3272 n1_2771_3272 1.074286e+00
R1807 n1_2771_3272 n1_4833_3272 1.178286e+01
R1808 n1_4833_3272 n1_5021_3272 1.074286e+00
R1809 n1_5021_3272 n1_7083_3272 1.178286e+01
R1810 n1_7083_3272 n1_7271_3272 1.074286e+00
R1811 n1_7271_3272 n1_9333_3272 1.178286e+01
R1812 n1_9333_3272 n1_9521_3272 1.074286e+00
R1813 n1_11583_3272 n1_11771_3272 1.074286e+00
R1814 n1_11771_3272 n1_13833_3272 1.178286e+01
R1815 n1_13833_3272 n1_14021_3272 1.074286e+00
R1816 n1_14021_3272 n1_16083_3272 1.178286e+01
R1817 n1_16083_3272 n1_16271_3272 1.074286e+00
R1818 n1_16271_3272 n1_18333_3272 1.178286e+01
R1819 n1_18333_3272 n1_18521_3272 1.074286e+00
R1820 n1_18521_3272 n1_20583_3272 1.178286e+01
R1821 n1_20583_3272 n1_20771_3272 1.074286e+00
R1822 n1_333_3455 n1_521_3455 1.074286e+00
R1823 n1_521_3455 n1_2583_3455 1.178286e+01
R1824 n1_2583_3455 n1_2771_3455 1.074286e+00
R1825 n1_2771_3455 n1_4833_3455 1.178286e+01
R1826 n1_4833_3455 n1_5021_3455 1.074286e+00
R1827 n1_5021_3455 n1_7083_3455 1.178286e+01
R1828 n1_7083_3455 n1_7271_3455 1.074286e+00
R1829 n1_7271_3455 n1_9333_3455 1.178286e+01
R1830 n1_9333_3455 n1_9521_3455 1.074286e+00
R1831 n1_11583_3455 n1_11771_3455 1.074286e+00
R1832 n1_11771_3455 n1_13833_3455 1.178286e+01
R1833 n1_13833_3455 n1_14021_3455 1.074286e+00
R1834 n1_14021_3455 n1_16083_3455 1.178286e+01
R1835 n1_16083_3455 n1_16271_3455 1.074286e+00
R1836 n1_16271_3455 n1_18333_3455 1.178286e+01
R1837 n1_18333_3455 n1_18521_3455 1.074286e+00
R1838 n1_18521_3455 n1_20583_3455 1.178286e+01
R1839 n1_20583_3455 n1_20771_3455 1.074286e+00
R1840 n1_333_3488 n1_521_3488 1.074286e+00
R1841 n1_521_3488 n1_2583_3488 1.178286e+01
R1842 n1_2583_3488 n1_2771_3488 1.074286e+00
R1843 n1_2771_3488 n1_4833_3488 1.178286e+01
R1844 n1_4833_3488 n1_5021_3488 1.074286e+00
R1845 n1_5021_3488 n1_7083_3488 1.178286e+01
R1846 n1_7083_3488 n1_7271_3488 1.074286e+00
R1847 n1_7271_3488 n1_9333_3488 1.178286e+01
R1848 n1_9333_3488 n1_9521_3488 1.074286e+00
R1849 n1_11583_3488 n1_11771_3488 1.074286e+00
R1850 n1_11771_3488 n1_13833_3488 1.178286e+01
R1851 n1_13833_3488 n1_14021_3488 1.074286e+00
R1852 n1_14021_3488 n1_16083_3488 1.178286e+01
R1853 n1_16083_3488 n1_16271_3488 1.074286e+00
R1854 n1_16271_3488 n1_18333_3488 1.178286e+01
R1855 n1_18333_3488 n1_18521_3488 1.074286e+00
R1856 n1_18521_3488 n1_20583_3488 1.178286e+01
R1857 n1_20583_3488 n1_20771_3488 1.074286e+00
R1858 n1_333_3671 n1_521_3671 1.074286e+00
R1859 n1_521_3671 n1_2583_3671 1.178286e+01
R1860 n1_2583_3671 n1_2771_3671 1.074286e+00
R1861 n1_2771_3671 n1_4833_3671 1.178286e+01
R1862 n1_4833_3671 n1_5021_3671 1.074286e+00
R1863 n1_5021_3671 n1_7083_3671 1.178286e+01
R1864 n1_7083_3671 n1_7271_3671 1.074286e+00
R1865 n1_7271_3671 n1_9333_3671 1.178286e+01
R1866 n1_9333_3671 n1_9521_3671 1.074286e+00
R1867 n1_11583_3671 n1_11771_3671 1.074286e+00
R1868 n1_11771_3671 n1_13833_3671 1.178286e+01
R1869 n1_13833_3671 n1_14021_3671 1.074286e+00
R1870 n1_14021_3671 n1_16083_3671 1.178286e+01
R1871 n1_16083_3671 n1_16271_3671 1.074286e+00
R1872 n1_16271_3671 n1_18333_3671 1.178286e+01
R1873 n1_18333_3671 n1_18521_3671 1.074286e+00
R1874 n1_18521_3671 n1_20583_3671 1.178286e+01
R1875 n1_20583_3671 n1_20771_3671 1.074286e+00
R1876 n1_333_3704 n1_521_3704 1.074286e+00
R1877 n1_521_3704 n1_2583_3704 1.178286e+01
R1878 n1_2583_3704 n1_2771_3704 1.074286e+00
R1879 n1_2771_3704 n1_4833_3704 1.178286e+01
R1880 n1_4833_3704 n1_5021_3704 1.074286e+00
R1881 n1_5021_3704 n1_7083_3704 1.178286e+01
R1882 n1_7083_3704 n1_7271_3704 1.074286e+00
R1883 n1_7271_3704 n1_9333_3704 1.178286e+01
R1884 n1_9333_3704 n1_9521_3704 1.074286e+00
R1885 n1_11583_3704 n1_11771_3704 1.074286e+00
R1886 n1_11771_3704 n1_13833_3704 1.178286e+01
R1887 n1_13833_3704 n1_14021_3704 1.074286e+00
R1888 n1_14021_3704 n1_16083_3704 1.178286e+01
R1889 n1_16083_3704 n1_16271_3704 1.074286e+00
R1890 n1_16271_3704 n1_18333_3704 1.178286e+01
R1891 n1_18333_3704 n1_18521_3704 1.074286e+00
R1892 n1_18521_3704 n1_20583_3704 1.178286e+01
R1893 n1_20583_3704 n1_20771_3704 1.074286e+00
R1894 n1_521_3887 n1_2771_3887 1.285714e+01
R1895 n1_2771_3887 n1_5021_3887 1.285714e+01
R1896 n1_5021_3887 n1_7271_3887 1.285714e+01
R1897 n1_7271_3887 n1_9521_3887 1.285714e+01
R1898 n1_11771_3887 n1_14021_3887 1.285714e+01
R1899 n1_14021_3887 n1_16271_3887 1.285714e+01
R1900 n1_16271_3887 n1_18521_3887 1.285714e+01
R1901 n1_18521_3887 n1_20771_3887 1.285714e+01
R1902 n1_521_3920 n1_2771_3920 1.285714e+01
R1903 n1_2771_3920 n1_5021_3920 1.285714e+01
R1904 n1_5021_3920 n1_7271_3920 1.285714e+01
R1905 n1_7271_3920 n1_9521_3920 1.285714e+01
R1906 n1_11771_3920 n1_14021_3920 1.285714e+01
R1907 n1_14021_3920 n1_16271_3920 1.285714e+01
R1908 n1_16271_3920 n1_18521_3920 1.285714e+01
R1909 n1_18521_3920 n1_20771_3920 1.285714e+01
R1910 n1_333_4103 n1_521_4103 1.074286e+00
R1911 n1_521_4103 n1_2583_4103 1.178286e+01
R1912 n1_2583_4103 n1_2771_4103 1.074286e+00
R1913 n1_2771_4103 n1_4833_4103 1.178286e+01
R1914 n1_4833_4103 n1_5021_4103 1.074286e+00
R1915 n1_5021_4103 n1_7083_4103 1.178286e+01
R1916 n1_7083_4103 n1_7271_4103 1.074286e+00
R1917 n1_7271_4103 n1_9333_4103 1.178286e+01
R1918 n1_9333_4103 n1_9521_4103 1.074286e+00
R1919 n1_11583_4103 n1_11771_4103 1.074286e+00
R1920 n1_11771_4103 n1_13833_4103 1.178286e+01
R1921 n1_13833_4103 n1_14021_4103 1.074286e+00
R1922 n1_14021_4103 n1_16083_4103 1.178286e+01
R1923 n1_16083_4103 n1_16271_4103 1.074286e+00
R1924 n1_16271_4103 n1_18333_4103 1.178286e+01
R1925 n1_18333_4103 n1_18521_4103 1.074286e+00
R1926 n1_18521_4103 n1_20583_4103 1.178286e+01
R1927 n1_20583_4103 n1_20771_4103 1.074286e+00
R1928 n1_333_4136 n1_521_4136 1.074286e+00
R1929 n1_521_4136 n1_2583_4136 1.178286e+01
R1930 n1_2583_4136 n1_2771_4136 1.074286e+00
R1931 n1_2771_4136 n1_4833_4136 1.178286e+01
R1932 n1_4833_4136 n1_5021_4136 1.074286e+00
R1933 n1_5021_4136 n1_7083_4136 1.178286e+01
R1934 n1_7083_4136 n1_7271_4136 1.074286e+00
R1935 n1_7271_4136 n1_9333_4136 1.178286e+01
R1936 n1_9333_4136 n1_9521_4136 1.074286e+00
R1937 n1_11583_4136 n1_11771_4136 1.074286e+00
R1938 n1_11771_4136 n1_13833_4136 1.178286e+01
R1939 n1_13833_4136 n1_14021_4136 1.074286e+00
R1940 n1_14021_4136 n1_16083_4136 1.178286e+01
R1941 n1_16083_4136 n1_16271_4136 1.074286e+00
R1942 n1_16271_4136 n1_18333_4136 1.178286e+01
R1943 n1_18333_4136 n1_18521_4136 1.074286e+00
R1944 n1_18521_4136 n1_20583_4136 1.178286e+01
R1945 n1_20583_4136 n1_20771_4136 1.074286e+00
R1946 n1_333_4319 n1_521_4319 1.074286e+00
R1947 n1_521_4319 n1_2583_4319 1.178286e+01
R1948 n1_2583_4319 n1_2771_4319 1.074286e+00
R1949 n1_2771_4319 n1_4833_4319 1.178286e+01
R1950 n1_4833_4319 n1_5021_4319 1.074286e+00
R1951 n1_5021_4319 n1_7083_4319 1.178286e+01
R1952 n1_7083_4319 n1_7271_4319 1.074286e+00
R1953 n1_7271_4319 n1_9333_4319 1.178286e+01
R1954 n1_9333_4319 n1_9521_4319 1.074286e+00
R1955 n1_11583_4319 n1_11771_4319 1.074286e+00
R1956 n1_11771_4319 n1_13833_4319 1.178286e+01
R1957 n1_13833_4319 n1_14021_4319 1.074286e+00
R1958 n1_14021_4319 n1_16083_4319 1.178286e+01
R1959 n1_16083_4319 n1_16271_4319 1.074286e+00
R1960 n1_16271_4319 n1_18333_4319 1.178286e+01
R1961 n1_18333_4319 n1_18521_4319 1.074286e+00
R1962 n1_18521_4319 n1_20583_4319 1.178286e+01
R1963 n1_20583_4319 n1_20771_4319 1.074286e+00
R1964 n1_333_4352 n1_521_4352 1.074286e+00
R1965 n1_521_4352 n1_2583_4352 1.178286e+01
R1966 n1_2583_4352 n1_2771_4352 1.074286e+00
R1967 n1_2771_4352 n1_4833_4352 1.178286e+01
R1968 n1_4833_4352 n1_5021_4352 1.074286e+00
R1969 n1_5021_4352 n1_7083_4352 1.178286e+01
R1970 n1_7083_4352 n1_7271_4352 1.074286e+00
R1971 n1_7271_4352 n1_9333_4352 1.178286e+01
R1972 n1_9333_4352 n1_9521_4352 1.074286e+00
R1973 n1_11583_4352 n1_11771_4352 1.074286e+00
R1974 n1_11771_4352 n1_13833_4352 1.178286e+01
R1975 n1_13833_4352 n1_14021_4352 1.074286e+00
R1976 n1_14021_4352 n1_16083_4352 1.178286e+01
R1977 n1_16083_4352 n1_16271_4352 1.074286e+00
R1978 n1_16271_4352 n1_18333_4352 1.178286e+01
R1979 n1_18333_4352 n1_18521_4352 1.074286e+00
R1980 n1_18521_4352 n1_20583_4352 1.178286e+01
R1981 n1_20583_4352 n1_20771_4352 1.074286e+00
R1982 n1_333_4535 n1_521_4535 1.074286e+00
R1983 n1_521_4535 n1_2583_4535 1.178286e+01
R1984 n1_2583_4535 n1_2771_4535 1.074286e+00
R1985 n1_2771_4535 n1_4833_4535 1.178286e+01
R1986 n1_4833_4535 n1_5021_4535 1.074286e+00
R1987 n1_5021_4535 n1_7083_4535 1.178286e+01
R1988 n1_7083_4535 n1_7271_4535 1.074286e+00
R1989 n1_7271_4535 n1_9333_4535 1.178286e+01
R1990 n1_9333_4535 n1_9521_4535 1.074286e+00
R1991 n1_11583_4535 n1_11771_4535 1.074286e+00
R1992 n1_11771_4535 n1_13833_4535 1.178286e+01
R1993 n1_13833_4535 n1_14021_4535 1.074286e+00
R1994 n1_14021_4535 n1_16083_4535 1.178286e+01
R1995 n1_16083_4535 n1_16271_4535 1.074286e+00
R1996 n1_16271_4535 n1_18333_4535 1.178286e+01
R1997 n1_18333_4535 n1_18521_4535 1.074286e+00
R1998 n1_18521_4535 n1_20583_4535 1.178286e+01
R1999 n1_20583_4535 n1_20771_4535 1.074286e+00
R2000 n1_333_4568 n1_521_4568 1.074286e+00
R2001 n1_521_4568 n1_2583_4568 1.178286e+01
R2002 n1_2583_4568 n1_2771_4568 1.074286e+00
R2003 n1_2771_4568 n1_4833_4568 1.178286e+01
R2004 n1_4833_4568 n1_5021_4568 1.074286e+00
R2005 n1_5021_4568 n1_7083_4568 1.178286e+01
R2006 n1_7083_4568 n1_7271_4568 1.074286e+00
R2007 n1_7271_4568 n1_9333_4568 1.178286e+01
R2008 n1_9333_4568 n1_9521_4568 1.074286e+00
R2009 n1_11583_4568 n1_11771_4568 1.074286e+00
R2010 n1_11771_4568 n1_13833_4568 1.178286e+01
R2011 n1_13833_4568 n1_14021_4568 1.074286e+00
R2012 n1_14021_4568 n1_16083_4568 1.178286e+01
R2013 n1_16083_4568 n1_16271_4568 1.074286e+00
R2014 n1_16271_4568 n1_18333_4568 1.178286e+01
R2015 n1_18333_4568 n1_18521_4568 1.074286e+00
R2016 n1_18521_4568 n1_20583_4568 1.178286e+01
R2017 n1_20583_4568 n1_20771_4568 1.074286e+00
R2018 n1_333_4751 n1_521_4751 1.074286e+00
R2019 n1_521_4751 n1_2583_4751 1.178286e+01
R2020 n1_2583_4751 n1_2771_4751 1.074286e+00
R2021 n1_2771_4751 n1_4833_4751 1.178286e+01
R2022 n1_4833_4751 n1_5021_4751 1.074286e+00
R2023 n1_5021_4751 n1_7083_4751 1.178286e+01
R2024 n1_7083_4751 n1_7271_4751 1.074286e+00
R2025 n1_7271_4751 n1_9333_4751 1.178286e+01
R2026 n1_9333_4751 n1_9521_4751 1.074286e+00
R2027 n1_11583_4751 n1_11771_4751 1.074286e+00
R2028 n1_11771_4751 n1_13833_4751 1.178286e+01
R2029 n1_13833_4751 n1_14021_4751 1.074286e+00
R2030 n1_14021_4751 n1_16083_4751 1.178286e+01
R2031 n1_16083_4751 n1_16271_4751 1.074286e+00
R2032 n1_16271_4751 n1_18333_4751 1.178286e+01
R2033 n1_18333_4751 n1_18521_4751 1.074286e+00
R2034 n1_18521_4751 n1_20583_4751 1.178286e+01
R2035 n1_20583_4751 n1_20771_4751 1.074286e+00
R2036 n1_333_4784 n1_521_4784 1.074286e+00
R2037 n1_521_4784 n1_2583_4784 1.178286e+01
R2038 n1_2583_4784 n1_2771_4784 1.074286e+00
R2039 n1_2771_4784 n1_4833_4784 1.178286e+01
R2040 n1_4833_4784 n1_5021_4784 1.074286e+00
R2041 n1_5021_4784 n1_7083_4784 1.178286e+01
R2042 n1_7083_4784 n1_7271_4784 1.074286e+00
R2043 n1_7271_4784 n1_9333_4784 1.178286e+01
R2044 n1_9333_4784 n1_9521_4784 1.074286e+00
R2045 n1_11583_4784 n1_11771_4784 1.074286e+00
R2046 n1_11771_4784 n1_13833_4784 1.178286e+01
R2047 n1_13833_4784 n1_14021_4784 1.074286e+00
R2048 n1_14021_4784 n1_16083_4784 1.178286e+01
R2049 n1_16083_4784 n1_16271_4784 1.074286e+00
R2050 n1_16271_4784 n1_18333_4784 1.178286e+01
R2051 n1_18333_4784 n1_18521_4784 1.074286e+00
R2052 n1_18521_4784 n1_20583_4784 1.178286e+01
R2053 n1_20583_4784 n1_20771_4784 1.074286e+00
R2054 n1_333_4967 n1_380_4967 2.685714e-01
R2055 n1_380_4967 n1_2583_4967 1.258857e+01
R2056 n1_2583_4967 n1_2630_4967 2.685714e-01
R2057 n1_2630_4967 n1_4833_4967 1.258857e+01
R2058 n1_4833_4967 n1_4880_4967 2.685714e-01
R2059 n1_4880_4967 n1_7083_4967 1.258857e+01
R2060 n1_7083_4967 n1_7130_4967 2.685714e-01
R2061 n1_7130_4967 n1_9333_4967 1.258857e+01
R2062 n1_9333_4967 n1_9380_4967 2.685714e-01
R2063 n1_11583_4967 n1_11630_4967 2.685714e-01
R2064 n1_11630_4967 n1_13833_4967 1.258857e+01
R2065 n1_13833_4967 n1_13880_4967 2.685714e-01
R2066 n1_13880_4967 n1_16083_4967 1.258857e+01
R2067 n1_16083_4967 n1_16130_4967 2.685714e-01
R2068 n1_16130_4967 n1_18333_4967 1.258857e+01
R2069 n1_18333_4967 n1_18380_4967 2.685714e-01
R2070 n1_18380_4967 n1_20583_4967 1.258857e+01
R2071 n1_20583_4967 n1_20630_4967 2.685714e-01
R2072 n1_333_5000 n1_380_5000 2.685714e-01
R2073 n1_380_5000 n1_521_5000 8.057143e-01
R2074 n1_521_5000 n1_2583_5000 1.178286e+01
R2075 n1_2583_5000 n1_2630_5000 2.685714e-01
R2076 n1_2630_5000 n1_2771_5000 8.057143e-01
R2077 n1_2771_5000 n1_4833_5000 1.178286e+01
R2078 n1_4833_5000 n1_4880_5000 2.685714e-01
R2079 n1_4880_5000 n1_5021_5000 8.057143e-01
R2080 n1_5021_5000 n1_7083_5000 1.178286e+01
R2081 n1_7083_5000 n1_7130_5000 2.685714e-01
R2082 n1_7130_5000 n1_7271_5000 8.057143e-01
R2083 n1_7271_5000 n1_9333_5000 1.178286e+01
R2084 n1_9333_5000 n1_9380_5000 2.685714e-01
R2085 n1_9380_5000 n1_9521_5000 8.057143e-01
R2086 n1_11583_5000 n1_11630_5000 2.685714e-01
R2087 n1_11630_5000 n1_11771_5000 8.057143e-01
R2088 n1_11771_5000 n1_13833_5000 1.178286e+01
R2089 n1_13833_5000 n1_13880_5000 2.685714e-01
R2090 n1_13880_5000 n1_14021_5000 8.057143e-01
R2091 n1_14021_5000 n1_16083_5000 1.178286e+01
R2092 n1_16083_5000 n1_16130_5000 2.685714e-01
R2093 n1_16130_5000 n1_16271_5000 8.057143e-01
R2094 n1_16271_5000 n1_18333_5000 1.178286e+01
R2095 n1_18333_5000 n1_18380_5000 2.685714e-01
R2096 n1_18380_5000 n1_18521_5000 8.057143e-01
R2097 n1_18521_5000 n1_20583_5000 1.178286e+01
R2098 n1_20583_5000 n1_20630_5000 2.685714e-01
R2099 n1_20630_5000 n1_20771_5000 8.057143e-01
R2100 n1_333_5183 n1_521_5183 1.074286e+00
R2101 n1_521_5183 n1_2583_5183 1.178286e+01
R2102 n1_2583_5183 n1_2771_5183 1.074286e+00
R2103 n1_2771_5183 n1_4833_5183 1.178286e+01
R2104 n1_4833_5183 n1_5021_5183 1.074286e+00
R2105 n1_5021_5183 n1_7083_5183 1.178286e+01
R2106 n1_7083_5183 n1_7271_5183 1.074286e+00
R2107 n1_7271_5183 n1_9333_5183 1.178286e+01
R2108 n1_9333_5183 n1_9521_5183 1.074286e+00
R2109 n1_11583_5183 n1_11771_5183 1.074286e+00
R2110 n1_11771_5183 n1_13833_5183 1.178286e+01
R2111 n1_13833_5183 n1_14021_5183 1.074286e+00
R2112 n1_14021_5183 n1_16083_5183 1.178286e+01
R2113 n1_16083_5183 n1_16271_5183 1.074286e+00
R2114 n1_16271_5183 n1_18333_5183 1.178286e+01
R2115 n1_18333_5183 n1_18521_5183 1.074286e+00
R2116 n1_18521_5183 n1_20583_5183 1.178286e+01
R2117 n1_20583_5183 n1_20771_5183 1.074286e+00
R2118 n1_333_5216 n1_521_5216 1.074286e+00
R2119 n1_521_5216 n1_2583_5216 1.178286e+01
R2120 n1_2583_5216 n1_2771_5216 1.074286e+00
R2121 n1_2771_5216 n1_4833_5216 1.178286e+01
R2122 n1_4833_5216 n1_5021_5216 1.074286e+00
R2123 n1_5021_5216 n1_7083_5216 1.178286e+01
R2124 n1_7083_5216 n1_7271_5216 1.074286e+00
R2125 n1_7271_5216 n1_9333_5216 1.178286e+01
R2126 n1_9333_5216 n1_9521_5216 1.074286e+00
R2127 n1_11583_5216 n1_11771_5216 1.074286e+00
R2128 n1_11771_5216 n1_13833_5216 1.178286e+01
R2129 n1_13833_5216 n1_14021_5216 1.074286e+00
R2130 n1_14021_5216 n1_16083_5216 1.178286e+01
R2131 n1_16083_5216 n1_16271_5216 1.074286e+00
R2132 n1_16271_5216 n1_18333_5216 1.178286e+01
R2133 n1_18333_5216 n1_18521_5216 1.074286e+00
R2134 n1_18521_5216 n1_20583_5216 1.178286e+01
R2135 n1_20583_5216 n1_20771_5216 1.074286e+00
R2136 n1_333_5399 n1_521_5399 1.074286e+00
R2137 n1_521_5399 n1_2583_5399 1.178286e+01
R2138 n1_2583_5399 n1_2771_5399 1.074286e+00
R2139 n1_2771_5399 n1_4833_5399 1.178286e+01
R2140 n1_4833_5399 n1_5021_5399 1.074286e+00
R2141 n1_5021_5399 n1_7083_5399 1.178286e+01
R2142 n1_7083_5399 n1_7271_5399 1.074286e+00
R2143 n1_7271_5399 n1_9333_5399 1.178286e+01
R2144 n1_9333_5399 n1_9521_5399 1.074286e+00
R2145 n1_11583_5399 n1_11771_5399 1.074286e+00
R2146 n1_11771_5399 n1_13833_5399 1.178286e+01
R2147 n1_13833_5399 n1_14021_5399 1.074286e+00
R2148 n1_14021_5399 n1_16083_5399 1.178286e+01
R2149 n1_16083_5399 n1_16271_5399 1.074286e+00
R2150 n1_16271_5399 n1_18333_5399 1.178286e+01
R2151 n1_18333_5399 n1_18521_5399 1.074286e+00
R2152 n1_18521_5399 n1_20583_5399 1.178286e+01
R2153 n1_20583_5399 n1_20771_5399 1.074286e+00
R2154 n1_333_5432 n1_521_5432 1.074286e+00
R2155 n1_521_5432 n1_2583_5432 1.178286e+01
R2156 n1_2583_5432 n1_2771_5432 1.074286e+00
R2157 n1_2771_5432 n1_4833_5432 1.178286e+01
R2158 n1_4833_5432 n1_5021_5432 1.074286e+00
R2159 n1_5021_5432 n1_7083_5432 1.178286e+01
R2160 n1_7083_5432 n1_7271_5432 1.074286e+00
R2161 n1_7271_5432 n1_9333_5432 1.178286e+01
R2162 n1_9333_5432 n1_9521_5432 1.074286e+00
R2163 n1_11583_5432 n1_11771_5432 1.074286e+00
R2164 n1_11771_5432 n1_13833_5432 1.178286e+01
R2165 n1_13833_5432 n1_14021_5432 1.074286e+00
R2166 n1_14021_5432 n1_16083_5432 1.178286e+01
R2167 n1_16083_5432 n1_16271_5432 1.074286e+00
R2168 n1_16271_5432 n1_18333_5432 1.178286e+01
R2169 n1_18333_5432 n1_18521_5432 1.074286e+00
R2170 n1_18521_5432 n1_20583_5432 1.178286e+01
R2171 n1_20583_5432 n1_20771_5432 1.074286e+00
R2172 n1_333_5615 n1_521_5615 1.074286e+00
R2173 n1_521_5615 n1_2583_5615 1.178286e+01
R2174 n1_2583_5615 n1_2771_5615 1.074286e+00
R2175 n1_2771_5615 n1_4833_5615 1.178286e+01
R2176 n1_4833_5615 n1_5021_5615 1.074286e+00
R2177 n1_5021_5615 n1_7083_5615 1.178286e+01
R2178 n1_7083_5615 n1_7271_5615 1.074286e+00
R2179 n1_7271_5615 n1_9333_5615 1.178286e+01
R2180 n1_9333_5615 n1_9521_5615 1.074286e+00
R2181 n1_11583_5615 n1_11771_5615 1.074286e+00
R2182 n1_11771_5615 n1_13833_5615 1.178286e+01
R2183 n1_13833_5615 n1_14021_5615 1.074286e+00
R2184 n1_14021_5615 n1_16083_5615 1.178286e+01
R2185 n1_16083_5615 n1_16271_5615 1.074286e+00
R2186 n1_16271_5615 n1_18333_5615 1.178286e+01
R2187 n1_18333_5615 n1_18521_5615 1.074286e+00
R2188 n1_18521_5615 n1_20583_5615 1.178286e+01
R2189 n1_20583_5615 n1_20771_5615 1.074286e+00
R2190 n1_333_5648 n1_521_5648 1.074286e+00
R2191 n1_521_5648 n1_2583_5648 1.178286e+01
R2192 n1_2583_5648 n1_2771_5648 1.074286e+00
R2193 n1_2771_5648 n1_4833_5648 1.178286e+01
R2194 n1_4833_5648 n1_5021_5648 1.074286e+00
R2195 n1_5021_5648 n1_7083_5648 1.178286e+01
R2196 n1_7083_5648 n1_7271_5648 1.074286e+00
R2197 n1_7271_5648 n1_9333_5648 1.178286e+01
R2198 n1_9333_5648 n1_9521_5648 1.074286e+00
R2199 n1_11583_5648 n1_11771_5648 1.074286e+00
R2200 n1_11771_5648 n1_13833_5648 1.178286e+01
R2201 n1_13833_5648 n1_14021_5648 1.074286e+00
R2202 n1_14021_5648 n1_16083_5648 1.178286e+01
R2203 n1_16083_5648 n1_16271_5648 1.074286e+00
R2204 n1_16271_5648 n1_18333_5648 1.178286e+01
R2205 n1_18333_5648 n1_18521_5648 1.074286e+00
R2206 n1_18521_5648 n1_20583_5648 1.178286e+01
R2207 n1_20583_5648 n1_20771_5648 1.074286e+00
R2208 n1_333_5831 n1_521_5831 1.074286e+00
R2209 n1_521_5831 n1_2583_5831 1.178286e+01
R2210 n1_2583_5831 n1_2771_5831 1.074286e+00
R2211 n1_2771_5831 n1_4833_5831 1.178286e+01
R2212 n1_4833_5831 n1_5021_5831 1.074286e+00
R2213 n1_5021_5831 n1_7083_5831 1.178286e+01
R2214 n1_7083_5831 n1_7271_5831 1.074286e+00
R2215 n1_7271_5831 n1_9333_5831 1.178286e+01
R2216 n1_9333_5831 n1_9521_5831 1.074286e+00
R2217 n1_11583_5831 n1_11771_5831 1.074286e+00
R2218 n1_11771_5831 n1_13833_5831 1.178286e+01
R2219 n1_13833_5831 n1_14021_5831 1.074286e+00
R2220 n1_14021_5831 n1_16083_5831 1.178286e+01
R2221 n1_16083_5831 n1_16271_5831 1.074286e+00
R2222 n1_16271_5831 n1_18333_5831 1.178286e+01
R2223 n1_18333_5831 n1_18521_5831 1.074286e+00
R2224 n1_18521_5831 n1_20583_5831 1.178286e+01
R2225 n1_20583_5831 n1_20771_5831 1.074286e+00
R2226 n1_333_5864 n1_521_5864 1.074286e+00
R2227 n1_521_5864 n1_2583_5864 1.178286e+01
R2228 n1_2583_5864 n1_2771_5864 1.074286e+00
R2229 n1_2771_5864 n1_4833_5864 1.178286e+01
R2230 n1_4833_5864 n1_5021_5864 1.074286e+00
R2231 n1_5021_5864 n1_7083_5864 1.178286e+01
R2232 n1_7083_5864 n1_7271_5864 1.074286e+00
R2233 n1_7271_5864 n1_9333_5864 1.178286e+01
R2234 n1_9333_5864 n1_9521_5864 1.074286e+00
R2235 n1_11583_5864 n1_11771_5864 1.074286e+00
R2236 n1_11771_5864 n1_13833_5864 1.178286e+01
R2237 n1_13833_5864 n1_14021_5864 1.074286e+00
R2238 n1_14021_5864 n1_16083_5864 1.178286e+01
R2239 n1_16083_5864 n1_16271_5864 1.074286e+00
R2240 n1_16271_5864 n1_18333_5864 1.178286e+01
R2241 n1_18333_5864 n1_18521_5864 1.074286e+00
R2242 n1_18521_5864 n1_20583_5864 1.178286e+01
R2243 n1_20583_5864 n1_20771_5864 1.074286e+00
R2244 n1_521_6047 n1_2771_6047 1.285714e+01
R2245 n1_2771_6047 n1_5021_6047 1.285714e+01
R2246 n1_5021_6047 n1_7271_6047 1.285714e+01
R2247 n1_7271_6047 n1_9521_6047 1.285714e+01
R2248 n1_11771_6047 n1_14021_6047 1.285714e+01
R2249 n1_14021_6047 n1_16271_6047 1.285714e+01
R2250 n1_16271_6047 n1_18521_6047 1.285714e+01
R2251 n1_18521_6047 n1_20771_6047 1.285714e+01
R2252 n1_521_6080 n1_2771_6080 1.285714e+01
R2253 n1_2771_6080 n1_5021_6080 1.285714e+01
R2254 n1_5021_6080 n1_7271_6080 1.285714e+01
R2255 n1_7271_6080 n1_9521_6080 1.285714e+01
R2256 n1_11771_6080 n1_14021_6080 1.285714e+01
R2257 n1_14021_6080 n1_16271_6080 1.285714e+01
R2258 n1_16271_6080 n1_18521_6080 1.285714e+01
R2259 n1_18521_6080 n1_20771_6080 1.285714e+01
R2260 n1_333_6263 n1_521_6263 1.074286e+00
R2261 n1_521_6263 n1_2583_6263 1.178286e+01
R2262 n1_2583_6263 n1_2771_6263 1.074286e+00
R2263 n1_2771_6263 n1_4833_6263 1.178286e+01
R2264 n1_4833_6263 n1_5021_6263 1.074286e+00
R2265 n1_5021_6263 n1_7083_6263 1.178286e+01
R2266 n1_7083_6263 n1_7271_6263 1.074286e+00
R2267 n1_7271_6263 n1_9333_6263 1.178286e+01
R2268 n1_9333_6263 n1_9521_6263 1.074286e+00
R2269 n1_11583_6263 n1_11771_6263 1.074286e+00
R2270 n1_11771_6263 n1_13833_6263 1.178286e+01
R2271 n1_13833_6263 n1_14021_6263 1.074286e+00
R2272 n1_14021_6263 n1_16083_6263 1.178286e+01
R2273 n1_16083_6263 n1_16271_6263 1.074286e+00
R2274 n1_16271_6263 n1_18333_6263 1.178286e+01
R2275 n1_18333_6263 n1_18521_6263 1.074286e+00
R2276 n1_18521_6263 n1_20583_6263 1.178286e+01
R2277 n1_20583_6263 n1_20771_6263 1.074286e+00
R2278 n1_333_6296 n1_521_6296 1.074286e+00
R2279 n1_521_6296 n1_2583_6296 1.178286e+01
R2280 n1_2583_6296 n1_2771_6296 1.074286e+00
R2281 n1_2771_6296 n1_4833_6296 1.178286e+01
R2282 n1_4833_6296 n1_5021_6296 1.074286e+00
R2283 n1_5021_6296 n1_7083_6296 1.178286e+01
R2284 n1_7083_6296 n1_7271_6296 1.074286e+00
R2285 n1_7271_6296 n1_9333_6296 1.178286e+01
R2286 n1_9333_6296 n1_9521_6296 1.074286e+00
R2287 n1_11583_6296 n1_11771_6296 1.074286e+00
R2288 n1_11771_6296 n1_13833_6296 1.178286e+01
R2289 n1_13833_6296 n1_14021_6296 1.074286e+00
R2290 n1_14021_6296 n1_16083_6296 1.178286e+01
R2291 n1_16083_6296 n1_16271_6296 1.074286e+00
R2292 n1_16271_6296 n1_18333_6296 1.178286e+01
R2293 n1_18333_6296 n1_18521_6296 1.074286e+00
R2294 n1_18521_6296 n1_20583_6296 1.178286e+01
R2295 n1_20583_6296 n1_20771_6296 1.074286e+00
R2296 n1_333_6479 n1_521_6479 1.074286e+00
R2297 n1_521_6479 n1_2583_6479 1.178286e+01
R2298 n1_2583_6479 n1_2771_6479 1.074286e+00
R2299 n1_2771_6479 n1_4833_6479 1.178286e+01
R2300 n1_4833_6479 n1_5021_6479 1.074286e+00
R2301 n1_5021_6479 n1_7083_6479 1.178286e+01
R2302 n1_7083_6479 n1_7271_6479 1.074286e+00
R2303 n1_7271_6479 n1_9333_6479 1.178286e+01
R2304 n1_9333_6479 n1_9521_6479 1.074286e+00
R2305 n1_11583_6479 n1_11771_6479 1.074286e+00
R2306 n1_11771_6479 n1_13833_6479 1.178286e+01
R2307 n1_13833_6479 n1_14021_6479 1.074286e+00
R2308 n1_14021_6479 n1_16083_6479 1.178286e+01
R2309 n1_16083_6479 n1_16271_6479 1.074286e+00
R2310 n1_16271_6479 n1_18333_6479 1.178286e+01
R2311 n1_18333_6479 n1_18521_6479 1.074286e+00
R2312 n1_18521_6479 n1_20583_6479 1.178286e+01
R2313 n1_20583_6479 n1_20771_6479 1.074286e+00
R2314 n1_333_6512 n1_521_6512 1.074286e+00
R2315 n1_521_6512 n1_2583_6512 1.178286e+01
R2316 n1_2583_6512 n1_2771_6512 1.074286e+00
R2317 n1_2771_6512 n1_4833_6512 1.178286e+01
R2318 n1_4833_6512 n1_5021_6512 1.074286e+00
R2319 n1_5021_6512 n1_7083_6512 1.178286e+01
R2320 n1_7083_6512 n1_7271_6512 1.074286e+00
R2321 n1_7271_6512 n1_9333_6512 1.178286e+01
R2322 n1_9333_6512 n1_9521_6512 1.074286e+00
R2323 n1_11583_6512 n1_11771_6512 1.074286e+00
R2324 n1_11771_6512 n1_13833_6512 1.178286e+01
R2325 n1_13833_6512 n1_14021_6512 1.074286e+00
R2326 n1_14021_6512 n1_16083_6512 1.178286e+01
R2327 n1_16083_6512 n1_16271_6512 1.074286e+00
R2328 n1_16271_6512 n1_18333_6512 1.178286e+01
R2329 n1_18333_6512 n1_18521_6512 1.074286e+00
R2330 n1_18521_6512 n1_20583_6512 1.178286e+01
R2331 n1_20583_6512 n1_20771_6512 1.074286e+00
R2332 n1_333_6695 n1_521_6695 1.074286e+00
R2333 n1_521_6695 n1_2583_6695 1.178286e+01
R2334 n1_2583_6695 n1_2771_6695 1.074286e+00
R2335 n1_2771_6695 n1_4833_6695 1.178286e+01
R2336 n1_4833_6695 n1_5021_6695 1.074286e+00
R2337 n1_5021_6695 n1_7083_6695 1.178286e+01
R2338 n1_7083_6695 n1_7271_6695 1.074286e+00
R2339 n1_7271_6695 n1_9333_6695 1.178286e+01
R2340 n1_9333_6695 n1_9521_6695 1.074286e+00
R2341 n1_11583_6695 n1_11771_6695 1.074286e+00
R2342 n1_11771_6695 n1_13833_6695 1.178286e+01
R2343 n1_13833_6695 n1_14021_6695 1.074286e+00
R2344 n1_14021_6695 n1_16083_6695 1.178286e+01
R2345 n1_16083_6695 n1_16271_6695 1.074286e+00
R2346 n1_16271_6695 n1_18333_6695 1.178286e+01
R2347 n1_18333_6695 n1_18521_6695 1.074286e+00
R2348 n1_18521_6695 n1_20583_6695 1.178286e+01
R2349 n1_20583_6695 n1_20771_6695 1.074286e+00
R2350 n1_333_6728 n1_521_6728 1.074286e+00
R2351 n1_521_6728 n1_2583_6728 1.178286e+01
R2352 n1_2583_6728 n1_2771_6728 1.074286e+00
R2353 n1_2771_6728 n1_4833_6728 1.178286e+01
R2354 n1_4833_6728 n1_5021_6728 1.074286e+00
R2355 n1_5021_6728 n1_7083_6728 1.178286e+01
R2356 n1_7083_6728 n1_7271_6728 1.074286e+00
R2357 n1_7271_6728 n1_9333_6728 1.178286e+01
R2358 n1_9333_6728 n1_9521_6728 1.074286e+00
R2359 n1_11583_6728 n1_11771_6728 1.074286e+00
R2360 n1_11771_6728 n1_13833_6728 1.178286e+01
R2361 n1_13833_6728 n1_14021_6728 1.074286e+00
R2362 n1_14021_6728 n1_16083_6728 1.178286e+01
R2363 n1_16083_6728 n1_16271_6728 1.074286e+00
R2364 n1_16271_6728 n1_18333_6728 1.178286e+01
R2365 n1_18333_6728 n1_18521_6728 1.074286e+00
R2366 n1_18521_6728 n1_20583_6728 1.178286e+01
R2367 n1_20583_6728 n1_20771_6728 1.074286e+00
R2368 n1_333_6911 n1_521_6911 1.074286e+00
R2369 n1_521_6911 n1_2583_6911 1.178286e+01
R2370 n1_2583_6911 n1_2771_6911 1.074286e+00
R2371 n1_2771_6911 n1_4833_6911 1.178286e+01
R2372 n1_4833_6911 n1_5021_6911 1.074286e+00
R2373 n1_5021_6911 n1_7083_6911 1.178286e+01
R2374 n1_7083_6911 n1_7271_6911 1.074286e+00
R2375 n1_7271_6911 n1_9333_6911 1.178286e+01
R2376 n1_9333_6911 n1_9521_6911 1.074286e+00
R2377 n1_11583_6911 n1_11771_6911 1.074286e+00
R2378 n1_11771_6911 n1_13833_6911 1.178286e+01
R2379 n1_13833_6911 n1_14021_6911 1.074286e+00
R2380 n1_14021_6911 n1_16083_6911 1.178286e+01
R2381 n1_16083_6911 n1_16271_6911 1.074286e+00
R2382 n1_16271_6911 n1_18333_6911 1.178286e+01
R2383 n1_18333_6911 n1_18521_6911 1.074286e+00
R2384 n1_18521_6911 n1_20583_6911 1.178286e+01
R2385 n1_20583_6911 n1_20771_6911 1.074286e+00
R2386 n1_333_6944 n1_521_6944 1.074286e+00
R2387 n1_521_6944 n1_2583_6944 1.178286e+01
R2388 n1_2583_6944 n1_2771_6944 1.074286e+00
R2389 n1_2771_6944 n1_4833_6944 1.178286e+01
R2390 n1_4833_6944 n1_5021_6944 1.074286e+00
R2391 n1_5021_6944 n1_7083_6944 1.178286e+01
R2392 n1_7083_6944 n1_7271_6944 1.074286e+00
R2393 n1_7271_6944 n1_9333_6944 1.178286e+01
R2394 n1_9333_6944 n1_9521_6944 1.074286e+00
R2395 n1_11583_6944 n1_11771_6944 1.074286e+00
R2396 n1_11771_6944 n1_13833_6944 1.178286e+01
R2397 n1_13833_6944 n1_14021_6944 1.074286e+00
R2398 n1_14021_6944 n1_16083_6944 1.178286e+01
R2399 n1_16083_6944 n1_16271_6944 1.074286e+00
R2400 n1_16271_6944 n1_18333_6944 1.178286e+01
R2401 n1_18333_6944 n1_18521_6944 1.074286e+00
R2402 n1_18521_6944 n1_20583_6944 1.178286e+01
R2403 n1_20583_6944 n1_20771_6944 1.074286e+00
R2404 n1_333_7127 n1_521_7127 1.074286e+00
R2405 n1_521_7127 n1_2583_7127 1.178286e+01
R2406 n1_2583_7127 n1_2771_7127 1.074286e+00
R2407 n1_2771_7127 n1_4833_7127 1.178286e+01
R2408 n1_4833_7127 n1_5021_7127 1.074286e+00
R2409 n1_5021_7127 n1_7083_7127 1.178286e+01
R2410 n1_7083_7127 n1_7271_7127 1.074286e+00
R2411 n1_7271_7127 n1_9333_7127 1.178286e+01
R2412 n1_9333_7127 n1_9521_7127 1.074286e+00
R2413 n1_11583_7127 n1_11771_7127 1.074286e+00
R2414 n1_11771_7127 n1_13833_7127 1.178286e+01
R2415 n1_13833_7127 n1_14021_7127 1.074286e+00
R2416 n1_14021_7127 n1_16083_7127 1.178286e+01
R2417 n1_16083_7127 n1_16271_7127 1.074286e+00
R2418 n1_16271_7127 n1_18333_7127 1.178286e+01
R2419 n1_18333_7127 n1_18521_7127 1.074286e+00
R2420 n1_18521_7127 n1_20583_7127 1.178286e+01
R2421 n1_20583_7127 n1_20771_7127 1.074286e+00
R2422 n1_333_7160 n1_380_7160 2.685714e-01
R2423 n1_380_7160 n1_521_7160 8.057143e-01
R2424 n1_521_7160 n1_2583_7160 1.178286e+01
R2425 n1_2583_7160 n1_2630_7160 2.685714e-01
R2426 n1_2630_7160 n1_2771_7160 8.057143e-01
R2427 n1_2771_7160 n1_4833_7160 1.178286e+01
R2428 n1_4833_7160 n1_4880_7160 2.685714e-01
R2429 n1_4880_7160 n1_5021_7160 8.057143e-01
R2430 n1_5021_7160 n1_7083_7160 1.178286e+01
R2431 n1_7083_7160 n1_7130_7160 2.685714e-01
R2432 n1_7130_7160 n1_7271_7160 8.057143e-01
R2433 n1_7271_7160 n1_9333_7160 1.178286e+01
R2434 n1_9333_7160 n1_9380_7160 2.685714e-01
R2435 n1_9380_7160 n1_9521_7160 8.057143e-01
R2436 n1_11583_7160 n1_11630_7160 2.685714e-01
R2437 n1_11630_7160 n1_11771_7160 8.057143e-01
R2438 n1_11771_7160 n1_13833_7160 1.178286e+01
R2439 n1_13833_7160 n1_13880_7160 2.685714e-01
R2440 n1_13880_7160 n1_14021_7160 8.057143e-01
R2441 n1_14021_7160 n1_16083_7160 1.178286e+01
R2442 n1_16083_7160 n1_16130_7160 2.685714e-01
R2443 n1_16130_7160 n1_16271_7160 8.057143e-01
R2444 n1_16271_7160 n1_18333_7160 1.178286e+01
R2445 n1_18333_7160 n1_18380_7160 2.685714e-01
R2446 n1_18380_7160 n1_18521_7160 8.057143e-01
R2447 n1_18521_7160 n1_20583_7160 1.178286e+01
R2448 n1_20583_7160 n1_20630_7160 2.685714e-01
R2449 n1_20630_7160 n1_20771_7160 8.057143e-01
R2450 n1_333_7343 n1_521_7343 1.074286e+00
R2451 n1_521_7343 n1_2583_7343 1.178286e+01
R2452 n1_2583_7343 n1_2771_7343 1.074286e+00
R2453 n1_2771_7343 n1_4833_7343 1.178286e+01
R2454 n1_4833_7343 n1_5021_7343 1.074286e+00
R2455 n1_5021_7343 n1_7083_7343 1.178286e+01
R2456 n1_7083_7343 n1_7271_7343 1.074286e+00
R2457 n1_7271_7343 n1_9333_7343 1.178286e+01
R2458 n1_9333_7343 n1_9521_7343 1.074286e+00
R2459 n1_11583_7343 n1_11771_7343 1.074286e+00
R2460 n1_11771_7343 n1_13833_7343 1.178286e+01
R2461 n1_13833_7343 n1_14021_7343 1.074286e+00
R2462 n1_14021_7343 n1_16083_7343 1.178286e+01
R2463 n1_16083_7343 n1_16271_7343 1.074286e+00
R2464 n1_16271_7343 n1_18333_7343 1.178286e+01
R2465 n1_18333_7343 n1_18521_7343 1.074286e+00
R2466 n1_18521_7343 n1_20583_7343 1.178286e+01
R2467 n1_20583_7343 n1_20771_7343 1.074286e+00
R2468 n1_333_7376 n1_521_7376 1.074286e+00
R2469 n1_521_7376 n1_2583_7376 1.178286e+01
R2470 n1_2583_7376 n1_2771_7376 1.074286e+00
R2471 n1_2771_7376 n1_4833_7376 1.178286e+01
R2472 n1_4833_7376 n1_5021_7376 1.074286e+00
R2473 n1_5021_7376 n1_7083_7376 1.178286e+01
R2474 n1_7083_7376 n1_7271_7376 1.074286e+00
R2475 n1_7271_7376 n1_9333_7376 1.178286e+01
R2476 n1_9333_7376 n1_9521_7376 1.074286e+00
R2477 n1_11583_7376 n1_11771_7376 1.074286e+00
R2478 n1_11771_7376 n1_13833_7376 1.178286e+01
R2479 n1_13833_7376 n1_14021_7376 1.074286e+00
R2480 n1_14021_7376 n1_16083_7376 1.178286e+01
R2481 n1_16083_7376 n1_16271_7376 1.074286e+00
R2482 n1_16271_7376 n1_18333_7376 1.178286e+01
R2483 n1_18333_7376 n1_18521_7376 1.074286e+00
R2484 n1_18521_7376 n1_20583_7376 1.178286e+01
R2485 n1_20583_7376 n1_20771_7376 1.074286e+00
R2486 n1_333_7559 n1_521_7559 1.074286e+00
R2487 n1_521_7559 n1_2583_7559 1.178286e+01
R2488 n1_2583_7559 n1_2771_7559 1.074286e+00
R2489 n1_2771_7559 n1_4833_7559 1.178286e+01
R2490 n1_4833_7559 n1_5021_7559 1.074286e+00
R2491 n1_5021_7559 n1_7083_7559 1.178286e+01
R2492 n1_7083_7559 n1_7271_7559 1.074286e+00
R2493 n1_7271_7559 n1_9333_7559 1.178286e+01
R2494 n1_9333_7559 n1_9521_7559 1.074286e+00
R2495 n1_11583_7559 n1_11771_7559 1.074286e+00
R2496 n1_11771_7559 n1_13833_7559 1.178286e+01
R2497 n1_13833_7559 n1_14021_7559 1.074286e+00
R2498 n1_14021_7559 n1_16083_7559 1.178286e+01
R2499 n1_16083_7559 n1_16271_7559 1.074286e+00
R2500 n1_16271_7559 n1_18333_7559 1.178286e+01
R2501 n1_18333_7559 n1_18521_7559 1.074286e+00
R2502 n1_18521_7559 n1_20583_7559 1.178286e+01
R2503 n1_20583_7559 n1_20771_7559 1.074286e+00
R2504 n1_333_7592 n1_521_7592 1.074286e+00
R2505 n1_521_7592 n1_2583_7592 1.178286e+01
R2506 n1_2583_7592 n1_2771_7592 1.074286e+00
R2507 n1_2771_7592 n1_4833_7592 1.178286e+01
R2508 n1_4833_7592 n1_5021_7592 1.074286e+00
R2509 n1_5021_7592 n1_7083_7592 1.178286e+01
R2510 n1_7083_7592 n1_7271_7592 1.074286e+00
R2511 n1_7271_7592 n1_9333_7592 1.178286e+01
R2512 n1_9333_7592 n1_9521_7592 1.074286e+00
R2513 n1_11583_7592 n1_11771_7592 1.074286e+00
R2514 n1_11771_7592 n1_13833_7592 1.178286e+01
R2515 n1_13833_7592 n1_14021_7592 1.074286e+00
R2516 n1_14021_7592 n1_16083_7592 1.178286e+01
R2517 n1_16083_7592 n1_16271_7592 1.074286e+00
R2518 n1_16271_7592 n1_18333_7592 1.178286e+01
R2519 n1_18333_7592 n1_18521_7592 1.074286e+00
R2520 n1_18521_7592 n1_20583_7592 1.178286e+01
R2521 n1_20583_7592 n1_20771_7592 1.074286e+00
R2522 n1_333_7775 n1_521_7775 1.074286e+00
R2523 n1_521_7775 n1_2583_7775 1.178286e+01
R2524 n1_2583_7775 n1_2771_7775 1.074286e+00
R2525 n1_2771_7775 n1_4833_7775 1.178286e+01
R2526 n1_4833_7775 n1_5021_7775 1.074286e+00
R2527 n1_5021_7775 n1_7083_7775 1.178286e+01
R2528 n1_7083_7775 n1_7271_7775 1.074286e+00
R2529 n1_7271_7775 n1_9333_7775 1.178286e+01
R2530 n1_9333_7775 n1_9521_7775 1.074286e+00
R2531 n1_11583_7775 n1_11771_7775 1.074286e+00
R2532 n1_11771_7775 n1_13833_7775 1.178286e+01
R2533 n1_13833_7775 n1_14021_7775 1.074286e+00
R2534 n1_14021_7775 n1_16083_7775 1.178286e+01
R2535 n1_16083_7775 n1_16271_7775 1.074286e+00
R2536 n1_16271_7775 n1_18333_7775 1.178286e+01
R2537 n1_18333_7775 n1_18521_7775 1.074286e+00
R2538 n1_18521_7775 n1_20583_7775 1.178286e+01
R2539 n1_20583_7775 n1_20771_7775 1.074286e+00
R2540 n1_333_7808 n1_521_7808 1.074286e+00
R2541 n1_521_7808 n1_2583_7808 1.178286e+01
R2542 n1_2583_7808 n1_2771_7808 1.074286e+00
R2543 n1_2771_7808 n1_4833_7808 1.178286e+01
R2544 n1_4833_7808 n1_5021_7808 1.074286e+00
R2545 n1_5021_7808 n1_7083_7808 1.178286e+01
R2546 n1_7083_7808 n1_7271_7808 1.074286e+00
R2547 n1_7271_7808 n1_9333_7808 1.178286e+01
R2548 n1_9333_7808 n1_9521_7808 1.074286e+00
R2549 n1_11583_7808 n1_11771_7808 1.074286e+00
R2550 n1_11771_7808 n1_13833_7808 1.178286e+01
R2551 n1_13833_7808 n1_14021_7808 1.074286e+00
R2552 n1_14021_7808 n1_16083_7808 1.178286e+01
R2553 n1_16083_7808 n1_16271_7808 1.074286e+00
R2554 n1_16271_7808 n1_18333_7808 1.178286e+01
R2555 n1_18333_7808 n1_18521_7808 1.074286e+00
R2556 n1_18521_7808 n1_20583_7808 1.178286e+01
R2557 n1_20583_7808 n1_20771_7808 1.074286e+00
R2558 n1_333_7991 n1_521_7991 1.074286e+00
R2559 n1_521_7991 n1_2583_7991 1.178286e+01
R2560 n1_2583_7991 n1_2771_7991 1.074286e+00
R2561 n1_2771_7991 n1_4833_7991 1.178286e+01
R2562 n1_4833_7991 n1_5021_7991 1.074286e+00
R2563 n1_5021_7991 n1_7083_7991 1.178286e+01
R2564 n1_7083_7991 n1_7271_7991 1.074286e+00
R2565 n1_7271_7991 n1_9333_7991 1.178286e+01
R2566 n1_9333_7991 n1_9521_7991 1.074286e+00
R2567 n1_11583_7991 n1_11771_7991 1.074286e+00
R2568 n1_11771_7991 n1_13833_7991 1.178286e+01
R2569 n1_13833_7991 n1_14021_7991 1.074286e+00
R2570 n1_14021_7991 n1_16083_7991 1.178286e+01
R2571 n1_16083_7991 n1_16271_7991 1.074286e+00
R2572 n1_16271_7991 n1_18333_7991 1.178286e+01
R2573 n1_18333_7991 n1_18521_7991 1.074286e+00
R2574 n1_18521_7991 n1_20583_7991 1.178286e+01
R2575 n1_20583_7991 n1_20771_7991 1.074286e+00
R2576 n1_333_8024 n1_521_8024 1.074286e+00
R2577 n1_521_8024 n1_2583_8024 1.178286e+01
R2578 n1_2583_8024 n1_2771_8024 1.074286e+00
R2579 n1_2771_8024 n1_4833_8024 1.178286e+01
R2580 n1_4833_8024 n1_5021_8024 1.074286e+00
R2581 n1_5021_8024 n1_7083_8024 1.178286e+01
R2582 n1_7083_8024 n1_7271_8024 1.074286e+00
R2583 n1_7271_8024 n1_9333_8024 1.178286e+01
R2584 n1_9333_8024 n1_9521_8024 1.074286e+00
R2585 n1_11583_8024 n1_11771_8024 1.074286e+00
R2586 n1_11771_8024 n1_13833_8024 1.178286e+01
R2587 n1_13833_8024 n1_14021_8024 1.074286e+00
R2588 n1_14021_8024 n1_16083_8024 1.178286e+01
R2589 n1_16083_8024 n1_16271_8024 1.074286e+00
R2590 n1_16271_8024 n1_18333_8024 1.178286e+01
R2591 n1_18333_8024 n1_18521_8024 1.074286e+00
R2592 n1_18521_8024 n1_20583_8024 1.178286e+01
R2593 n1_20583_8024 n1_20771_8024 1.074286e+00
R2594 n1_333_8207 n1_521_8207 1.074286e+00
R2595 n1_521_8207 n1_2583_8207 1.178286e+01
R2596 n1_2583_8207 n1_2771_8207 1.074286e+00
R2597 n1_2771_8207 n1_4833_8207 1.178286e+01
R2598 n1_4833_8207 n1_5021_8207 1.074286e+00
R2599 n1_5021_8207 n1_7083_8207 1.178286e+01
R2600 n1_7083_8207 n1_7271_8207 1.074286e+00
R2601 n1_7271_8207 n1_9333_8207 1.178286e+01
R2602 n1_9333_8207 n1_9521_8207 1.074286e+00
R2603 n1_11583_8207 n1_11771_8207 1.074286e+00
R2604 n1_11771_8207 n1_13833_8207 1.178286e+01
R2605 n1_13833_8207 n1_14021_8207 1.074286e+00
R2606 n1_14021_8207 n1_16083_8207 1.178286e+01
R2607 n1_16083_8207 n1_16271_8207 1.074286e+00
R2608 n1_16271_8207 n1_18333_8207 1.178286e+01
R2609 n1_18333_8207 n1_18521_8207 1.074286e+00
R2610 n1_18521_8207 n1_20583_8207 1.178286e+01
R2611 n1_20583_8207 n1_20771_8207 1.074286e+00
R2612 n1_333_8240 n1_521_8240 1.074286e+00
R2613 n1_521_8240 n1_2583_8240 1.178286e+01
R2614 n1_2583_8240 n1_2771_8240 1.074286e+00
R2615 n1_2771_8240 n1_4833_8240 1.178286e+01
R2616 n1_4833_8240 n1_5021_8240 1.074286e+00
R2617 n1_5021_8240 n1_7083_8240 1.178286e+01
R2618 n1_7083_8240 n1_7271_8240 1.074286e+00
R2619 n1_7271_8240 n1_9333_8240 1.178286e+01
R2620 n1_9333_8240 n1_9521_8240 1.074286e+00
R2621 n1_11583_8240 n1_11771_8240 1.074286e+00
R2622 n1_11771_8240 n1_13833_8240 1.178286e+01
R2623 n1_13833_8240 n1_14021_8240 1.074286e+00
R2624 n1_14021_8240 n1_16083_8240 1.178286e+01
R2625 n1_16083_8240 n1_16271_8240 1.074286e+00
R2626 n1_16271_8240 n1_18333_8240 1.178286e+01
R2627 n1_18333_8240 n1_18521_8240 1.074286e+00
R2628 n1_18521_8240 n1_20583_8240 1.178286e+01
R2629 n1_20583_8240 n1_20771_8240 1.074286e+00
R2630 n1_521_8423 n1_2771_8423 1.285714e+01
R2631 n1_2771_8423 n1_5021_8423 1.285714e+01
R2632 n1_5021_8423 n1_7271_8423 1.285714e+01
R2633 n1_7271_8423 n1_9521_8423 1.285714e+01
R2634 n1_11771_8423 n1_14021_8423 1.285714e+01
R2635 n1_14021_8423 n1_16271_8423 1.285714e+01
R2636 n1_16271_8423 n1_18521_8423 1.285714e+01
R2637 n1_18521_8423 n1_20771_8423 1.285714e+01
R2638 n1_333_8456 n1_521_8456 1.074286e+00
R2639 n1_521_8456 n1_2583_8456 1.178286e+01
R2640 n1_2583_8456 n1_2771_8456 1.074286e+00
R2641 n1_2771_8456 n1_4833_8456 1.178286e+01
R2642 n1_4833_8456 n1_5021_8456 1.074286e+00
R2643 n1_5021_8456 n1_7083_8456 1.178286e+01
R2644 n1_7083_8456 n1_7271_8456 1.074286e+00
R2645 n1_7271_8456 n1_9333_8456 1.178286e+01
R2646 n1_9333_8456 n1_9521_8456 1.074286e+00
R2647 n1_11583_8456 n1_11771_8456 1.074286e+00
R2648 n1_11771_8456 n1_13833_8456 1.178286e+01
R2649 n1_13833_8456 n1_14021_8456 1.074286e+00
R2650 n1_14021_8456 n1_16083_8456 1.178286e+01
R2651 n1_16083_8456 n1_16271_8456 1.074286e+00
R2652 n1_16271_8456 n1_18333_8456 1.178286e+01
R2653 n1_18333_8456 n1_18521_8456 1.074286e+00
R2654 n1_18521_8456 n1_20583_8456 1.178286e+01
R2655 n1_20583_8456 n1_20771_8456 1.074286e+00
R2656 n1_333_8639 n1_521_8639 1.074286e+00
R2657 n1_521_8639 n1_2583_8639 1.178286e+01
R2658 n1_2583_8639 n1_2771_8639 1.074286e+00
R2659 n1_2771_8639 n1_4833_8639 1.178286e+01
R2660 n1_4833_8639 n1_5021_8639 1.074286e+00
R2661 n1_5021_8639 n1_7083_8639 1.178286e+01
R2662 n1_7083_8639 n1_7271_8639 1.074286e+00
R2663 n1_7271_8639 n1_9333_8639 1.178286e+01
R2664 n1_9333_8639 n1_9521_8639 1.074286e+00
R2665 n1_11583_8639 n1_11771_8639 1.074286e+00
R2666 n1_11771_8639 n1_13833_8639 1.178286e+01
R2667 n1_13833_8639 n1_14021_8639 1.074286e+00
R2668 n1_14021_8639 n1_16083_8639 1.178286e+01
R2669 n1_16083_8639 n1_16271_8639 1.074286e+00
R2670 n1_16271_8639 n1_18333_8639 1.178286e+01
R2671 n1_18333_8639 n1_18521_8639 1.074286e+00
R2672 n1_18521_8639 n1_20583_8639 1.178286e+01
R2673 n1_20583_8639 n1_20771_8639 1.074286e+00
R2674 n1_333_8672 n1_521_8672 1.074286e+00
R2675 n1_521_8672 n1_2583_8672 1.178286e+01
R2676 n1_2583_8672 n1_2771_8672 1.074286e+00
R2677 n1_2771_8672 n1_4833_8672 1.178286e+01
R2678 n1_4833_8672 n1_5021_8672 1.074286e+00
R2679 n1_5021_8672 n1_7083_8672 1.178286e+01
R2680 n1_7083_8672 n1_7271_8672 1.074286e+00
R2681 n1_7271_8672 n1_9333_8672 1.178286e+01
R2682 n1_9333_8672 n1_9521_8672 1.074286e+00
R2683 n1_11583_8672 n1_11771_8672 1.074286e+00
R2684 n1_11771_8672 n1_13833_8672 1.178286e+01
R2685 n1_13833_8672 n1_14021_8672 1.074286e+00
R2686 n1_14021_8672 n1_16083_8672 1.178286e+01
R2687 n1_16083_8672 n1_16271_8672 1.074286e+00
R2688 n1_16271_8672 n1_18333_8672 1.178286e+01
R2689 n1_18333_8672 n1_18521_8672 1.074286e+00
R2690 n1_18521_8672 n1_20583_8672 1.178286e+01
R2691 n1_20583_8672 n1_20771_8672 1.074286e+00
R2692 n1_333_8855 n1_521_8855 1.074286e+00
R2693 n1_521_8855 n1_2583_8855 1.178286e+01
R2694 n1_2583_8855 n1_2771_8855 1.074286e+00
R2695 n1_2771_8855 n1_4833_8855 1.178286e+01
R2696 n1_4833_8855 n1_5021_8855 1.074286e+00
R2697 n1_5021_8855 n1_7083_8855 1.178286e+01
R2698 n1_7083_8855 n1_7271_8855 1.074286e+00
R2699 n1_7271_8855 n1_9333_8855 1.178286e+01
R2700 n1_9333_8855 n1_9521_8855 1.074286e+00
R2701 n1_11583_8855 n1_11771_8855 1.074286e+00
R2702 n1_11771_8855 n1_13833_8855 1.178286e+01
R2703 n1_13833_8855 n1_14021_8855 1.074286e+00
R2704 n1_14021_8855 n1_16083_8855 1.178286e+01
R2705 n1_16083_8855 n1_16271_8855 1.074286e+00
R2706 n1_16271_8855 n1_18333_8855 1.178286e+01
R2707 n1_18333_8855 n1_18521_8855 1.074286e+00
R2708 n1_18521_8855 n1_20583_8855 1.178286e+01
R2709 n1_20583_8855 n1_20771_8855 1.074286e+00
R2710 n1_333_8888 n1_521_8888 1.074286e+00
R2711 n1_521_8888 n1_2583_8888 1.178286e+01
R2712 n1_2583_8888 n1_2771_8888 1.074286e+00
R2713 n1_2771_8888 n1_4833_8888 1.178286e+01
R2714 n1_4833_8888 n1_5021_8888 1.074286e+00
R2715 n1_5021_8888 n1_7083_8888 1.178286e+01
R2716 n1_7083_8888 n1_7271_8888 1.074286e+00
R2717 n1_7271_8888 n1_9333_8888 1.178286e+01
R2718 n1_9333_8888 n1_9521_8888 1.074286e+00
R2719 n1_11583_8888 n1_11771_8888 1.074286e+00
R2720 n1_11771_8888 n1_13833_8888 1.178286e+01
R2721 n1_13833_8888 n1_14021_8888 1.074286e+00
R2722 n1_14021_8888 n1_16083_8888 1.178286e+01
R2723 n1_16083_8888 n1_16271_8888 1.074286e+00
R2724 n1_16271_8888 n1_18333_8888 1.178286e+01
R2725 n1_18333_8888 n1_18521_8888 1.074286e+00
R2726 n1_18521_8888 n1_20583_8888 1.178286e+01
R2727 n1_20583_8888 n1_20771_8888 1.074286e+00
R2728 n1_333_9071 n1_521_9071 1.074286e+00
R2729 n1_521_9071 n1_2583_9071 1.178286e+01
R2730 n1_2583_9071 n1_2771_9071 1.074286e+00
R2731 n1_2771_9071 n1_4833_9071 1.178286e+01
R2732 n1_4833_9071 n1_5021_9071 1.074286e+00
R2733 n1_5021_9071 n1_7083_9071 1.178286e+01
R2734 n1_7083_9071 n1_7271_9071 1.074286e+00
R2735 n1_7271_9071 n1_9333_9071 1.178286e+01
R2736 n1_9333_9071 n1_9521_9071 1.074286e+00
R2737 n1_11583_9071 n1_11771_9071 1.074286e+00
R2738 n1_11771_9071 n1_13833_9071 1.178286e+01
R2739 n1_13833_9071 n1_14021_9071 1.074286e+00
R2740 n1_14021_9071 n1_16083_9071 1.178286e+01
R2741 n1_16083_9071 n1_16271_9071 1.074286e+00
R2742 n1_16271_9071 n1_18333_9071 1.178286e+01
R2743 n1_18333_9071 n1_18521_9071 1.074286e+00
R2744 n1_18521_9071 n1_20583_9071 1.178286e+01
R2745 n1_20583_9071 n1_20771_9071 1.074286e+00
R2746 n1_333_9104 n1_521_9104 1.074286e+00
R2747 n1_521_9104 n1_2583_9104 1.178286e+01
R2748 n1_2583_9104 n1_2771_9104 1.074286e+00
R2749 n1_2771_9104 n1_4833_9104 1.178286e+01
R2750 n1_4833_9104 n1_5021_9104 1.074286e+00
R2751 n1_5021_9104 n1_7083_9104 1.178286e+01
R2752 n1_7083_9104 n1_7271_9104 1.074286e+00
R2753 n1_7271_9104 n1_9333_9104 1.178286e+01
R2754 n1_9333_9104 n1_9521_9104 1.074286e+00
R2755 n1_11583_9104 n1_11771_9104 1.074286e+00
R2756 n1_11771_9104 n1_13833_9104 1.178286e+01
R2757 n1_13833_9104 n1_14021_9104 1.074286e+00
R2758 n1_14021_9104 n1_16083_9104 1.178286e+01
R2759 n1_16083_9104 n1_16271_9104 1.074286e+00
R2760 n1_16271_9104 n1_18333_9104 1.178286e+01
R2761 n1_18333_9104 n1_18521_9104 1.074286e+00
R2762 n1_18521_9104 n1_20583_9104 1.178286e+01
R2763 n1_20583_9104 n1_20771_9104 1.074286e+00
R2764 n1_333_12095 n1_521_12095 1.074286e+00
R2765 n1_521_12095 n1_2583_12095 1.178286e+01
R2766 n1_2583_12095 n1_2771_12095 1.074286e+00
R2767 n1_2771_12095 n1_4833_12095 1.178286e+01
R2768 n1_4833_12095 n1_5021_12095 1.074286e+00
R2769 n1_5021_12095 n1_7083_12095 1.178286e+01
R2770 n1_7083_12095 n1_7271_12095 1.074286e+00
R2771 n1_7271_12095 n1_9333_12095 1.178286e+01
R2772 n1_9333_12095 n1_9521_12095 1.074286e+00
R2773 n1_11583_12095 n1_11771_12095 1.074286e+00
R2774 n1_11771_12095 n1_13833_12095 1.178286e+01
R2775 n1_13833_12095 n1_14021_12095 1.074286e+00
R2776 n1_14021_12095 n1_16083_12095 1.178286e+01
R2777 n1_16083_12095 n1_16271_12095 1.074286e+00
R2778 n1_16271_12095 n1_18333_12095 1.178286e+01
R2779 n1_18333_12095 n1_18521_12095 1.074286e+00
R2780 n1_18521_12095 n1_20583_12095 1.178286e+01
R2781 n1_20583_12095 n1_20771_12095 1.074286e+00
R2782 n1_333_12128 n1_521_12128 1.074286e+00
R2783 n1_521_12128 n1_2583_12128 1.178286e+01
R2784 n1_2583_12128 n1_2771_12128 1.074286e+00
R2785 n1_2771_12128 n1_4833_12128 1.178286e+01
R2786 n1_4833_12128 n1_5021_12128 1.074286e+00
R2787 n1_5021_12128 n1_7083_12128 1.178286e+01
R2788 n1_7083_12128 n1_7271_12128 1.074286e+00
R2789 n1_7271_12128 n1_9333_12128 1.178286e+01
R2790 n1_9333_12128 n1_9521_12128 1.074286e+00
R2791 n1_11583_12128 n1_11771_12128 1.074286e+00
R2792 n1_11771_12128 n1_13833_12128 1.178286e+01
R2793 n1_13833_12128 n1_14021_12128 1.074286e+00
R2794 n1_14021_12128 n1_16083_12128 1.178286e+01
R2795 n1_16083_12128 n1_16271_12128 1.074286e+00
R2796 n1_16271_12128 n1_18333_12128 1.178286e+01
R2797 n1_18333_12128 n1_18521_12128 1.074286e+00
R2798 n1_18521_12128 n1_20583_12128 1.178286e+01
R2799 n1_20583_12128 n1_20771_12128 1.074286e+00
R2800 n1_333_12311 n1_521_12311 1.074286e+00
R2801 n1_521_12311 n1_2583_12311 1.178286e+01
R2802 n1_2583_12311 n1_2771_12311 1.074286e+00
R2803 n1_2771_12311 n1_4833_12311 1.178286e+01
R2804 n1_4833_12311 n1_5021_12311 1.074286e+00
R2805 n1_5021_12311 n1_7083_12311 1.178286e+01
R2806 n1_7083_12311 n1_7271_12311 1.074286e+00
R2807 n1_7271_12311 n1_9333_12311 1.178286e+01
R2808 n1_9333_12311 n1_9521_12311 1.074286e+00
R2809 n1_11583_12311 n1_11771_12311 1.074286e+00
R2810 n1_11771_12311 n1_13833_12311 1.178286e+01
R2811 n1_13833_12311 n1_14021_12311 1.074286e+00
R2812 n1_14021_12311 n1_16083_12311 1.178286e+01
R2813 n1_16083_12311 n1_16271_12311 1.074286e+00
R2814 n1_16271_12311 n1_18333_12311 1.178286e+01
R2815 n1_18333_12311 n1_18521_12311 1.074286e+00
R2816 n1_18521_12311 n1_20583_12311 1.178286e+01
R2817 n1_20583_12311 n1_20771_12311 1.074286e+00
R2818 n1_333_12344 n1_521_12344 1.074286e+00
R2819 n1_521_12344 n1_2583_12344 1.178286e+01
R2820 n1_2583_12344 n1_2771_12344 1.074286e+00
R2821 n1_2771_12344 n1_4833_12344 1.178286e+01
R2822 n1_4833_12344 n1_5021_12344 1.074286e+00
R2823 n1_5021_12344 n1_7083_12344 1.178286e+01
R2824 n1_7083_12344 n1_7271_12344 1.074286e+00
R2825 n1_7271_12344 n1_9333_12344 1.178286e+01
R2826 n1_9333_12344 n1_9521_12344 1.074286e+00
R2827 n1_11583_12344 n1_11771_12344 1.074286e+00
R2828 n1_11771_12344 n1_13833_12344 1.178286e+01
R2829 n1_13833_12344 n1_14021_12344 1.074286e+00
R2830 n1_14021_12344 n1_16083_12344 1.178286e+01
R2831 n1_16083_12344 n1_16271_12344 1.074286e+00
R2832 n1_16271_12344 n1_18333_12344 1.178286e+01
R2833 n1_18333_12344 n1_18521_12344 1.074286e+00
R2834 n1_18521_12344 n1_20583_12344 1.178286e+01
R2835 n1_20583_12344 n1_20771_12344 1.074286e+00
R2836 n1_333_12527 n1_521_12527 1.074286e+00
R2837 n1_521_12527 n1_2583_12527 1.178286e+01
R2838 n1_2583_12527 n1_2771_12527 1.074286e+00
R2839 n1_2771_12527 n1_4833_12527 1.178286e+01
R2840 n1_4833_12527 n1_5021_12527 1.074286e+00
R2841 n1_5021_12527 n1_7083_12527 1.178286e+01
R2842 n1_7083_12527 n1_7271_12527 1.074286e+00
R2843 n1_7271_12527 n1_9333_12527 1.178286e+01
R2844 n1_9333_12527 n1_9521_12527 1.074286e+00
R2845 n1_11583_12527 n1_11771_12527 1.074286e+00
R2846 n1_11771_12527 n1_13833_12527 1.178286e+01
R2847 n1_13833_12527 n1_14021_12527 1.074286e+00
R2848 n1_14021_12527 n1_16083_12527 1.178286e+01
R2849 n1_16083_12527 n1_16271_12527 1.074286e+00
R2850 n1_16271_12527 n1_18333_12527 1.178286e+01
R2851 n1_18333_12527 n1_18521_12527 1.074286e+00
R2852 n1_18521_12527 n1_20583_12527 1.178286e+01
R2853 n1_20583_12527 n1_20771_12527 1.074286e+00
R2854 n1_333_12560 n1_521_12560 1.074286e+00
R2855 n1_521_12560 n1_2583_12560 1.178286e+01
R2856 n1_2583_12560 n1_2771_12560 1.074286e+00
R2857 n1_2771_12560 n1_4833_12560 1.178286e+01
R2858 n1_4833_12560 n1_5021_12560 1.074286e+00
R2859 n1_5021_12560 n1_7083_12560 1.178286e+01
R2860 n1_7083_12560 n1_7271_12560 1.074286e+00
R2861 n1_7271_12560 n1_9333_12560 1.178286e+01
R2862 n1_9333_12560 n1_9521_12560 1.074286e+00
R2863 n1_11583_12560 n1_11771_12560 1.074286e+00
R2864 n1_11771_12560 n1_13833_12560 1.178286e+01
R2865 n1_13833_12560 n1_14021_12560 1.074286e+00
R2866 n1_14021_12560 n1_16083_12560 1.178286e+01
R2867 n1_16083_12560 n1_16271_12560 1.074286e+00
R2868 n1_16271_12560 n1_18333_12560 1.178286e+01
R2869 n1_18333_12560 n1_18521_12560 1.074286e+00
R2870 n1_18521_12560 n1_20583_12560 1.178286e+01
R2871 n1_20583_12560 n1_20771_12560 1.074286e+00
R2872 n1_333_12743 n1_521_12743 1.074286e+00
R2873 n1_521_12743 n1_2583_12743 1.178286e+01
R2874 n1_2583_12743 n1_2771_12743 1.074286e+00
R2875 n1_2771_12743 n1_4833_12743 1.178286e+01
R2876 n1_4833_12743 n1_5021_12743 1.074286e+00
R2877 n1_5021_12743 n1_7083_12743 1.178286e+01
R2878 n1_7083_12743 n1_7271_12743 1.074286e+00
R2879 n1_7271_12743 n1_9333_12743 1.178286e+01
R2880 n1_9333_12743 n1_9521_12743 1.074286e+00
R2881 n1_11583_12743 n1_11771_12743 1.074286e+00
R2882 n1_11771_12743 n1_13833_12743 1.178286e+01
R2883 n1_13833_12743 n1_14021_12743 1.074286e+00
R2884 n1_14021_12743 n1_16083_12743 1.178286e+01
R2885 n1_16083_12743 n1_16271_12743 1.074286e+00
R2886 n1_16271_12743 n1_18333_12743 1.178286e+01
R2887 n1_18333_12743 n1_18521_12743 1.074286e+00
R2888 n1_18521_12743 n1_20583_12743 1.178286e+01
R2889 n1_20583_12743 n1_20771_12743 1.074286e+00
R2890 n1_521_12776 n1_2771_12776 1.285714e+01
R2891 n1_2771_12776 n1_5021_12776 1.285714e+01
R2892 n1_5021_12776 n1_7271_12776 1.285714e+01
R2893 n1_7271_12776 n1_9521_12776 1.285714e+01
R2894 n1_11771_12776 n1_14021_12776 1.285714e+01
R2895 n1_14021_12776 n1_16271_12776 1.285714e+01
R2896 n1_16271_12776 n1_18521_12776 1.285714e+01
R2897 n1_18521_12776 n1_20771_12776 1.285714e+01
R2898 n1_333_12959 n1_521_12959 1.074286e+00
R2899 n1_521_12959 n1_2583_12959 1.178286e+01
R2900 n1_2583_12959 n1_2771_12959 1.074286e+00
R2901 n1_2771_12959 n1_4833_12959 1.178286e+01
R2902 n1_4833_12959 n1_5021_12959 1.074286e+00
R2903 n1_5021_12959 n1_7083_12959 1.178286e+01
R2904 n1_7083_12959 n1_7271_12959 1.074286e+00
R2905 n1_7271_12959 n1_9333_12959 1.178286e+01
R2906 n1_9333_12959 n1_9521_12959 1.074286e+00
R2907 n1_11583_12959 n1_11771_12959 1.074286e+00
R2908 n1_11771_12959 n1_13833_12959 1.178286e+01
R2909 n1_13833_12959 n1_14021_12959 1.074286e+00
R2910 n1_14021_12959 n1_16083_12959 1.178286e+01
R2911 n1_16083_12959 n1_16271_12959 1.074286e+00
R2912 n1_16271_12959 n1_18333_12959 1.178286e+01
R2913 n1_18333_12959 n1_18521_12959 1.074286e+00
R2914 n1_18521_12959 n1_20583_12959 1.178286e+01
R2915 n1_20583_12959 n1_20771_12959 1.074286e+00
R2916 n1_333_12992 n1_521_12992 1.074286e+00
R2917 n1_521_12992 n1_2583_12992 1.178286e+01
R2918 n1_2583_12992 n1_2771_12992 1.074286e+00
R2919 n1_2771_12992 n1_4833_12992 1.178286e+01
R2920 n1_4833_12992 n1_5021_12992 1.074286e+00
R2921 n1_5021_12992 n1_7083_12992 1.178286e+01
R2922 n1_7083_12992 n1_7271_12992 1.074286e+00
R2923 n1_7271_12992 n1_9333_12992 1.178286e+01
R2924 n1_9333_12992 n1_9521_12992 1.074286e+00
R2925 n1_11583_12992 n1_11771_12992 1.074286e+00
R2926 n1_11771_12992 n1_13833_12992 1.178286e+01
R2927 n1_13833_12992 n1_14021_12992 1.074286e+00
R2928 n1_14021_12992 n1_16083_12992 1.178286e+01
R2929 n1_16083_12992 n1_16271_12992 1.074286e+00
R2930 n1_16271_12992 n1_18333_12992 1.178286e+01
R2931 n1_18333_12992 n1_18521_12992 1.074286e+00
R2932 n1_18521_12992 n1_20583_12992 1.178286e+01
R2933 n1_20583_12992 n1_20771_12992 1.074286e+00
R2934 n1_333_13175 n1_521_13175 1.074286e+00
R2935 n1_521_13175 n1_2583_13175 1.178286e+01
R2936 n1_2583_13175 n1_2771_13175 1.074286e+00
R2937 n1_2771_13175 n1_4833_13175 1.178286e+01
R2938 n1_4833_13175 n1_5021_13175 1.074286e+00
R2939 n1_5021_13175 n1_7083_13175 1.178286e+01
R2940 n1_7083_13175 n1_7271_13175 1.074286e+00
R2941 n1_7271_13175 n1_9333_13175 1.178286e+01
R2942 n1_9333_13175 n1_9521_13175 1.074286e+00
R2943 n1_11583_13175 n1_11771_13175 1.074286e+00
R2944 n1_11771_13175 n1_13833_13175 1.178286e+01
R2945 n1_13833_13175 n1_14021_13175 1.074286e+00
R2946 n1_14021_13175 n1_16083_13175 1.178286e+01
R2947 n1_16083_13175 n1_16271_13175 1.074286e+00
R2948 n1_16271_13175 n1_18333_13175 1.178286e+01
R2949 n1_18333_13175 n1_18521_13175 1.074286e+00
R2950 n1_18521_13175 n1_20583_13175 1.178286e+01
R2951 n1_20583_13175 n1_20771_13175 1.074286e+00
R2952 n1_333_13208 n1_521_13208 1.074286e+00
R2953 n1_521_13208 n1_2583_13208 1.178286e+01
R2954 n1_2583_13208 n1_2771_13208 1.074286e+00
R2955 n1_2771_13208 n1_4833_13208 1.178286e+01
R2956 n1_4833_13208 n1_5021_13208 1.074286e+00
R2957 n1_5021_13208 n1_7083_13208 1.178286e+01
R2958 n1_7083_13208 n1_7271_13208 1.074286e+00
R2959 n1_7271_13208 n1_9333_13208 1.178286e+01
R2960 n1_9333_13208 n1_9521_13208 1.074286e+00
R2961 n1_11583_13208 n1_11771_13208 1.074286e+00
R2962 n1_11771_13208 n1_13833_13208 1.178286e+01
R2963 n1_13833_13208 n1_14021_13208 1.074286e+00
R2964 n1_14021_13208 n1_16083_13208 1.178286e+01
R2965 n1_16083_13208 n1_16271_13208 1.074286e+00
R2966 n1_16271_13208 n1_18333_13208 1.178286e+01
R2967 n1_18333_13208 n1_18521_13208 1.074286e+00
R2968 n1_18521_13208 n1_20583_13208 1.178286e+01
R2969 n1_20583_13208 n1_20771_13208 1.074286e+00
R2970 n1_333_13391 n1_521_13391 1.074286e+00
R2971 n1_521_13391 n1_2583_13391 1.178286e+01
R2972 n1_2583_13391 n1_2771_13391 1.074286e+00
R2973 n1_2771_13391 n1_4833_13391 1.178286e+01
R2974 n1_4833_13391 n1_5021_13391 1.074286e+00
R2975 n1_5021_13391 n1_7083_13391 1.178286e+01
R2976 n1_7083_13391 n1_7271_13391 1.074286e+00
R2977 n1_7271_13391 n1_9333_13391 1.178286e+01
R2978 n1_9333_13391 n1_9521_13391 1.074286e+00
R2979 n1_11583_13391 n1_11771_13391 1.074286e+00
R2980 n1_11771_13391 n1_13833_13391 1.178286e+01
R2981 n1_13833_13391 n1_14021_13391 1.074286e+00
R2982 n1_14021_13391 n1_16083_13391 1.178286e+01
R2983 n1_16083_13391 n1_16271_13391 1.074286e+00
R2984 n1_16271_13391 n1_18333_13391 1.178286e+01
R2985 n1_18333_13391 n1_18521_13391 1.074286e+00
R2986 n1_18521_13391 n1_20583_13391 1.178286e+01
R2987 n1_20583_13391 n1_20771_13391 1.074286e+00
R2988 n1_333_13424 n1_521_13424 1.074286e+00
R2989 n1_521_13424 n1_2583_13424 1.178286e+01
R2990 n1_2583_13424 n1_2771_13424 1.074286e+00
R2991 n1_2771_13424 n1_4833_13424 1.178286e+01
R2992 n1_4833_13424 n1_5021_13424 1.074286e+00
R2993 n1_5021_13424 n1_7083_13424 1.178286e+01
R2994 n1_7083_13424 n1_7271_13424 1.074286e+00
R2995 n1_7271_13424 n1_9333_13424 1.178286e+01
R2996 n1_9333_13424 n1_9521_13424 1.074286e+00
R2997 n1_11583_13424 n1_11771_13424 1.074286e+00
R2998 n1_11771_13424 n1_13833_13424 1.178286e+01
R2999 n1_13833_13424 n1_14021_13424 1.074286e+00
R3000 n1_14021_13424 n1_16083_13424 1.178286e+01
R3001 n1_16083_13424 n1_16271_13424 1.074286e+00
R3002 n1_16271_13424 n1_18333_13424 1.178286e+01
R3003 n1_18333_13424 n1_18521_13424 1.074286e+00
R3004 n1_18521_13424 n1_20583_13424 1.178286e+01
R3005 n1_20583_13424 n1_20771_13424 1.074286e+00
R3006 n1_333_13607 n1_521_13607 1.074286e+00
R3007 n1_521_13607 n1_2583_13607 1.178286e+01
R3008 n1_2583_13607 n1_2771_13607 1.074286e+00
R3009 n1_2771_13607 n1_4833_13607 1.178286e+01
R3010 n1_4833_13607 n1_5021_13607 1.074286e+00
R3011 n1_5021_13607 n1_7083_13607 1.178286e+01
R3012 n1_7083_13607 n1_7271_13607 1.074286e+00
R3013 n1_7271_13607 n1_9333_13607 1.178286e+01
R3014 n1_9333_13607 n1_9521_13607 1.074286e+00
R3015 n1_11583_13607 n1_11771_13607 1.074286e+00
R3016 n1_11771_13607 n1_13833_13607 1.178286e+01
R3017 n1_13833_13607 n1_14021_13607 1.074286e+00
R3018 n1_14021_13607 n1_16083_13607 1.178286e+01
R3019 n1_16083_13607 n1_16271_13607 1.074286e+00
R3020 n1_16271_13607 n1_18333_13607 1.178286e+01
R3021 n1_18333_13607 n1_18521_13607 1.074286e+00
R3022 n1_18521_13607 n1_20583_13607 1.178286e+01
R3023 n1_20583_13607 n1_20771_13607 1.074286e+00
R3024 n1_333_13640 n1_521_13640 1.074286e+00
R3025 n1_521_13640 n1_2583_13640 1.178286e+01
R3026 n1_2583_13640 n1_2771_13640 1.074286e+00
R3027 n1_2771_13640 n1_4833_13640 1.178286e+01
R3028 n1_4833_13640 n1_5021_13640 1.074286e+00
R3029 n1_5021_13640 n1_7083_13640 1.178286e+01
R3030 n1_7083_13640 n1_7271_13640 1.074286e+00
R3031 n1_7271_13640 n1_9333_13640 1.178286e+01
R3032 n1_9333_13640 n1_9521_13640 1.074286e+00
R3033 n1_11583_13640 n1_11771_13640 1.074286e+00
R3034 n1_11771_13640 n1_13833_13640 1.178286e+01
R3035 n1_13833_13640 n1_14021_13640 1.074286e+00
R3036 n1_14021_13640 n1_16083_13640 1.178286e+01
R3037 n1_16083_13640 n1_16271_13640 1.074286e+00
R3038 n1_16271_13640 n1_18333_13640 1.178286e+01
R3039 n1_18333_13640 n1_18521_13640 1.074286e+00
R3040 n1_18521_13640 n1_20583_13640 1.178286e+01
R3041 n1_20583_13640 n1_20771_13640 1.074286e+00
R3042 n1_333_13823 n1_521_13823 1.074286e+00
R3043 n1_521_13823 n1_2583_13823 1.178286e+01
R3044 n1_2583_13823 n1_2771_13823 1.074286e+00
R3045 n1_2771_13823 n1_4833_13823 1.178286e+01
R3046 n1_4833_13823 n1_5021_13823 1.074286e+00
R3047 n1_5021_13823 n1_7083_13823 1.178286e+01
R3048 n1_7083_13823 n1_7271_13823 1.074286e+00
R3049 n1_7271_13823 n1_9333_13823 1.178286e+01
R3050 n1_9333_13823 n1_9521_13823 1.074286e+00
R3051 n1_11583_13823 n1_11771_13823 1.074286e+00
R3052 n1_11771_13823 n1_13833_13823 1.178286e+01
R3053 n1_13833_13823 n1_14021_13823 1.074286e+00
R3054 n1_14021_13823 n1_16083_13823 1.178286e+01
R3055 n1_16083_13823 n1_16271_13823 1.074286e+00
R3056 n1_16271_13823 n1_18333_13823 1.178286e+01
R3057 n1_18333_13823 n1_18521_13823 1.074286e+00
R3058 n1_18521_13823 n1_20583_13823 1.178286e+01
R3059 n1_20583_13823 n1_20771_13823 1.074286e+00
R3060 n1_333_13856 n1_521_13856 1.074286e+00
R3061 n1_521_13856 n1_2583_13856 1.178286e+01
R3062 n1_2583_13856 n1_2771_13856 1.074286e+00
R3063 n1_2771_13856 n1_4833_13856 1.178286e+01
R3064 n1_4833_13856 n1_5021_13856 1.074286e+00
R3065 n1_5021_13856 n1_7083_13856 1.178286e+01
R3066 n1_7083_13856 n1_7271_13856 1.074286e+00
R3067 n1_7271_13856 n1_9333_13856 1.178286e+01
R3068 n1_9333_13856 n1_9521_13856 1.074286e+00
R3069 n1_11583_13856 n1_11771_13856 1.074286e+00
R3070 n1_11771_13856 n1_13833_13856 1.178286e+01
R3071 n1_13833_13856 n1_14021_13856 1.074286e+00
R3072 n1_14021_13856 n1_16083_13856 1.178286e+01
R3073 n1_16083_13856 n1_16271_13856 1.074286e+00
R3074 n1_16271_13856 n1_18333_13856 1.178286e+01
R3075 n1_18333_13856 n1_18521_13856 1.074286e+00
R3076 n1_18521_13856 n1_20583_13856 1.178286e+01
R3077 n1_20583_13856 n1_20771_13856 1.074286e+00
R3078 n1_333_14039 n1_380_14039 2.685714e-01
R3079 n1_380_14039 n1_521_14039 8.057143e-01
R3080 n1_521_14039 n1_2583_14039 1.178286e+01
R3081 n1_2583_14039 n1_2630_14039 2.685714e-01
R3082 n1_2630_14039 n1_2771_14039 8.057143e-01
R3083 n1_2771_14039 n1_4833_14039 1.178286e+01
R3084 n1_4833_14039 n1_4880_14039 2.685714e-01
R3085 n1_4880_14039 n1_5021_14039 8.057143e-01
R3086 n1_5021_14039 n1_7083_14039 1.178286e+01
R3087 n1_7083_14039 n1_7130_14039 2.685714e-01
R3088 n1_7130_14039 n1_7271_14039 8.057143e-01
R3089 n1_7271_14039 n1_9333_14039 1.178286e+01
R3090 n1_9333_14039 n1_9380_14039 2.685714e-01
R3091 n1_9380_14039 n1_9521_14039 8.057143e-01
R3092 n1_11583_14039 n1_11630_14039 2.685714e-01
R3093 n1_11630_14039 n1_11771_14039 8.057143e-01
R3094 n1_11771_14039 n1_13833_14039 1.178286e+01
R3095 n1_13833_14039 n1_13880_14039 2.685714e-01
R3096 n1_13880_14039 n1_14021_14039 8.057143e-01
R3097 n1_14021_14039 n1_16083_14039 1.178286e+01
R3098 n1_16083_14039 n1_16130_14039 2.685714e-01
R3099 n1_16130_14039 n1_16271_14039 8.057143e-01
R3100 n1_16271_14039 n1_18333_14039 1.178286e+01
R3101 n1_18333_14039 n1_18380_14039 2.685714e-01
R3102 n1_18380_14039 n1_18521_14039 8.057143e-01
R3103 n1_18521_14039 n1_20583_14039 1.178286e+01
R3104 n1_20583_14039 n1_20630_14039 2.685714e-01
R3105 n1_20630_14039 n1_20771_14039 8.057143e-01
R3106 n1_333_14072 n1_521_14072 1.074286e+00
R3107 n1_521_14072 n1_2583_14072 1.178286e+01
R3108 n1_2583_14072 n1_2771_14072 1.074286e+00
R3109 n1_2771_14072 n1_4833_14072 1.178286e+01
R3110 n1_4833_14072 n1_5021_14072 1.074286e+00
R3111 n1_5021_14072 n1_7083_14072 1.178286e+01
R3112 n1_7083_14072 n1_7271_14072 1.074286e+00
R3113 n1_7271_14072 n1_9333_14072 1.178286e+01
R3114 n1_9333_14072 n1_9521_14072 1.074286e+00
R3115 n1_11583_14072 n1_11771_14072 1.074286e+00
R3116 n1_11771_14072 n1_13833_14072 1.178286e+01
R3117 n1_13833_14072 n1_14021_14072 1.074286e+00
R3118 n1_14021_14072 n1_16083_14072 1.178286e+01
R3119 n1_16083_14072 n1_16271_14072 1.074286e+00
R3120 n1_16271_14072 n1_18333_14072 1.178286e+01
R3121 n1_18333_14072 n1_18521_14072 1.074286e+00
R3122 n1_18521_14072 n1_20583_14072 1.178286e+01
R3123 n1_20583_14072 n1_20771_14072 1.074286e+00
R3124 n1_333_14255 n1_521_14255 1.074286e+00
R3125 n1_521_14255 n1_2583_14255 1.178286e+01
R3126 n1_2583_14255 n1_2771_14255 1.074286e+00
R3127 n1_2771_14255 n1_4833_14255 1.178286e+01
R3128 n1_4833_14255 n1_5021_14255 1.074286e+00
R3129 n1_5021_14255 n1_7083_14255 1.178286e+01
R3130 n1_7083_14255 n1_7271_14255 1.074286e+00
R3131 n1_7271_14255 n1_9333_14255 1.178286e+01
R3132 n1_9333_14255 n1_9521_14255 1.074286e+00
R3133 n1_11583_14255 n1_11771_14255 1.074286e+00
R3134 n1_11771_14255 n1_13833_14255 1.178286e+01
R3135 n1_13833_14255 n1_14021_14255 1.074286e+00
R3136 n1_14021_14255 n1_16083_14255 1.178286e+01
R3137 n1_16083_14255 n1_16271_14255 1.074286e+00
R3138 n1_16271_14255 n1_18333_14255 1.178286e+01
R3139 n1_18333_14255 n1_18521_14255 1.074286e+00
R3140 n1_18521_14255 n1_20583_14255 1.178286e+01
R3141 n1_20583_14255 n1_20771_14255 1.074286e+00
R3142 n1_333_14288 n1_521_14288 1.074286e+00
R3143 n1_521_14288 n1_2583_14288 1.178286e+01
R3144 n1_2583_14288 n1_2771_14288 1.074286e+00
R3145 n1_2771_14288 n1_4833_14288 1.178286e+01
R3146 n1_4833_14288 n1_5021_14288 1.074286e+00
R3147 n1_5021_14288 n1_7083_14288 1.178286e+01
R3148 n1_7083_14288 n1_7271_14288 1.074286e+00
R3149 n1_7271_14288 n1_9333_14288 1.178286e+01
R3150 n1_9333_14288 n1_9521_14288 1.074286e+00
R3151 n1_11583_14288 n1_11771_14288 1.074286e+00
R3152 n1_11771_14288 n1_13833_14288 1.178286e+01
R3153 n1_13833_14288 n1_14021_14288 1.074286e+00
R3154 n1_14021_14288 n1_16083_14288 1.178286e+01
R3155 n1_16083_14288 n1_16271_14288 1.074286e+00
R3156 n1_16271_14288 n1_18333_14288 1.178286e+01
R3157 n1_18333_14288 n1_18521_14288 1.074286e+00
R3158 n1_18521_14288 n1_20583_14288 1.178286e+01
R3159 n1_20583_14288 n1_20771_14288 1.074286e+00
R3160 n1_333_14471 n1_521_14471 1.074286e+00
R3161 n1_521_14471 n1_2583_14471 1.178286e+01
R3162 n1_2583_14471 n1_2771_14471 1.074286e+00
R3163 n1_2771_14471 n1_4833_14471 1.178286e+01
R3164 n1_4833_14471 n1_5021_14471 1.074286e+00
R3165 n1_5021_14471 n1_7083_14471 1.178286e+01
R3166 n1_7083_14471 n1_7271_14471 1.074286e+00
R3167 n1_7271_14471 n1_9333_14471 1.178286e+01
R3168 n1_9333_14471 n1_9521_14471 1.074286e+00
R3169 n1_11583_14471 n1_11771_14471 1.074286e+00
R3170 n1_11771_14471 n1_13833_14471 1.178286e+01
R3171 n1_13833_14471 n1_14021_14471 1.074286e+00
R3172 n1_14021_14471 n1_16083_14471 1.178286e+01
R3173 n1_16083_14471 n1_16271_14471 1.074286e+00
R3174 n1_16271_14471 n1_18333_14471 1.178286e+01
R3175 n1_18333_14471 n1_18521_14471 1.074286e+00
R3176 n1_18521_14471 n1_20583_14471 1.178286e+01
R3177 n1_20583_14471 n1_20771_14471 1.074286e+00
R3178 n1_333_14504 n1_521_14504 1.074286e+00
R3179 n1_521_14504 n1_2583_14504 1.178286e+01
R3180 n1_2583_14504 n1_2771_14504 1.074286e+00
R3181 n1_2771_14504 n1_4833_14504 1.178286e+01
R3182 n1_4833_14504 n1_5021_14504 1.074286e+00
R3183 n1_5021_14504 n1_7083_14504 1.178286e+01
R3184 n1_7083_14504 n1_7271_14504 1.074286e+00
R3185 n1_7271_14504 n1_9333_14504 1.178286e+01
R3186 n1_9333_14504 n1_9521_14504 1.074286e+00
R3187 n1_11583_14504 n1_11771_14504 1.074286e+00
R3188 n1_11771_14504 n1_13833_14504 1.178286e+01
R3189 n1_13833_14504 n1_14021_14504 1.074286e+00
R3190 n1_14021_14504 n1_16083_14504 1.178286e+01
R3191 n1_16083_14504 n1_16271_14504 1.074286e+00
R3192 n1_16271_14504 n1_18333_14504 1.178286e+01
R3193 n1_18333_14504 n1_18521_14504 1.074286e+00
R3194 n1_18521_14504 n1_20583_14504 1.178286e+01
R3195 n1_20583_14504 n1_20771_14504 1.074286e+00
R3196 n1_333_14687 n1_521_14687 1.074286e+00
R3197 n1_521_14687 n1_2583_14687 1.178286e+01
R3198 n1_2583_14687 n1_2771_14687 1.074286e+00
R3199 n1_2771_14687 n1_4833_14687 1.178286e+01
R3200 n1_4833_14687 n1_5021_14687 1.074286e+00
R3201 n1_5021_14687 n1_7083_14687 1.178286e+01
R3202 n1_7083_14687 n1_7271_14687 1.074286e+00
R3203 n1_7271_14687 n1_9333_14687 1.178286e+01
R3204 n1_9333_14687 n1_9521_14687 1.074286e+00
R3205 n1_11583_14687 n1_11771_14687 1.074286e+00
R3206 n1_11771_14687 n1_13833_14687 1.178286e+01
R3207 n1_13833_14687 n1_14021_14687 1.074286e+00
R3208 n1_14021_14687 n1_16083_14687 1.178286e+01
R3209 n1_16083_14687 n1_16271_14687 1.074286e+00
R3210 n1_16271_14687 n1_18333_14687 1.178286e+01
R3211 n1_18333_14687 n1_18521_14687 1.074286e+00
R3212 n1_18521_14687 n1_20583_14687 1.178286e+01
R3213 n1_20583_14687 n1_20771_14687 1.074286e+00
R3214 n1_333_14720 n1_521_14720 1.074286e+00
R3215 n1_521_14720 n1_2583_14720 1.178286e+01
R3216 n1_2583_14720 n1_2771_14720 1.074286e+00
R3217 n1_2771_14720 n1_4833_14720 1.178286e+01
R3218 n1_4833_14720 n1_5021_14720 1.074286e+00
R3219 n1_5021_14720 n1_7083_14720 1.178286e+01
R3220 n1_7083_14720 n1_7271_14720 1.074286e+00
R3221 n1_7271_14720 n1_9333_14720 1.178286e+01
R3222 n1_9333_14720 n1_9521_14720 1.074286e+00
R3223 n1_11583_14720 n1_11771_14720 1.074286e+00
R3224 n1_11771_14720 n1_13833_14720 1.178286e+01
R3225 n1_13833_14720 n1_14021_14720 1.074286e+00
R3226 n1_14021_14720 n1_16083_14720 1.178286e+01
R3227 n1_16083_14720 n1_16271_14720 1.074286e+00
R3228 n1_16271_14720 n1_18333_14720 1.178286e+01
R3229 n1_18333_14720 n1_18521_14720 1.074286e+00
R3230 n1_18521_14720 n1_20583_14720 1.178286e+01
R3231 n1_20583_14720 n1_20771_14720 1.074286e+00
R3232 n1_333_14903 n1_521_14903 1.074286e+00
R3233 n1_521_14903 n1_2583_14903 1.178286e+01
R3234 n1_2583_14903 n1_2771_14903 1.074286e+00
R3235 n1_2771_14903 n1_4833_14903 1.178286e+01
R3236 n1_4833_14903 n1_5021_14903 1.074286e+00
R3237 n1_5021_14903 n1_7083_14903 1.178286e+01
R3238 n1_7083_14903 n1_7271_14903 1.074286e+00
R3239 n1_7271_14903 n1_9333_14903 1.178286e+01
R3240 n1_9333_14903 n1_9521_14903 1.074286e+00
R3241 n1_11583_14903 n1_11771_14903 1.074286e+00
R3242 n1_11771_14903 n1_13833_14903 1.178286e+01
R3243 n1_13833_14903 n1_14021_14903 1.074286e+00
R3244 n1_14021_14903 n1_16083_14903 1.178286e+01
R3245 n1_16083_14903 n1_16271_14903 1.074286e+00
R3246 n1_16271_14903 n1_18333_14903 1.178286e+01
R3247 n1_18333_14903 n1_18521_14903 1.074286e+00
R3248 n1_18521_14903 n1_20583_14903 1.178286e+01
R3249 n1_20583_14903 n1_20771_14903 1.074286e+00
R3250 n1_333_14936 n1_521_14936 1.074286e+00
R3251 n1_521_14936 n1_2583_14936 1.178286e+01
R3252 n1_2583_14936 n1_2771_14936 1.074286e+00
R3253 n1_2771_14936 n1_4833_14936 1.178286e+01
R3254 n1_4833_14936 n1_5021_14936 1.074286e+00
R3255 n1_5021_14936 n1_7083_14936 1.178286e+01
R3256 n1_7083_14936 n1_7271_14936 1.074286e+00
R3257 n1_7271_14936 n1_9333_14936 1.178286e+01
R3258 n1_9333_14936 n1_9521_14936 1.074286e+00
R3259 n1_11583_14936 n1_11771_14936 1.074286e+00
R3260 n1_11771_14936 n1_13833_14936 1.178286e+01
R3261 n1_13833_14936 n1_14021_14936 1.074286e+00
R3262 n1_14021_14936 n1_16083_14936 1.178286e+01
R3263 n1_16083_14936 n1_16271_14936 1.074286e+00
R3264 n1_16271_14936 n1_18333_14936 1.178286e+01
R3265 n1_18333_14936 n1_18521_14936 1.074286e+00
R3266 n1_18521_14936 n1_20583_14936 1.178286e+01
R3267 n1_20583_14936 n1_20771_14936 1.074286e+00
R3268 n1_521_15119 n1_2771_15119 1.285714e+01
R3269 n1_2771_15119 n1_5021_15119 1.285714e+01
R3270 n1_5021_15119 n1_7271_15119 1.285714e+01
R3271 n1_7271_15119 n1_9521_15119 1.285714e+01
R3272 n1_11771_15119 n1_14021_15119 1.285714e+01
R3273 n1_14021_15119 n1_16271_15119 1.285714e+01
R3274 n1_16271_15119 n1_18521_15119 1.285714e+01
R3275 n1_18521_15119 n1_20771_15119 1.285714e+01
R3276 n1_521_15152 n1_2771_15152 1.285714e+01
R3277 n1_2771_15152 n1_5021_15152 1.285714e+01
R3278 n1_5021_15152 n1_7271_15152 1.285714e+01
R3279 n1_7271_15152 n1_9521_15152 1.285714e+01
R3280 n1_11771_15152 n1_14021_15152 1.285714e+01
R3281 n1_14021_15152 n1_16271_15152 1.285714e+01
R3282 n1_16271_15152 n1_18521_15152 1.285714e+01
R3283 n1_18521_15152 n1_20771_15152 1.285714e+01
R3284 n1_333_15335 n1_521_15335 1.074286e+00
R3285 n1_521_15335 n1_2583_15335 1.178286e+01
R3286 n1_2583_15335 n1_2771_15335 1.074286e+00
R3287 n1_2771_15335 n1_4833_15335 1.178286e+01
R3288 n1_4833_15335 n1_5021_15335 1.074286e+00
R3289 n1_5021_15335 n1_7083_15335 1.178286e+01
R3290 n1_7083_15335 n1_7271_15335 1.074286e+00
R3291 n1_7271_15335 n1_9333_15335 1.178286e+01
R3292 n1_9333_15335 n1_9521_15335 1.074286e+00
R3293 n1_11583_15335 n1_11771_15335 1.074286e+00
R3294 n1_11771_15335 n1_13833_15335 1.178286e+01
R3295 n1_13833_15335 n1_14021_15335 1.074286e+00
R3296 n1_14021_15335 n1_16083_15335 1.178286e+01
R3297 n1_16083_15335 n1_16271_15335 1.074286e+00
R3298 n1_16271_15335 n1_18333_15335 1.178286e+01
R3299 n1_18333_15335 n1_18521_15335 1.074286e+00
R3300 n1_18521_15335 n1_20583_15335 1.178286e+01
R3301 n1_20583_15335 n1_20771_15335 1.074286e+00
R3302 n1_333_15368 n1_521_15368 1.074286e+00
R3303 n1_521_15368 n1_2583_15368 1.178286e+01
R3304 n1_2583_15368 n1_2771_15368 1.074286e+00
R3305 n1_2771_15368 n1_4833_15368 1.178286e+01
R3306 n1_4833_15368 n1_5021_15368 1.074286e+00
R3307 n1_5021_15368 n1_7083_15368 1.178286e+01
R3308 n1_7083_15368 n1_7271_15368 1.074286e+00
R3309 n1_7271_15368 n1_9333_15368 1.178286e+01
R3310 n1_9333_15368 n1_9521_15368 1.074286e+00
R3311 n1_11583_15368 n1_11771_15368 1.074286e+00
R3312 n1_11771_15368 n1_13833_15368 1.178286e+01
R3313 n1_13833_15368 n1_14021_15368 1.074286e+00
R3314 n1_14021_15368 n1_16083_15368 1.178286e+01
R3315 n1_16083_15368 n1_16271_15368 1.074286e+00
R3316 n1_16271_15368 n1_18333_15368 1.178286e+01
R3317 n1_18333_15368 n1_18521_15368 1.074286e+00
R3318 n1_18521_15368 n1_20583_15368 1.178286e+01
R3319 n1_20583_15368 n1_20771_15368 1.074286e+00
R3320 n1_333_15551 n1_521_15551 1.074286e+00
R3321 n1_521_15551 n1_2583_15551 1.178286e+01
R3322 n1_2583_15551 n1_2771_15551 1.074286e+00
R3323 n1_2771_15551 n1_4833_15551 1.178286e+01
R3324 n1_4833_15551 n1_5021_15551 1.074286e+00
R3325 n1_5021_15551 n1_7083_15551 1.178286e+01
R3326 n1_7083_15551 n1_7271_15551 1.074286e+00
R3327 n1_7271_15551 n1_9333_15551 1.178286e+01
R3328 n1_9333_15551 n1_9521_15551 1.074286e+00
R3329 n1_11583_15551 n1_11771_15551 1.074286e+00
R3330 n1_11771_15551 n1_13833_15551 1.178286e+01
R3331 n1_13833_15551 n1_14021_15551 1.074286e+00
R3332 n1_14021_15551 n1_16083_15551 1.178286e+01
R3333 n1_16083_15551 n1_16271_15551 1.074286e+00
R3334 n1_16271_15551 n1_18333_15551 1.178286e+01
R3335 n1_18333_15551 n1_18521_15551 1.074286e+00
R3336 n1_18521_15551 n1_20583_15551 1.178286e+01
R3337 n1_20583_15551 n1_20771_15551 1.074286e+00
R3338 n1_333_15584 n1_521_15584 1.074286e+00
R3339 n1_521_15584 n1_2583_15584 1.178286e+01
R3340 n1_2583_15584 n1_2771_15584 1.074286e+00
R3341 n1_2771_15584 n1_4833_15584 1.178286e+01
R3342 n1_4833_15584 n1_5021_15584 1.074286e+00
R3343 n1_5021_15584 n1_7083_15584 1.178286e+01
R3344 n1_7083_15584 n1_7271_15584 1.074286e+00
R3345 n1_7271_15584 n1_9333_15584 1.178286e+01
R3346 n1_9333_15584 n1_9521_15584 1.074286e+00
R3347 n1_11583_15584 n1_11771_15584 1.074286e+00
R3348 n1_11771_15584 n1_13833_15584 1.178286e+01
R3349 n1_13833_15584 n1_14021_15584 1.074286e+00
R3350 n1_14021_15584 n1_16083_15584 1.178286e+01
R3351 n1_16083_15584 n1_16271_15584 1.074286e+00
R3352 n1_16271_15584 n1_18333_15584 1.178286e+01
R3353 n1_18333_15584 n1_18521_15584 1.074286e+00
R3354 n1_18521_15584 n1_20583_15584 1.178286e+01
R3355 n1_20583_15584 n1_20771_15584 1.074286e+00
R3356 n1_333_15767 n1_521_15767 1.074286e+00
R3357 n1_521_15767 n1_2583_15767 1.178286e+01
R3358 n1_2583_15767 n1_2771_15767 1.074286e+00
R3359 n1_2771_15767 n1_4833_15767 1.178286e+01
R3360 n1_4833_15767 n1_5021_15767 1.074286e+00
R3361 n1_5021_15767 n1_7083_15767 1.178286e+01
R3362 n1_7083_15767 n1_7271_15767 1.074286e+00
R3363 n1_7271_15767 n1_9333_15767 1.178286e+01
R3364 n1_9333_15767 n1_9521_15767 1.074286e+00
R3365 n1_11583_15767 n1_11771_15767 1.074286e+00
R3366 n1_11771_15767 n1_13833_15767 1.178286e+01
R3367 n1_13833_15767 n1_14021_15767 1.074286e+00
R3368 n1_14021_15767 n1_16083_15767 1.178286e+01
R3369 n1_16083_15767 n1_16271_15767 1.074286e+00
R3370 n1_16271_15767 n1_18333_15767 1.178286e+01
R3371 n1_18333_15767 n1_18521_15767 1.074286e+00
R3372 n1_18521_15767 n1_20583_15767 1.178286e+01
R3373 n1_20583_15767 n1_20771_15767 1.074286e+00
R3374 n1_333_15800 n1_521_15800 1.074286e+00
R3375 n1_521_15800 n1_2583_15800 1.178286e+01
R3376 n1_2583_15800 n1_2771_15800 1.074286e+00
R3377 n1_2771_15800 n1_4833_15800 1.178286e+01
R3378 n1_4833_15800 n1_5021_15800 1.074286e+00
R3379 n1_5021_15800 n1_7083_15800 1.178286e+01
R3380 n1_7083_15800 n1_7271_15800 1.074286e+00
R3381 n1_7271_15800 n1_9333_15800 1.178286e+01
R3382 n1_9333_15800 n1_9521_15800 1.074286e+00
R3383 n1_11583_15800 n1_11771_15800 1.074286e+00
R3384 n1_11771_15800 n1_13833_15800 1.178286e+01
R3385 n1_13833_15800 n1_14021_15800 1.074286e+00
R3386 n1_14021_15800 n1_16083_15800 1.178286e+01
R3387 n1_16083_15800 n1_16271_15800 1.074286e+00
R3388 n1_16271_15800 n1_18333_15800 1.178286e+01
R3389 n1_18333_15800 n1_18521_15800 1.074286e+00
R3390 n1_18521_15800 n1_20583_15800 1.178286e+01
R3391 n1_20583_15800 n1_20771_15800 1.074286e+00
R3392 n1_333_15983 n1_521_15983 1.074286e+00
R3393 n1_521_15983 n1_2583_15983 1.178286e+01
R3394 n1_2583_15983 n1_2771_15983 1.074286e+00
R3395 n1_2771_15983 n1_4833_15983 1.178286e+01
R3396 n1_4833_15983 n1_5021_15983 1.074286e+00
R3397 n1_5021_15983 n1_7083_15983 1.178286e+01
R3398 n1_7083_15983 n1_7271_15983 1.074286e+00
R3399 n1_7271_15983 n1_9333_15983 1.178286e+01
R3400 n1_9333_15983 n1_9521_15983 1.074286e+00
R3401 n1_11583_15983 n1_11771_15983 1.074286e+00
R3402 n1_11771_15983 n1_13833_15983 1.178286e+01
R3403 n1_13833_15983 n1_14021_15983 1.074286e+00
R3404 n1_14021_15983 n1_16083_15983 1.178286e+01
R3405 n1_16083_15983 n1_16271_15983 1.074286e+00
R3406 n1_16271_15983 n1_18333_15983 1.178286e+01
R3407 n1_18333_15983 n1_18521_15983 1.074286e+00
R3408 n1_18521_15983 n1_20583_15983 1.178286e+01
R3409 n1_20583_15983 n1_20771_15983 1.074286e+00
R3410 n1_333_16016 n1_521_16016 1.074286e+00
R3411 n1_521_16016 n1_2583_16016 1.178286e+01
R3412 n1_2583_16016 n1_2771_16016 1.074286e+00
R3413 n1_2771_16016 n1_4833_16016 1.178286e+01
R3414 n1_4833_16016 n1_5021_16016 1.074286e+00
R3415 n1_5021_16016 n1_7083_16016 1.178286e+01
R3416 n1_7083_16016 n1_7271_16016 1.074286e+00
R3417 n1_7271_16016 n1_9333_16016 1.178286e+01
R3418 n1_9333_16016 n1_9521_16016 1.074286e+00
R3419 n1_11583_16016 n1_11771_16016 1.074286e+00
R3420 n1_11771_16016 n1_13833_16016 1.178286e+01
R3421 n1_13833_16016 n1_14021_16016 1.074286e+00
R3422 n1_14021_16016 n1_16083_16016 1.178286e+01
R3423 n1_16083_16016 n1_16271_16016 1.074286e+00
R3424 n1_16271_16016 n1_18333_16016 1.178286e+01
R3425 n1_18333_16016 n1_18521_16016 1.074286e+00
R3426 n1_18521_16016 n1_20583_16016 1.178286e+01
R3427 n1_20583_16016 n1_20771_16016 1.074286e+00
R3428 n1_333_16199 n1_380_16199 2.685714e-01
R3429 n1_380_16199 n1_521_16199 8.057143e-01
R3430 n1_521_16199 n1_2583_16199 1.178286e+01
R3431 n1_2583_16199 n1_2630_16199 2.685714e-01
R3432 n1_2630_16199 n1_2771_16199 8.057143e-01
R3433 n1_2771_16199 n1_4833_16199 1.178286e+01
R3434 n1_4833_16199 n1_4880_16199 2.685714e-01
R3435 n1_4880_16199 n1_5021_16199 8.057143e-01
R3436 n1_5021_16199 n1_7083_16199 1.178286e+01
R3437 n1_7083_16199 n1_7130_16199 2.685714e-01
R3438 n1_7130_16199 n1_7271_16199 8.057143e-01
R3439 n1_7271_16199 n1_9333_16199 1.178286e+01
R3440 n1_9333_16199 n1_9380_16199 2.685714e-01
R3441 n1_9380_16199 n1_9521_16199 8.057143e-01
R3442 n1_11583_16199 n1_11630_16199 2.685714e-01
R3443 n1_11630_16199 n1_11771_16199 8.057143e-01
R3444 n1_11771_16199 n1_13833_16199 1.178286e+01
R3445 n1_13833_16199 n1_13880_16199 2.685714e-01
R3446 n1_13880_16199 n1_14021_16199 8.057143e-01
R3447 n1_14021_16199 n1_16083_16199 1.178286e+01
R3448 n1_16083_16199 n1_16130_16199 2.685714e-01
R3449 n1_16130_16199 n1_16271_16199 8.057143e-01
R3450 n1_16271_16199 n1_18333_16199 1.178286e+01
R3451 n1_18333_16199 n1_18380_16199 2.685714e-01
R3452 n1_18380_16199 n1_18521_16199 8.057143e-01
R3453 n1_18521_16199 n1_20583_16199 1.178286e+01
R3454 n1_20583_16199 n1_20630_16199 2.685714e-01
R3455 n1_20630_16199 n1_20771_16199 8.057143e-01
R3456 n1_333_16232 n1_380_16232 2.685714e-01
R3457 n1_380_16232 n1_2583_16232 1.258857e+01
R3458 n1_2583_16232 n1_2630_16232 2.685714e-01
R3459 n1_2630_16232 n1_4833_16232 1.258857e+01
R3460 n1_4833_16232 n1_4880_16232 2.685714e-01
R3461 n1_4880_16232 n1_7083_16232 1.258857e+01
R3462 n1_7083_16232 n1_7130_16232 2.685714e-01
R3463 n1_7130_16232 n1_9333_16232 1.258857e+01
R3464 n1_9333_16232 n1_9380_16232 2.685714e-01
R3465 n1_11583_16232 n1_11630_16232 2.685714e-01
R3466 n1_11630_16232 n1_13833_16232 1.258857e+01
R3467 n1_13833_16232 n1_13880_16232 2.685714e-01
R3468 n1_13880_16232 n1_16083_16232 1.258857e+01
R3469 n1_16083_16232 n1_16130_16232 2.685714e-01
R3470 n1_16130_16232 n1_18333_16232 1.258857e+01
R3471 n1_18333_16232 n1_18380_16232 2.685714e-01
R3472 n1_18380_16232 n1_20583_16232 1.258857e+01
R3473 n1_20583_16232 n1_20630_16232 2.685714e-01
R3474 n1_333_16415 n1_521_16415 1.074286e+00
R3475 n1_521_16415 n1_2583_16415 1.178286e+01
R3476 n1_2583_16415 n1_2771_16415 1.074286e+00
R3477 n1_2771_16415 n1_4833_16415 1.178286e+01
R3478 n1_4833_16415 n1_5021_16415 1.074286e+00
R3479 n1_5021_16415 n1_7083_16415 1.178286e+01
R3480 n1_7083_16415 n1_7271_16415 1.074286e+00
R3481 n1_7271_16415 n1_9333_16415 1.178286e+01
R3482 n1_9333_16415 n1_9521_16415 1.074286e+00
R3483 n1_11583_16415 n1_11771_16415 1.074286e+00
R3484 n1_11771_16415 n1_13833_16415 1.178286e+01
R3485 n1_13833_16415 n1_14021_16415 1.074286e+00
R3486 n1_14021_16415 n1_16083_16415 1.178286e+01
R3487 n1_16083_16415 n1_16271_16415 1.074286e+00
R3488 n1_16271_16415 n1_18333_16415 1.178286e+01
R3489 n1_18333_16415 n1_18521_16415 1.074286e+00
R3490 n1_18521_16415 n1_20583_16415 1.178286e+01
R3491 n1_20583_16415 n1_20771_16415 1.074286e+00
R3492 n1_333_16448 n1_521_16448 1.074286e+00
R3493 n1_521_16448 n1_2583_16448 1.178286e+01
R3494 n1_2583_16448 n1_2771_16448 1.074286e+00
R3495 n1_2771_16448 n1_4833_16448 1.178286e+01
R3496 n1_4833_16448 n1_5021_16448 1.074286e+00
R3497 n1_5021_16448 n1_7083_16448 1.178286e+01
R3498 n1_7083_16448 n1_7271_16448 1.074286e+00
R3499 n1_7271_16448 n1_9333_16448 1.178286e+01
R3500 n1_9333_16448 n1_9521_16448 1.074286e+00
R3501 n1_11583_16448 n1_11771_16448 1.074286e+00
R3502 n1_11771_16448 n1_13833_16448 1.178286e+01
R3503 n1_13833_16448 n1_14021_16448 1.074286e+00
R3504 n1_14021_16448 n1_16083_16448 1.178286e+01
R3505 n1_16083_16448 n1_16271_16448 1.074286e+00
R3506 n1_16271_16448 n1_18333_16448 1.178286e+01
R3507 n1_18333_16448 n1_18521_16448 1.074286e+00
R3508 n1_18521_16448 n1_20583_16448 1.178286e+01
R3509 n1_20583_16448 n1_20771_16448 1.074286e+00
R3510 n1_333_16631 n1_521_16631 1.074286e+00
R3511 n1_521_16631 n1_2583_16631 1.178286e+01
R3512 n1_2583_16631 n1_2771_16631 1.074286e+00
R3513 n1_2771_16631 n1_4833_16631 1.178286e+01
R3514 n1_4833_16631 n1_5021_16631 1.074286e+00
R3515 n1_5021_16631 n1_7083_16631 1.178286e+01
R3516 n1_7083_16631 n1_7271_16631 1.074286e+00
R3517 n1_7271_16631 n1_9333_16631 1.178286e+01
R3518 n1_9333_16631 n1_9521_16631 1.074286e+00
R3519 n1_11583_16631 n1_11771_16631 1.074286e+00
R3520 n1_11771_16631 n1_13833_16631 1.178286e+01
R3521 n1_13833_16631 n1_14021_16631 1.074286e+00
R3522 n1_14021_16631 n1_16083_16631 1.178286e+01
R3523 n1_16083_16631 n1_16271_16631 1.074286e+00
R3524 n1_16271_16631 n1_18333_16631 1.178286e+01
R3525 n1_18333_16631 n1_18521_16631 1.074286e+00
R3526 n1_18521_16631 n1_20583_16631 1.178286e+01
R3527 n1_20583_16631 n1_20771_16631 1.074286e+00
R3528 n1_333_16664 n1_521_16664 1.074286e+00
R3529 n1_521_16664 n1_2583_16664 1.178286e+01
R3530 n1_2583_16664 n1_2771_16664 1.074286e+00
R3531 n1_2771_16664 n1_4833_16664 1.178286e+01
R3532 n1_4833_16664 n1_5021_16664 1.074286e+00
R3533 n1_5021_16664 n1_7083_16664 1.178286e+01
R3534 n1_7083_16664 n1_7271_16664 1.074286e+00
R3535 n1_7271_16664 n1_9333_16664 1.178286e+01
R3536 n1_9333_16664 n1_9521_16664 1.074286e+00
R3537 n1_11583_16664 n1_11771_16664 1.074286e+00
R3538 n1_11771_16664 n1_13833_16664 1.178286e+01
R3539 n1_13833_16664 n1_14021_16664 1.074286e+00
R3540 n1_14021_16664 n1_16083_16664 1.178286e+01
R3541 n1_16083_16664 n1_16271_16664 1.074286e+00
R3542 n1_16271_16664 n1_18333_16664 1.178286e+01
R3543 n1_18333_16664 n1_18521_16664 1.074286e+00
R3544 n1_18521_16664 n1_20583_16664 1.178286e+01
R3545 n1_20583_16664 n1_20771_16664 1.074286e+00
R3546 n1_333_16847 n1_521_16847 1.074286e+00
R3547 n1_521_16847 n1_2583_16847 1.178286e+01
R3548 n1_2583_16847 n1_2771_16847 1.074286e+00
R3549 n1_2771_16847 n1_4833_16847 1.178286e+01
R3550 n1_4833_16847 n1_5021_16847 1.074286e+00
R3551 n1_5021_16847 n1_7083_16847 1.178286e+01
R3552 n1_7083_16847 n1_7271_16847 1.074286e+00
R3553 n1_7271_16847 n1_9333_16847 1.178286e+01
R3554 n1_9333_16847 n1_9521_16847 1.074286e+00
R3555 n1_11583_16847 n1_11771_16847 1.074286e+00
R3556 n1_11771_16847 n1_13833_16847 1.178286e+01
R3557 n1_13833_16847 n1_14021_16847 1.074286e+00
R3558 n1_14021_16847 n1_16083_16847 1.178286e+01
R3559 n1_16083_16847 n1_16271_16847 1.074286e+00
R3560 n1_16271_16847 n1_18333_16847 1.178286e+01
R3561 n1_18333_16847 n1_18521_16847 1.074286e+00
R3562 n1_18521_16847 n1_20583_16847 1.178286e+01
R3563 n1_20583_16847 n1_20771_16847 1.074286e+00
R3564 n1_333_16880 n1_521_16880 1.074286e+00
R3565 n1_521_16880 n1_2583_16880 1.178286e+01
R3566 n1_2583_16880 n1_2771_16880 1.074286e+00
R3567 n1_2771_16880 n1_4833_16880 1.178286e+01
R3568 n1_4833_16880 n1_5021_16880 1.074286e+00
R3569 n1_5021_16880 n1_7083_16880 1.178286e+01
R3570 n1_7083_16880 n1_7271_16880 1.074286e+00
R3571 n1_7271_16880 n1_9333_16880 1.178286e+01
R3572 n1_9333_16880 n1_9521_16880 1.074286e+00
R3573 n1_11583_16880 n1_11771_16880 1.074286e+00
R3574 n1_11771_16880 n1_13833_16880 1.178286e+01
R3575 n1_13833_16880 n1_14021_16880 1.074286e+00
R3576 n1_14021_16880 n1_16083_16880 1.178286e+01
R3577 n1_16083_16880 n1_16271_16880 1.074286e+00
R3578 n1_16271_16880 n1_18333_16880 1.178286e+01
R3579 n1_18333_16880 n1_18521_16880 1.074286e+00
R3580 n1_18521_16880 n1_20583_16880 1.178286e+01
R3581 n1_20583_16880 n1_20771_16880 1.074286e+00
R3582 n1_333_17063 n1_521_17063 1.074286e+00
R3583 n1_521_17063 n1_2583_17063 1.178286e+01
R3584 n1_2583_17063 n1_2771_17063 1.074286e+00
R3585 n1_2771_17063 n1_4833_17063 1.178286e+01
R3586 n1_4833_17063 n1_5021_17063 1.074286e+00
R3587 n1_5021_17063 n1_7083_17063 1.178286e+01
R3588 n1_7083_17063 n1_7271_17063 1.074286e+00
R3589 n1_7271_17063 n1_9333_17063 1.178286e+01
R3590 n1_9333_17063 n1_9521_17063 1.074286e+00
R3591 n1_11583_17063 n1_11771_17063 1.074286e+00
R3592 n1_11771_17063 n1_13833_17063 1.178286e+01
R3593 n1_13833_17063 n1_14021_17063 1.074286e+00
R3594 n1_14021_17063 n1_16083_17063 1.178286e+01
R3595 n1_16083_17063 n1_16271_17063 1.074286e+00
R3596 n1_16271_17063 n1_18333_17063 1.178286e+01
R3597 n1_18333_17063 n1_18521_17063 1.074286e+00
R3598 n1_18521_17063 n1_20583_17063 1.178286e+01
R3599 n1_20583_17063 n1_20771_17063 1.074286e+00
R3600 n1_333_17096 n1_521_17096 1.074286e+00
R3601 n1_521_17096 n1_2583_17096 1.178286e+01
R3602 n1_2583_17096 n1_2771_17096 1.074286e+00
R3603 n1_2771_17096 n1_4833_17096 1.178286e+01
R3604 n1_4833_17096 n1_5021_17096 1.074286e+00
R3605 n1_5021_17096 n1_7083_17096 1.178286e+01
R3606 n1_7083_17096 n1_7271_17096 1.074286e+00
R3607 n1_7271_17096 n1_9333_17096 1.178286e+01
R3608 n1_9333_17096 n1_9521_17096 1.074286e+00
R3609 n1_11583_17096 n1_11771_17096 1.074286e+00
R3610 n1_11771_17096 n1_13833_17096 1.178286e+01
R3611 n1_13833_17096 n1_14021_17096 1.074286e+00
R3612 n1_14021_17096 n1_16083_17096 1.178286e+01
R3613 n1_16083_17096 n1_16271_17096 1.074286e+00
R3614 n1_16271_17096 n1_18333_17096 1.178286e+01
R3615 n1_18333_17096 n1_18521_17096 1.074286e+00
R3616 n1_18521_17096 n1_20583_17096 1.178286e+01
R3617 n1_20583_17096 n1_20771_17096 1.074286e+00
R3618 n1_521_17279 n1_2771_17279 1.285714e+01
R3619 n1_2771_17279 n1_5021_17279 1.285714e+01
R3620 n1_5021_17279 n1_7271_17279 1.285714e+01
R3621 n1_7271_17279 n1_9521_17279 1.285714e+01
R3622 n1_11771_17279 n1_14021_17279 1.285714e+01
R3623 n1_14021_17279 n1_16271_17279 1.285714e+01
R3624 n1_16271_17279 n1_18521_17279 1.285714e+01
R3625 n1_18521_17279 n1_20771_17279 1.285714e+01
R3626 n1_521_17312 n1_2771_17312 1.285714e+01
R3627 n1_2771_17312 n1_5021_17312 1.285714e+01
R3628 n1_5021_17312 n1_7271_17312 1.285714e+01
R3629 n1_7271_17312 n1_9521_17312 1.285714e+01
R3630 n1_11771_17312 n1_14021_17312 1.285714e+01
R3631 n1_14021_17312 n1_16271_17312 1.285714e+01
R3632 n1_16271_17312 n1_18521_17312 1.285714e+01
R3633 n1_18521_17312 n1_20771_17312 1.285714e+01
R3634 n1_333_17495 n1_521_17495 1.074286e+00
R3635 n1_521_17495 n1_2583_17495 1.178286e+01
R3636 n1_2583_17495 n1_2771_17495 1.074286e+00
R3637 n1_2771_17495 n1_4833_17495 1.178286e+01
R3638 n1_4833_17495 n1_5021_17495 1.074286e+00
R3639 n1_5021_17495 n1_7083_17495 1.178286e+01
R3640 n1_7083_17495 n1_7271_17495 1.074286e+00
R3641 n1_7271_17495 n1_9333_17495 1.178286e+01
R3642 n1_9333_17495 n1_9521_17495 1.074286e+00
R3643 n1_11583_17495 n1_11771_17495 1.074286e+00
R3644 n1_11771_17495 n1_13833_17495 1.178286e+01
R3645 n1_13833_17495 n1_14021_17495 1.074286e+00
R3646 n1_14021_17495 n1_16083_17495 1.178286e+01
R3647 n1_16083_17495 n1_16271_17495 1.074286e+00
R3648 n1_16271_17495 n1_18333_17495 1.178286e+01
R3649 n1_18333_17495 n1_18521_17495 1.074286e+00
R3650 n1_18521_17495 n1_20583_17495 1.178286e+01
R3651 n1_20583_17495 n1_20771_17495 1.074286e+00
R3652 n1_333_17528 n1_521_17528 1.074286e+00
R3653 n1_521_17528 n1_2583_17528 1.178286e+01
R3654 n1_2583_17528 n1_2771_17528 1.074286e+00
R3655 n1_2771_17528 n1_4833_17528 1.178286e+01
R3656 n1_4833_17528 n1_5021_17528 1.074286e+00
R3657 n1_5021_17528 n1_7083_17528 1.178286e+01
R3658 n1_7083_17528 n1_7271_17528 1.074286e+00
R3659 n1_7271_17528 n1_9333_17528 1.178286e+01
R3660 n1_9333_17528 n1_9521_17528 1.074286e+00
R3661 n1_11583_17528 n1_11771_17528 1.074286e+00
R3662 n1_11771_17528 n1_13833_17528 1.178286e+01
R3663 n1_13833_17528 n1_14021_17528 1.074286e+00
R3664 n1_14021_17528 n1_16083_17528 1.178286e+01
R3665 n1_16083_17528 n1_16271_17528 1.074286e+00
R3666 n1_16271_17528 n1_18333_17528 1.178286e+01
R3667 n1_18333_17528 n1_18521_17528 1.074286e+00
R3668 n1_18521_17528 n1_20583_17528 1.178286e+01
R3669 n1_20583_17528 n1_20771_17528 1.074286e+00
R3670 n1_333_17711 n1_521_17711 1.074286e+00
R3671 n1_521_17711 n1_2583_17711 1.178286e+01
R3672 n1_2583_17711 n1_2771_17711 1.074286e+00
R3673 n1_2771_17711 n1_4833_17711 1.178286e+01
R3674 n1_4833_17711 n1_5021_17711 1.074286e+00
R3675 n1_5021_17711 n1_7083_17711 1.178286e+01
R3676 n1_7083_17711 n1_7271_17711 1.074286e+00
R3677 n1_7271_17711 n1_9333_17711 1.178286e+01
R3678 n1_9333_17711 n1_9521_17711 1.074286e+00
R3679 n1_11583_17711 n1_11771_17711 1.074286e+00
R3680 n1_11771_17711 n1_13833_17711 1.178286e+01
R3681 n1_13833_17711 n1_14021_17711 1.074286e+00
R3682 n1_14021_17711 n1_16083_17711 1.178286e+01
R3683 n1_16083_17711 n1_16271_17711 1.074286e+00
R3684 n1_16271_17711 n1_18333_17711 1.178286e+01
R3685 n1_18333_17711 n1_18521_17711 1.074286e+00
R3686 n1_18521_17711 n1_20583_17711 1.178286e+01
R3687 n1_20583_17711 n1_20771_17711 1.074286e+00
R3688 n1_333_17744 n1_521_17744 1.074286e+00
R3689 n1_521_17744 n1_2583_17744 1.178286e+01
R3690 n1_2583_17744 n1_2771_17744 1.074286e+00
R3691 n1_2771_17744 n1_4833_17744 1.178286e+01
R3692 n1_4833_17744 n1_5021_17744 1.074286e+00
R3693 n1_5021_17744 n1_7083_17744 1.178286e+01
R3694 n1_7083_17744 n1_7271_17744 1.074286e+00
R3695 n1_7271_17744 n1_9333_17744 1.178286e+01
R3696 n1_9333_17744 n1_9521_17744 1.074286e+00
R3697 n1_11583_17744 n1_11771_17744 1.074286e+00
R3698 n1_11771_17744 n1_13833_17744 1.178286e+01
R3699 n1_13833_17744 n1_14021_17744 1.074286e+00
R3700 n1_14021_17744 n1_16083_17744 1.178286e+01
R3701 n1_16083_17744 n1_16271_17744 1.074286e+00
R3702 n1_16271_17744 n1_18333_17744 1.178286e+01
R3703 n1_18333_17744 n1_18521_17744 1.074286e+00
R3704 n1_18521_17744 n1_20583_17744 1.178286e+01
R3705 n1_20583_17744 n1_20771_17744 1.074286e+00
R3706 n1_333_17927 n1_521_17927 1.074286e+00
R3707 n1_521_17927 n1_2583_17927 1.178286e+01
R3708 n1_2583_17927 n1_2771_17927 1.074286e+00
R3709 n1_2771_17927 n1_4833_17927 1.178286e+01
R3710 n1_4833_17927 n1_5021_17927 1.074286e+00
R3711 n1_5021_17927 n1_7083_17927 1.178286e+01
R3712 n1_7083_17927 n1_7271_17927 1.074286e+00
R3713 n1_7271_17927 n1_9333_17927 1.178286e+01
R3714 n1_9333_17927 n1_9521_17927 1.074286e+00
R3715 n1_11583_17927 n1_11771_17927 1.074286e+00
R3716 n1_11771_17927 n1_13833_17927 1.178286e+01
R3717 n1_13833_17927 n1_14021_17927 1.074286e+00
R3718 n1_14021_17927 n1_16083_17927 1.178286e+01
R3719 n1_16083_17927 n1_16271_17927 1.074286e+00
R3720 n1_16271_17927 n1_18333_17927 1.178286e+01
R3721 n1_18333_17927 n1_18521_17927 1.074286e+00
R3722 n1_18521_17927 n1_20583_17927 1.178286e+01
R3723 n1_20583_17927 n1_20771_17927 1.074286e+00
R3724 n1_333_17960 n1_521_17960 1.074286e+00
R3725 n1_521_17960 n1_2583_17960 1.178286e+01
R3726 n1_2583_17960 n1_2771_17960 1.074286e+00
R3727 n1_2771_17960 n1_4833_17960 1.178286e+01
R3728 n1_4833_17960 n1_5021_17960 1.074286e+00
R3729 n1_5021_17960 n1_7083_17960 1.178286e+01
R3730 n1_7083_17960 n1_7271_17960 1.074286e+00
R3731 n1_7271_17960 n1_9333_17960 1.178286e+01
R3732 n1_9333_17960 n1_9521_17960 1.074286e+00
R3733 n1_11583_17960 n1_11771_17960 1.074286e+00
R3734 n1_11771_17960 n1_13833_17960 1.178286e+01
R3735 n1_13833_17960 n1_14021_17960 1.074286e+00
R3736 n1_14021_17960 n1_16083_17960 1.178286e+01
R3737 n1_16083_17960 n1_16271_17960 1.074286e+00
R3738 n1_16271_17960 n1_18333_17960 1.178286e+01
R3739 n1_18333_17960 n1_18521_17960 1.074286e+00
R3740 n1_18521_17960 n1_20583_17960 1.178286e+01
R3741 n1_20583_17960 n1_20771_17960 1.074286e+00
R3742 n1_333_18143 n1_521_18143 1.074286e+00
R3743 n1_521_18143 n1_2583_18143 1.178286e+01
R3744 n1_2583_18143 n1_2771_18143 1.074286e+00
R3745 n1_2771_18143 n1_4833_18143 1.178286e+01
R3746 n1_4833_18143 n1_5021_18143 1.074286e+00
R3747 n1_5021_18143 n1_7083_18143 1.178286e+01
R3748 n1_7083_18143 n1_7271_18143 1.074286e+00
R3749 n1_7271_18143 n1_9333_18143 1.178286e+01
R3750 n1_9333_18143 n1_9521_18143 1.074286e+00
R3751 n1_11583_18143 n1_11771_18143 1.074286e+00
R3752 n1_11771_18143 n1_13833_18143 1.178286e+01
R3753 n1_13833_18143 n1_14021_18143 1.074286e+00
R3754 n1_14021_18143 n1_16083_18143 1.178286e+01
R3755 n1_16083_18143 n1_16271_18143 1.074286e+00
R3756 n1_16271_18143 n1_18333_18143 1.178286e+01
R3757 n1_18333_18143 n1_18521_18143 1.074286e+00
R3758 n1_18521_18143 n1_20583_18143 1.178286e+01
R3759 n1_20583_18143 n1_20771_18143 1.074286e+00
R3760 n1_333_18176 n1_521_18176 1.074286e+00
R3761 n1_521_18176 n1_2583_18176 1.178286e+01
R3762 n1_2583_18176 n1_2771_18176 1.074286e+00
R3763 n1_2771_18176 n1_4833_18176 1.178286e+01
R3764 n1_4833_18176 n1_5021_18176 1.074286e+00
R3765 n1_5021_18176 n1_7083_18176 1.178286e+01
R3766 n1_7083_18176 n1_7271_18176 1.074286e+00
R3767 n1_7271_18176 n1_9333_18176 1.178286e+01
R3768 n1_9333_18176 n1_9521_18176 1.074286e+00
R3769 n1_11583_18176 n1_11771_18176 1.074286e+00
R3770 n1_11771_18176 n1_13833_18176 1.178286e+01
R3771 n1_13833_18176 n1_14021_18176 1.074286e+00
R3772 n1_14021_18176 n1_16083_18176 1.178286e+01
R3773 n1_16083_18176 n1_16271_18176 1.074286e+00
R3774 n1_16271_18176 n1_18333_18176 1.178286e+01
R3775 n1_18333_18176 n1_18521_18176 1.074286e+00
R3776 n1_18521_18176 n1_20583_18176 1.178286e+01
R3777 n1_20583_18176 n1_20771_18176 1.074286e+00
R3778 n1_333_18359 n1_521_18359 1.074286e+00
R3779 n1_521_18359 n1_2583_18359 1.178286e+01
R3780 n1_2583_18359 n1_2771_18359 1.074286e+00
R3781 n1_2771_18359 n1_4833_18359 1.178286e+01
R3782 n1_4833_18359 n1_5021_18359 1.074286e+00
R3783 n1_5021_18359 n1_7083_18359 1.178286e+01
R3784 n1_7083_18359 n1_7271_18359 1.074286e+00
R3785 n1_7271_18359 n1_9333_18359 1.178286e+01
R3786 n1_9333_18359 n1_9521_18359 1.074286e+00
R3787 n1_11583_18359 n1_11771_18359 1.074286e+00
R3788 n1_11771_18359 n1_13833_18359 1.178286e+01
R3789 n1_13833_18359 n1_14021_18359 1.074286e+00
R3790 n1_14021_18359 n1_16083_18359 1.178286e+01
R3791 n1_16083_18359 n1_16271_18359 1.074286e+00
R3792 n1_16271_18359 n1_18333_18359 1.178286e+01
R3793 n1_18333_18359 n1_18521_18359 1.074286e+00
R3794 n1_18521_18359 n1_20583_18359 1.178286e+01
R3795 n1_20583_18359 n1_20771_18359 1.074286e+00
R3796 n1_333_18392 n1_380_18392 2.685714e-01
R3797 n1_380_18392 n1_521_18392 8.057143e-01
R3798 n1_521_18392 n1_2583_18392 1.178286e+01
R3799 n1_2583_18392 n1_2630_18392 2.685714e-01
R3800 n1_2630_18392 n1_2771_18392 8.057143e-01
R3801 n1_2771_18392 n1_4833_18392 1.178286e+01
R3802 n1_4833_18392 n1_4880_18392 2.685714e-01
R3803 n1_4880_18392 n1_5021_18392 8.057143e-01
R3804 n1_5021_18392 n1_7083_18392 1.178286e+01
R3805 n1_7083_18392 n1_7130_18392 2.685714e-01
R3806 n1_7130_18392 n1_7271_18392 8.057143e-01
R3807 n1_7271_18392 n1_9333_18392 1.178286e+01
R3808 n1_9333_18392 n1_9380_18392 2.685714e-01
R3809 n1_9380_18392 n1_9521_18392 8.057143e-01
R3810 n1_11583_18392 n1_11630_18392 2.685714e-01
R3811 n1_11630_18392 n1_11771_18392 8.057143e-01
R3812 n1_11771_18392 n1_13833_18392 1.178286e+01
R3813 n1_13833_18392 n1_13880_18392 2.685714e-01
R3814 n1_13880_18392 n1_14021_18392 8.057143e-01
R3815 n1_14021_18392 n1_16083_18392 1.178286e+01
R3816 n1_16083_18392 n1_16130_18392 2.685714e-01
R3817 n1_16130_18392 n1_16271_18392 8.057143e-01
R3818 n1_16271_18392 n1_18333_18392 1.178286e+01
R3819 n1_18333_18392 n1_18380_18392 2.685714e-01
R3820 n1_18380_18392 n1_18521_18392 8.057143e-01
R3821 n1_18521_18392 n1_20583_18392 1.178286e+01
R3822 n1_20583_18392 n1_20630_18392 2.685714e-01
R3823 n1_20630_18392 n1_20771_18392 8.057143e-01
R3824 n1_333_18575 n1_521_18575 1.074286e+00
R3825 n1_521_18575 n1_2400_18575 1.073714e+01
R3826 n1_2400_18575 n1_2583_18575 1.045714e+00
R3827 n1_2583_18575 n1_2771_18575 1.074286e+00
R3828 n1_2771_18575 n1_2864_18575 5.314286e-01
R3829 n1_2864_18575 n1_4650_18575 1.020571e+01
R3830 n1_4650_18575 n1_4833_18575 1.045714e+00
R3831 n1_4833_18575 n1_5021_18575 1.074286e+00
R3832 n1_5021_18575 n1_5114_18575 5.314286e-01
R3833 n1_5114_18575 n1_6900_18575 1.020571e+01
R3834 n1_6900_18575 n1_7083_18575 1.045714e+00
R3835 n1_7083_18575 n1_7271_18575 1.074286e+00
R3836 n1_7271_18575 n1_7364_18575 5.314286e-01
R3837 n1_7364_18575 n1_9150_18575 1.020571e+01
R3838 n1_9150_18575 n1_9333_18575 1.045714e+00
R3839 n1_9333_18575 n1_9521_18575 1.074286e+00
R3840 n1_9521_18575 n1_9614_18575 5.314286e-01
R3841 n1_11400_18575 n1_11583_18575 1.045714e+00
R3842 n1_11583_18575 n1_11771_18575 1.074286e+00
R3843 n1_11771_18575 n1_11864_18575 5.314286e-01
R3844 n1_11864_18575 n1_13650_18575 1.020571e+01
R3845 n1_13650_18575 n1_13833_18575 1.045714e+00
R3846 n1_13833_18575 n1_14021_18575 1.074286e+00
R3847 n1_14021_18575 n1_14114_18575 5.314286e-01
R3848 n1_14114_18575 n1_15900_18575 1.020571e+01
R3849 n1_15900_18575 n1_16083_18575 1.045714e+00
R3850 n1_16083_18575 n1_16271_18575 1.074286e+00
R3851 n1_16271_18575 n1_16364_18575 5.314286e-01
R3852 n1_16364_18575 n1_18150_18575 1.020571e+01
R3853 n1_18150_18575 n1_18333_18575 1.045714e+00
R3854 n1_18333_18575 n1_18521_18575 1.074286e+00
R3855 n1_18521_18575 n1_18614_18575 5.314286e-01
R3856 n1_18614_18575 n1_20583_18575 1.125143e+01
R3857 n1_20583_18575 n1_20771_18575 1.074286e+00
R3858 n1_333_18608 n1_521_18608 1.074286e+00
R3859 n1_521_18608 n1_2400_18608 1.073714e+01
R3860 n1_2400_18608 n1_2583_18608 1.045714e+00
R3861 n1_2583_18608 n1_2771_18608 1.074286e+00
R3862 n1_2771_18608 n1_2864_18608 5.314286e-01
R3863 n1_2864_18608 n1_4650_18608 1.020571e+01
R3864 n1_4650_18608 n1_4833_18608 1.045714e+00
R3865 n1_4833_18608 n1_5021_18608 1.074286e+00
R3866 n1_5021_18608 n1_5114_18608 5.314286e-01
R3867 n1_5114_18608 n1_6900_18608 1.020571e+01
R3868 n1_6900_18608 n1_7083_18608 1.045714e+00
R3869 n1_7083_18608 n1_7271_18608 1.074286e+00
R3870 n1_7271_18608 n1_7364_18608 5.314286e-01
R3871 n1_7364_18608 n1_9150_18608 1.020571e+01
R3872 n1_9150_18608 n1_9333_18608 1.045714e+00
R3873 n1_9333_18608 n1_9521_18608 1.074286e+00
R3874 n1_9521_18608 n1_9614_18608 5.314286e-01
R3875 n1_11400_18608 n1_11583_18608 1.045714e+00
R3876 n1_11583_18608 n1_11771_18608 1.074286e+00
R3877 n1_11771_18608 n1_11864_18608 5.314286e-01
R3878 n1_11864_18608 n1_13650_18608 1.020571e+01
R3879 n1_13650_18608 n1_13833_18608 1.045714e+00
R3880 n1_13833_18608 n1_14021_18608 1.074286e+00
R3881 n1_14021_18608 n1_14114_18608 5.314286e-01
R3882 n1_14114_18608 n1_15900_18608 1.020571e+01
R3883 n1_15900_18608 n1_16083_18608 1.045714e+00
R3884 n1_16083_18608 n1_16271_18608 1.074286e+00
R3885 n1_16271_18608 n1_16364_18608 5.314286e-01
R3886 n1_16364_18608 n1_18150_18608 1.020571e+01
R3887 n1_18150_18608 n1_18333_18608 1.045714e+00
R3888 n1_18333_18608 n1_18521_18608 1.074286e+00
R3889 n1_18521_18608 n1_18614_18608 5.314286e-01
R3890 n1_18614_18608 n1_20583_18608 1.125143e+01
R3891 n1_20583_18608 n1_20771_18608 1.074286e+00
R3892 n1_333_18791 n1_521_18791 1.074286e+00
R3893 n1_521_18791 n1_2400_18791 1.073714e+01
R3894 n1_2400_18791 n1_2583_18791 1.045714e+00
R3895 n1_2583_18791 n1_2771_18791 1.074286e+00
R3896 n1_2771_18791 n1_2864_18791 5.314286e-01
R3897 n1_2864_18791 n1_4650_18791 1.020571e+01
R3898 n1_4650_18791 n1_4833_18791 1.045714e+00
R3899 n1_4833_18791 n1_5021_18791 1.074286e+00
R3900 n1_5021_18791 n1_5114_18791 5.314286e-01
R3901 n1_5114_18791 n1_6900_18791 1.020571e+01
R3902 n1_6900_18791 n1_7083_18791 1.045714e+00
R3903 n1_7083_18791 n1_7271_18791 1.074286e+00
R3904 n1_7271_18791 n1_7364_18791 5.314286e-01
R3905 n1_7364_18791 n1_9150_18791 1.020571e+01
R3906 n1_9150_18791 n1_9333_18791 1.045714e+00
R3907 n1_9333_18791 n1_9521_18791 1.074286e+00
R3908 n1_9521_18791 n1_9614_18791 5.314286e-01
R3909 n1_11400_18791 n1_11583_18791 1.045714e+00
R3910 n1_11583_18791 n1_11771_18791 1.074286e+00
R3911 n1_11771_18791 n1_11864_18791 5.314286e-01
R3912 n1_11864_18791 n1_13650_18791 1.020571e+01
R3913 n1_13650_18791 n1_13833_18791 1.045714e+00
R3914 n1_13833_18791 n1_14021_18791 1.074286e+00
R3915 n1_14021_18791 n1_14114_18791 5.314286e-01
R3916 n1_14114_18791 n1_15900_18791 1.020571e+01
R3917 n1_15900_18791 n1_16083_18791 1.045714e+00
R3918 n1_16083_18791 n1_16271_18791 1.074286e+00
R3919 n1_16271_18791 n1_16364_18791 5.314286e-01
R3920 n1_16364_18791 n1_18150_18791 1.020571e+01
R3921 n1_18150_18791 n1_18333_18791 1.045714e+00
R3922 n1_18333_18791 n1_18521_18791 1.074286e+00
R3923 n1_18521_18791 n1_18614_18791 5.314286e-01
R3924 n1_18614_18791 n1_20583_18791 1.125143e+01
R3925 n1_20583_18791 n1_20771_18791 1.074286e+00
R3926 n1_333_18824 n1_521_18824 1.074286e+00
R3927 n1_521_18824 n1_2400_18824 1.073714e+01
R3928 n1_2400_18824 n1_2583_18824 1.045714e+00
R3929 n1_2583_18824 n1_2771_18824 1.074286e+00
R3930 n1_2771_18824 n1_2864_18824 5.314286e-01
R3931 n1_2864_18824 n1_4650_18824 1.020571e+01
R3932 n1_4650_18824 n1_4833_18824 1.045714e+00
R3933 n1_4833_18824 n1_5021_18824 1.074286e+00
R3934 n1_5021_18824 n1_5114_18824 5.314286e-01
R3935 n1_5114_18824 n1_6900_18824 1.020571e+01
R3936 n1_6900_18824 n1_7083_18824 1.045714e+00
R3937 n1_7083_18824 n1_7271_18824 1.074286e+00
R3938 n1_7271_18824 n1_7364_18824 5.314286e-01
R3939 n1_7364_18824 n1_9150_18824 1.020571e+01
R3940 n1_9150_18824 n1_9333_18824 1.045714e+00
R3941 n1_9333_18824 n1_9521_18824 1.074286e+00
R3942 n1_9521_18824 n1_9614_18824 5.314286e-01
R3943 n1_11400_18824 n1_11583_18824 1.045714e+00
R3944 n1_11583_18824 n1_11771_18824 1.074286e+00
R3945 n1_11771_18824 n1_11864_18824 5.314286e-01
R3946 n1_11864_18824 n1_13650_18824 1.020571e+01
R3947 n1_13650_18824 n1_13833_18824 1.045714e+00
R3948 n1_13833_18824 n1_14021_18824 1.074286e+00
R3949 n1_14021_18824 n1_14114_18824 5.314286e-01
R3950 n1_14114_18824 n1_15900_18824 1.020571e+01
R3951 n1_15900_18824 n1_16083_18824 1.045714e+00
R3952 n1_16083_18824 n1_16271_18824 1.074286e+00
R3953 n1_16271_18824 n1_16364_18824 5.314286e-01
R3954 n1_16364_18824 n1_18150_18824 1.020571e+01
R3955 n1_18150_18824 n1_18333_18824 1.045714e+00
R3956 n1_18333_18824 n1_18521_18824 1.074286e+00
R3957 n1_18521_18824 n1_18614_18824 5.314286e-01
R3958 n1_18614_18824 n1_20583_18824 1.125143e+01
R3959 n1_20583_18824 n1_20771_18824 1.074286e+00
R3960 n1_333_19007 n1_521_19007 1.074286e+00
R3961 n1_521_19007 n1_2400_19007 1.073714e+01
R3962 n1_2400_19007 n1_2583_19007 1.045714e+00
R3963 n1_2583_19007 n1_2771_19007 1.074286e+00
R3964 n1_2771_19007 n1_2864_19007 5.314286e-01
R3965 n1_2864_19007 n1_4650_19007 1.020571e+01
R3966 n1_4650_19007 n1_4833_19007 1.045714e+00
R3967 n1_4833_19007 n1_5021_19007 1.074286e+00
R3968 n1_5021_19007 n1_5114_19007 5.314286e-01
R3969 n1_5114_19007 n1_6900_19007 1.020571e+01
R3970 n1_6900_19007 n1_7083_19007 1.045714e+00
R3971 n1_7083_19007 n1_7271_19007 1.074286e+00
R3972 n1_7271_19007 n1_7364_19007 5.314286e-01
R3973 n1_7364_19007 n1_9150_19007 1.020571e+01
R3974 n1_9150_19007 n1_9333_19007 1.045714e+00
R3975 n1_9333_19007 n1_9521_19007 1.074286e+00
R3976 n1_9521_19007 n1_9614_19007 5.314286e-01
R3977 n1_11400_19007 n1_11583_19007 1.045714e+00
R3978 n1_11583_19007 n1_11771_19007 1.074286e+00
R3979 n1_11771_19007 n1_11864_19007 5.314286e-01
R3980 n1_11864_19007 n1_13650_19007 1.020571e+01
R3981 n1_13650_19007 n1_13833_19007 1.045714e+00
R3982 n1_13833_19007 n1_14021_19007 1.074286e+00
R3983 n1_14021_19007 n1_14114_19007 5.314286e-01
R3984 n1_14114_19007 n1_15900_19007 1.020571e+01
R3985 n1_15900_19007 n1_16083_19007 1.045714e+00
R3986 n1_16083_19007 n1_16271_19007 1.074286e+00
R3987 n1_16271_19007 n1_16364_19007 5.314286e-01
R3988 n1_16364_19007 n1_18150_19007 1.020571e+01
R3989 n1_18150_19007 n1_18333_19007 1.045714e+00
R3990 n1_18333_19007 n1_18521_19007 1.074286e+00
R3991 n1_18521_19007 n1_18614_19007 5.314286e-01
R3992 n1_18614_19007 n1_20583_19007 1.125143e+01
R3993 n1_20583_19007 n1_20771_19007 1.074286e+00
R3994 n1_333_19040 n1_521_19040 1.074286e+00
R3995 n1_521_19040 n1_2400_19040 1.073714e+01
R3996 n1_2400_19040 n1_2583_19040 1.045714e+00
R3997 n1_2583_19040 n1_2771_19040 1.074286e+00
R3998 n1_2771_19040 n1_2864_19040 5.314286e-01
R3999 n1_2864_19040 n1_4650_19040 1.020571e+01
R4000 n1_4650_19040 n1_4833_19040 1.045714e+00
R4001 n1_4833_19040 n1_5021_19040 1.074286e+00
R4002 n1_5021_19040 n1_5114_19040 5.314286e-01
R4003 n1_5114_19040 n1_6900_19040 1.020571e+01
R4004 n1_6900_19040 n1_7083_19040 1.045714e+00
R4005 n1_7083_19040 n1_7271_19040 1.074286e+00
R4006 n1_7271_19040 n1_7364_19040 5.314286e-01
R4007 n1_7364_19040 n1_9150_19040 1.020571e+01
R4008 n1_9150_19040 n1_9333_19040 1.045714e+00
R4009 n1_9333_19040 n1_9521_19040 1.074286e+00
R4010 n1_9521_19040 n1_9614_19040 5.314286e-01
R4011 n1_11400_19040 n1_11583_19040 1.045714e+00
R4012 n1_11583_19040 n1_11771_19040 1.074286e+00
R4013 n1_11771_19040 n1_11864_19040 5.314286e-01
R4014 n1_11864_19040 n1_13650_19040 1.020571e+01
R4015 n1_13650_19040 n1_13833_19040 1.045714e+00
R4016 n1_13833_19040 n1_14021_19040 1.074286e+00
R4017 n1_14021_19040 n1_14114_19040 5.314286e-01
R4018 n1_14114_19040 n1_15900_19040 1.020571e+01
R4019 n1_15900_19040 n1_16083_19040 1.045714e+00
R4020 n1_16083_19040 n1_16271_19040 1.074286e+00
R4021 n1_16271_19040 n1_16364_19040 5.314286e-01
R4022 n1_16364_19040 n1_18150_19040 1.020571e+01
R4023 n1_18150_19040 n1_18333_19040 1.045714e+00
R4024 n1_18333_19040 n1_18521_19040 1.074286e+00
R4025 n1_18521_19040 n1_18614_19040 5.314286e-01
R4026 n1_18614_19040 n1_20583_19040 1.125143e+01
R4027 n1_20583_19040 n1_20771_19040 1.074286e+00
R4028 n1_333_19223 n1_521_19223 1.074286e+00
R4029 n1_521_19223 n1_2400_19223 1.073714e+01
R4030 n1_2400_19223 n1_2583_19223 1.045714e+00
R4031 n1_2583_19223 n1_2771_19223 1.074286e+00
R4032 n1_2771_19223 n1_2864_19223 5.314286e-01
R4033 n1_2864_19223 n1_4650_19223 1.020571e+01
R4034 n1_4650_19223 n1_4833_19223 1.045714e+00
R4035 n1_4833_19223 n1_5021_19223 1.074286e+00
R4036 n1_5021_19223 n1_5114_19223 5.314286e-01
R4037 n1_5114_19223 n1_6900_19223 1.020571e+01
R4038 n1_6900_19223 n1_7083_19223 1.045714e+00
R4039 n1_7083_19223 n1_7271_19223 1.074286e+00
R4040 n1_7271_19223 n1_7364_19223 5.314286e-01
R4041 n1_7364_19223 n1_9150_19223 1.020571e+01
R4042 n1_9150_19223 n1_9333_19223 1.045714e+00
R4043 n1_9333_19223 n1_9521_19223 1.074286e+00
R4044 n1_9521_19223 n1_9614_19223 5.314286e-01
R4045 n1_11400_19223 n1_11583_19223 1.045714e+00
R4046 n1_11583_19223 n1_11771_19223 1.074286e+00
R4047 n1_11771_19223 n1_11864_19223 5.314286e-01
R4048 n1_11864_19223 n1_13650_19223 1.020571e+01
R4049 n1_13650_19223 n1_13833_19223 1.045714e+00
R4050 n1_13833_19223 n1_14021_19223 1.074286e+00
R4051 n1_14021_19223 n1_14114_19223 5.314286e-01
R4052 n1_14114_19223 n1_15900_19223 1.020571e+01
R4053 n1_15900_19223 n1_16083_19223 1.045714e+00
R4054 n1_16083_19223 n1_16271_19223 1.074286e+00
R4055 n1_16271_19223 n1_16364_19223 5.314286e-01
R4056 n1_16364_19223 n1_18150_19223 1.020571e+01
R4057 n1_18150_19223 n1_18333_19223 1.045714e+00
R4058 n1_18333_19223 n1_18521_19223 1.074286e+00
R4059 n1_18521_19223 n1_18614_19223 5.314286e-01
R4060 n1_18614_19223 n1_20583_19223 1.125143e+01
R4061 n1_20583_19223 n1_20771_19223 1.074286e+00
R4062 n1_333_19256 n1_521_19256 1.074286e+00
R4063 n1_521_19256 n1_2400_19256 1.073714e+01
R4064 n1_2400_19256 n1_2583_19256 1.045714e+00
R4065 n1_2583_19256 n1_2771_19256 1.074286e+00
R4066 n1_2771_19256 n1_2864_19256 5.314286e-01
R4067 n1_2864_19256 n1_4650_19256 1.020571e+01
R4068 n1_4650_19256 n1_4833_19256 1.045714e+00
R4069 n1_4833_19256 n1_5021_19256 1.074286e+00
R4070 n1_5021_19256 n1_5114_19256 5.314286e-01
R4071 n1_5114_19256 n1_6900_19256 1.020571e+01
R4072 n1_6900_19256 n1_7083_19256 1.045714e+00
R4073 n1_7083_19256 n1_7271_19256 1.074286e+00
R4074 n1_7271_19256 n1_7364_19256 5.314286e-01
R4075 n1_7364_19256 n1_9150_19256 1.020571e+01
R4076 n1_9150_19256 n1_9333_19256 1.045714e+00
R4077 n1_9333_19256 n1_9521_19256 1.074286e+00
R4078 n1_9521_19256 n1_9614_19256 5.314286e-01
R4079 n1_11400_19256 n1_11583_19256 1.045714e+00
R4080 n1_11583_19256 n1_11771_19256 1.074286e+00
R4081 n1_11771_19256 n1_11864_19256 5.314286e-01
R4082 n1_11864_19256 n1_13650_19256 1.020571e+01
R4083 n1_13650_19256 n1_13833_19256 1.045714e+00
R4084 n1_13833_19256 n1_14021_19256 1.074286e+00
R4085 n1_14021_19256 n1_14114_19256 5.314286e-01
R4086 n1_14114_19256 n1_15900_19256 1.020571e+01
R4087 n1_15900_19256 n1_16083_19256 1.045714e+00
R4088 n1_16083_19256 n1_16271_19256 1.074286e+00
R4089 n1_16271_19256 n1_16364_19256 5.314286e-01
R4090 n1_16364_19256 n1_18150_19256 1.020571e+01
R4091 n1_18150_19256 n1_18333_19256 1.045714e+00
R4092 n1_18333_19256 n1_18521_19256 1.074286e+00
R4093 n1_18521_19256 n1_18614_19256 5.314286e-01
R4094 n1_18614_19256 n1_20583_19256 1.125143e+01
R4095 n1_20583_19256 n1_20771_19256 1.074286e+00
R4096 n1_333_19439 n1_521_19439 1.074286e+00
R4097 n1_521_19439 n1_2400_19439 1.073714e+01
R4098 n1_2400_19439 n1_2583_19439 1.045714e+00
R4099 n1_2583_19439 n1_2771_19439 1.074286e+00
R4100 n1_2771_19439 n1_2864_19439 5.314286e-01
R4101 n1_2864_19439 n1_4650_19439 1.020571e+01
R4102 n1_4650_19439 n1_4833_19439 1.045714e+00
R4103 n1_4833_19439 n1_5021_19439 1.074286e+00
R4104 n1_5021_19439 n1_5114_19439 5.314286e-01
R4105 n1_5114_19439 n1_6900_19439 1.020571e+01
R4106 n1_6900_19439 n1_7083_19439 1.045714e+00
R4107 n1_7083_19439 n1_7271_19439 1.074286e+00
R4108 n1_7271_19439 n1_7364_19439 5.314286e-01
R4109 n1_7364_19439 n1_9150_19439 1.020571e+01
R4110 n1_9150_19439 n1_9333_19439 1.045714e+00
R4111 n1_9333_19439 n1_9521_19439 1.074286e+00
R4112 n1_9521_19439 n1_9614_19439 5.314286e-01
R4113 n1_11400_19439 n1_11583_19439 1.045714e+00
R4114 n1_11583_19439 n1_11771_19439 1.074286e+00
R4115 n1_11771_19439 n1_11864_19439 5.314286e-01
R4116 n1_11864_19439 n1_13650_19439 1.020571e+01
R4117 n1_13650_19439 n1_13833_19439 1.045714e+00
R4118 n1_13833_19439 n1_14021_19439 1.074286e+00
R4119 n1_14021_19439 n1_14114_19439 5.314286e-01
R4120 n1_14114_19439 n1_15900_19439 1.020571e+01
R4121 n1_15900_19439 n1_16083_19439 1.045714e+00
R4122 n1_16083_19439 n1_16271_19439 1.074286e+00
R4123 n1_16271_19439 n1_16364_19439 5.314286e-01
R4124 n1_16364_19439 n1_18150_19439 1.020571e+01
R4125 n1_18150_19439 n1_18333_19439 1.045714e+00
R4126 n1_18333_19439 n1_18521_19439 1.074286e+00
R4127 n1_18521_19439 n1_18614_19439 5.314286e-01
R4128 n1_18614_19439 n1_20583_19439 1.125143e+01
R4129 n1_20583_19439 n1_20771_19439 1.074286e+00
R4130 n1_333_19472 n1_521_19472 1.074286e+00
R4131 n1_521_19472 n1_2400_19472 1.073714e+01
R4132 n1_2400_19472 n1_2583_19472 1.045714e+00
R4133 n1_2583_19472 n1_2771_19472 1.074286e+00
R4134 n1_2771_19472 n1_2864_19472 5.314286e-01
R4135 n1_2864_19472 n1_4650_19472 1.020571e+01
R4136 n1_4650_19472 n1_4833_19472 1.045714e+00
R4137 n1_4833_19472 n1_5021_19472 1.074286e+00
R4138 n1_5021_19472 n1_5114_19472 5.314286e-01
R4139 n1_5114_19472 n1_6900_19472 1.020571e+01
R4140 n1_6900_19472 n1_7083_19472 1.045714e+00
R4141 n1_7083_19472 n1_7271_19472 1.074286e+00
R4142 n1_7271_19472 n1_7364_19472 5.314286e-01
R4143 n1_7364_19472 n1_9150_19472 1.020571e+01
R4144 n1_9150_19472 n1_9333_19472 1.045714e+00
R4145 n1_9333_19472 n1_9521_19472 1.074286e+00
R4146 n1_9521_19472 n1_9614_19472 5.314286e-01
R4147 n1_11400_19472 n1_11583_19472 1.045714e+00
R4148 n1_11583_19472 n1_11771_19472 1.074286e+00
R4149 n1_11771_19472 n1_11864_19472 5.314286e-01
R4150 n1_11864_19472 n1_13650_19472 1.020571e+01
R4151 n1_13650_19472 n1_13833_19472 1.045714e+00
R4152 n1_13833_19472 n1_14021_19472 1.074286e+00
R4153 n1_14021_19472 n1_14114_19472 5.314286e-01
R4154 n1_14114_19472 n1_15900_19472 1.020571e+01
R4155 n1_15900_19472 n1_16083_19472 1.045714e+00
R4156 n1_16083_19472 n1_16271_19472 1.074286e+00
R4157 n1_16271_19472 n1_16364_19472 5.314286e-01
R4158 n1_16364_19472 n1_18150_19472 1.020571e+01
R4159 n1_18150_19472 n1_18333_19472 1.045714e+00
R4160 n1_18333_19472 n1_18521_19472 1.074286e+00
R4161 n1_18521_19472 n1_18614_19472 5.314286e-01
R4162 n1_18614_19472 n1_20583_19472 1.125143e+01
R4163 n1_20583_19472 n1_20771_19472 1.074286e+00
R4164 n1_521_19655 n1_2400_19655 1.073714e+01
R4165 n1_2400_19655 n1_2771_19655 2.120000e+00
R4166 n1_2771_19655 n1_2864_19655 5.314286e-01
R4167 n1_2864_19655 n1_4650_19655 1.020571e+01
R4168 n1_4650_19655 n1_5021_19655 2.120000e+00
R4169 n1_5021_19655 n1_5114_19655 5.314286e-01
R4170 n1_5114_19655 n1_6900_19655 1.020571e+01
R4171 n1_6900_19655 n1_7271_19655 2.120000e+00
R4172 n1_7271_19655 n1_7364_19655 5.314286e-01
R4173 n1_7364_19655 n1_9150_19655 1.020571e+01
R4174 n1_9150_19655 n1_9521_19655 2.120000e+00
R4175 n1_9521_19655 n1_9614_19655 5.314286e-01
R4176 n1_11400_19655 n1_11771_19655 2.120000e+00
R4177 n1_11771_19655 n1_11864_19655 5.314286e-01
R4178 n1_11864_19655 n1_13650_19655 1.020571e+01
R4179 n1_13650_19655 n1_14021_19655 2.120000e+00
R4180 n1_14021_19655 n1_14114_19655 5.314286e-01
R4181 n1_14114_19655 n1_15900_19655 1.020571e+01
R4182 n1_15900_19655 n1_16271_19655 2.120000e+00
R4183 n1_16271_19655 n1_16364_19655 5.314286e-01
R4184 n1_16364_19655 n1_18150_19655 1.020571e+01
R4185 n1_18150_19655 n1_18521_19655 2.120000e+00
R4186 n1_18521_19655 n1_18614_19655 5.314286e-01
R4187 n1_18614_19655 n1_20771_19655 1.232571e+01
R4188 n1_521_19688 n1_2400_19688 1.073714e+01
R4189 n1_2400_19688 n1_2771_19688 2.120000e+00
R4190 n1_2771_19688 n1_2864_19688 5.314286e-01
R4191 n1_2864_19688 n1_4650_19688 1.020571e+01
R4192 n1_4650_19688 n1_5021_19688 2.120000e+00
R4193 n1_5021_19688 n1_5114_19688 5.314286e-01
R4194 n1_5114_19688 n1_6900_19688 1.020571e+01
R4195 n1_6900_19688 n1_7271_19688 2.120000e+00
R4196 n1_7271_19688 n1_7364_19688 5.314286e-01
R4197 n1_7364_19688 n1_9150_19688 1.020571e+01
R4198 n1_9150_19688 n1_9521_19688 2.120000e+00
R4199 n1_9521_19688 n1_9614_19688 5.314286e-01
R4200 n1_11400_19688 n1_11771_19688 2.120000e+00
R4201 n1_11771_19688 n1_11864_19688 5.314286e-01
R4202 n1_11864_19688 n1_13650_19688 1.020571e+01
R4203 n1_13650_19688 n1_14021_19688 2.120000e+00
R4204 n1_14021_19688 n1_14114_19688 5.314286e-01
R4205 n1_14114_19688 n1_15900_19688 1.020571e+01
R4206 n1_15900_19688 n1_16271_19688 2.120000e+00
R4207 n1_16271_19688 n1_16364_19688 5.314286e-01
R4208 n1_16364_19688 n1_18150_19688 1.020571e+01
R4209 n1_18150_19688 n1_18521_19688 2.120000e+00
R4210 n1_18521_19688 n1_18614_19688 5.314286e-01
R4211 n1_18614_19688 n1_20771_19688 1.232571e+01
R4212 n1_333_19871 n1_521_19871 1.074286e+00
R4213 n1_521_19871 n1_2400_19871 1.073714e+01
R4214 n1_2400_19871 n1_2583_19871 1.045714e+00
R4215 n1_2583_19871 n1_2771_19871 1.074286e+00
R4216 n1_2771_19871 n1_2864_19871 5.314286e-01
R4217 n1_2864_19871 n1_4650_19871 1.020571e+01
R4218 n1_4650_19871 n1_4833_19871 1.045714e+00
R4219 n1_4833_19871 n1_5021_19871 1.074286e+00
R4220 n1_5021_19871 n1_5114_19871 5.314286e-01
R4221 n1_5114_19871 n1_6900_19871 1.020571e+01
R4222 n1_6900_19871 n1_7083_19871 1.045714e+00
R4223 n1_7083_19871 n1_7271_19871 1.074286e+00
R4224 n1_7271_19871 n1_7364_19871 5.314286e-01
R4225 n1_7364_19871 n1_9150_19871 1.020571e+01
R4226 n1_9150_19871 n1_9333_19871 1.045714e+00
R4227 n1_9333_19871 n1_9521_19871 1.074286e+00
R4228 n1_9521_19871 n1_9614_19871 5.314286e-01
R4229 n1_11400_19871 n1_11583_19871 1.045714e+00
R4230 n1_11583_19871 n1_11771_19871 1.074286e+00
R4231 n1_11771_19871 n1_11864_19871 5.314286e-01
R4232 n1_11864_19871 n1_13650_19871 1.020571e+01
R4233 n1_13650_19871 n1_13833_19871 1.045714e+00
R4234 n1_13833_19871 n1_14021_19871 1.074286e+00
R4235 n1_14021_19871 n1_14114_19871 5.314286e-01
R4236 n1_14114_19871 n1_15900_19871 1.020571e+01
R4237 n1_15900_19871 n1_16083_19871 1.045714e+00
R4238 n1_16083_19871 n1_16271_19871 1.074286e+00
R4239 n1_16271_19871 n1_16364_19871 5.314286e-01
R4240 n1_16364_19871 n1_18150_19871 1.020571e+01
R4241 n1_18150_19871 n1_18333_19871 1.045714e+00
R4242 n1_18333_19871 n1_18521_19871 1.074286e+00
R4243 n1_18521_19871 n1_18614_19871 5.314286e-01
R4244 n1_18614_19871 n1_20583_19871 1.125143e+01
R4245 n1_20583_19871 n1_20771_19871 1.074286e+00
R4246 n1_333_19904 n1_521_19904 1.074286e+00
R4247 n1_521_19904 n1_2400_19904 1.073714e+01
R4248 n1_2400_19904 n1_2583_19904 1.045714e+00
R4249 n1_2583_19904 n1_2771_19904 1.074286e+00
R4250 n1_2771_19904 n1_2864_19904 5.314286e-01
R4251 n1_2864_19904 n1_4650_19904 1.020571e+01
R4252 n1_4650_19904 n1_4833_19904 1.045714e+00
R4253 n1_4833_19904 n1_5021_19904 1.074286e+00
R4254 n1_5021_19904 n1_5114_19904 5.314286e-01
R4255 n1_5114_19904 n1_6900_19904 1.020571e+01
R4256 n1_6900_19904 n1_7083_19904 1.045714e+00
R4257 n1_7083_19904 n1_7271_19904 1.074286e+00
R4258 n1_7271_19904 n1_7364_19904 5.314286e-01
R4259 n1_7364_19904 n1_9150_19904 1.020571e+01
R4260 n1_9150_19904 n1_9333_19904 1.045714e+00
R4261 n1_9333_19904 n1_9521_19904 1.074286e+00
R4262 n1_9521_19904 n1_9614_19904 5.314286e-01
R4263 n1_11400_19904 n1_11583_19904 1.045714e+00
R4264 n1_11583_19904 n1_11771_19904 1.074286e+00
R4265 n1_11771_19904 n1_11864_19904 5.314286e-01
R4266 n1_11864_19904 n1_13650_19904 1.020571e+01
R4267 n1_13650_19904 n1_13833_19904 1.045714e+00
R4268 n1_13833_19904 n1_14021_19904 1.074286e+00
R4269 n1_14021_19904 n1_14114_19904 5.314286e-01
R4270 n1_14114_19904 n1_15900_19904 1.020571e+01
R4271 n1_15900_19904 n1_16083_19904 1.045714e+00
R4272 n1_16083_19904 n1_16271_19904 1.074286e+00
R4273 n1_16271_19904 n1_16364_19904 5.314286e-01
R4274 n1_16364_19904 n1_18150_19904 1.020571e+01
R4275 n1_18150_19904 n1_18333_19904 1.045714e+00
R4276 n1_18333_19904 n1_18521_19904 1.074286e+00
R4277 n1_18521_19904 n1_18614_19904 5.314286e-01
R4278 n1_18614_19904 n1_20583_19904 1.125143e+01
R4279 n1_20583_19904 n1_20771_19904 1.074286e+00
R4280 n1_333_20087 n1_521_20087 1.074286e+00
R4281 n1_521_20087 n1_2400_20087 1.073714e+01
R4282 n1_2400_20087 n1_2583_20087 1.045714e+00
R4283 n1_2583_20087 n1_2771_20087 1.074286e+00
R4284 n1_2771_20087 n1_2864_20087 5.314286e-01
R4285 n1_2864_20087 n1_4650_20087 1.020571e+01
R4286 n1_4650_20087 n1_4833_20087 1.045714e+00
R4287 n1_4833_20087 n1_5021_20087 1.074286e+00
R4288 n1_5021_20087 n1_5114_20087 5.314286e-01
R4289 n1_5114_20087 n1_6900_20087 1.020571e+01
R4290 n1_6900_20087 n1_7083_20087 1.045714e+00
R4291 n1_7083_20087 n1_7271_20087 1.074286e+00
R4292 n1_7271_20087 n1_7364_20087 5.314286e-01
R4293 n1_7364_20087 n1_9150_20087 1.020571e+01
R4294 n1_9150_20087 n1_9333_20087 1.045714e+00
R4295 n1_9333_20087 n1_9521_20087 1.074286e+00
R4296 n1_9521_20087 n1_9614_20087 5.314286e-01
R4297 n1_11400_20087 n1_11583_20087 1.045714e+00
R4298 n1_11583_20087 n1_11771_20087 1.074286e+00
R4299 n1_11771_20087 n1_11864_20087 5.314286e-01
R4300 n1_11864_20087 n1_13650_20087 1.020571e+01
R4301 n1_13650_20087 n1_13833_20087 1.045714e+00
R4302 n1_13833_20087 n1_14021_20087 1.074286e+00
R4303 n1_14021_20087 n1_14114_20087 5.314286e-01
R4304 n1_14114_20087 n1_15900_20087 1.020571e+01
R4305 n1_15900_20087 n1_16083_20087 1.045714e+00
R4306 n1_16083_20087 n1_16271_20087 1.074286e+00
R4307 n1_16271_20087 n1_16364_20087 5.314286e-01
R4308 n1_16364_20087 n1_18150_20087 1.020571e+01
R4309 n1_18150_20087 n1_18333_20087 1.045714e+00
R4310 n1_18333_20087 n1_18521_20087 1.074286e+00
R4311 n1_18521_20087 n1_18614_20087 5.314286e-01
R4312 n1_18614_20087 n1_20583_20087 1.125143e+01
R4313 n1_20583_20087 n1_20771_20087 1.074286e+00
R4314 n1_333_20120 n1_521_20120 1.074286e+00
R4315 n1_521_20120 n1_2400_20120 1.073714e+01
R4316 n1_2400_20120 n1_2583_20120 1.045714e+00
R4317 n1_2583_20120 n1_2771_20120 1.074286e+00
R4318 n1_2771_20120 n1_2864_20120 5.314286e-01
R4319 n1_2864_20120 n1_4650_20120 1.020571e+01
R4320 n1_4650_20120 n1_4833_20120 1.045714e+00
R4321 n1_4833_20120 n1_5021_20120 1.074286e+00
R4322 n1_5021_20120 n1_5114_20120 5.314286e-01
R4323 n1_5114_20120 n1_6900_20120 1.020571e+01
R4324 n1_6900_20120 n1_7083_20120 1.045714e+00
R4325 n1_7083_20120 n1_7271_20120 1.074286e+00
R4326 n1_7271_20120 n1_7364_20120 5.314286e-01
R4327 n1_7364_20120 n1_9150_20120 1.020571e+01
R4328 n1_9150_20120 n1_9333_20120 1.045714e+00
R4329 n1_9333_20120 n1_9521_20120 1.074286e+00
R4330 n1_9521_20120 n1_9614_20120 5.314286e-01
R4331 n1_11400_20120 n1_11583_20120 1.045714e+00
R4332 n1_11583_20120 n1_11771_20120 1.074286e+00
R4333 n1_11771_20120 n1_11864_20120 5.314286e-01
R4334 n1_11864_20120 n1_13650_20120 1.020571e+01
R4335 n1_13650_20120 n1_13833_20120 1.045714e+00
R4336 n1_13833_20120 n1_14021_20120 1.074286e+00
R4337 n1_14021_20120 n1_14114_20120 5.314286e-01
R4338 n1_14114_20120 n1_15900_20120 1.020571e+01
R4339 n1_15900_20120 n1_16083_20120 1.045714e+00
R4340 n1_16083_20120 n1_16271_20120 1.074286e+00
R4341 n1_16271_20120 n1_16364_20120 5.314286e-01
R4342 n1_16364_20120 n1_18150_20120 1.020571e+01
R4343 n1_18150_20120 n1_18333_20120 1.045714e+00
R4344 n1_18333_20120 n1_18521_20120 1.074286e+00
R4345 n1_18521_20120 n1_18614_20120 5.314286e-01
R4346 n1_18614_20120 n1_20583_20120 1.125143e+01
R4347 n1_20583_20120 n1_20771_20120 1.074286e+00
R4348 n1_333_20303 n1_521_20303 1.074286e+00
R4349 n1_521_20303 n1_2400_20303 1.073714e+01
R4350 n1_2400_20303 n1_2583_20303 1.045714e+00
R4351 n1_2583_20303 n1_2771_20303 1.074286e+00
R4352 n1_2771_20303 n1_2864_20303 5.314286e-01
R4353 n1_2864_20303 n1_4650_20303 1.020571e+01
R4354 n1_4650_20303 n1_4833_20303 1.045714e+00
R4355 n1_4833_20303 n1_5021_20303 1.074286e+00
R4356 n1_5021_20303 n1_5114_20303 5.314286e-01
R4357 n1_5114_20303 n1_6900_20303 1.020571e+01
R4358 n1_6900_20303 n1_7083_20303 1.045714e+00
R4359 n1_7083_20303 n1_7271_20303 1.074286e+00
R4360 n1_7271_20303 n1_7364_20303 5.314286e-01
R4361 n1_7364_20303 n1_9150_20303 1.020571e+01
R4362 n1_9150_20303 n1_9333_20303 1.045714e+00
R4363 n1_9333_20303 n1_9521_20303 1.074286e+00
R4364 n1_9521_20303 n1_9614_20303 5.314286e-01
R4365 n1_11400_20303 n1_11583_20303 1.045714e+00
R4366 n1_11583_20303 n1_11771_20303 1.074286e+00
R4367 n1_11771_20303 n1_11864_20303 5.314286e-01
R4368 n1_11864_20303 n1_13650_20303 1.020571e+01
R4369 n1_13650_20303 n1_13833_20303 1.045714e+00
R4370 n1_13833_20303 n1_14021_20303 1.074286e+00
R4371 n1_14021_20303 n1_14114_20303 5.314286e-01
R4372 n1_14114_20303 n1_15900_20303 1.020571e+01
R4373 n1_15900_20303 n1_16083_20303 1.045714e+00
R4374 n1_16083_20303 n1_16271_20303 1.074286e+00
R4375 n1_16271_20303 n1_16364_20303 5.314286e-01
R4376 n1_16364_20303 n1_18150_20303 1.020571e+01
R4377 n1_18150_20303 n1_18333_20303 1.045714e+00
R4378 n1_18333_20303 n1_18521_20303 1.074286e+00
R4379 n1_18521_20303 n1_18614_20303 5.314286e-01
R4380 n1_18614_20303 n1_20583_20303 1.125143e+01
R4381 n1_20583_20303 n1_20771_20303 1.074286e+00
R4382 n1_333_20336 n1_521_20336 1.074286e+00
R4383 n1_521_20336 n1_2400_20336 1.073714e+01
R4384 n1_2400_20336 n1_2583_20336 1.045714e+00
R4385 n1_2583_20336 n1_2771_20336 1.074286e+00
R4386 n1_2771_20336 n1_2864_20336 5.314286e-01
R4387 n1_2864_20336 n1_4650_20336 1.020571e+01
R4388 n1_4650_20336 n1_4833_20336 1.045714e+00
R4389 n1_4833_20336 n1_5021_20336 1.074286e+00
R4390 n1_5021_20336 n1_5114_20336 5.314286e-01
R4391 n1_5114_20336 n1_6900_20336 1.020571e+01
R4392 n1_6900_20336 n1_7083_20336 1.045714e+00
R4393 n1_7083_20336 n1_7271_20336 1.074286e+00
R4394 n1_7271_20336 n1_7364_20336 5.314286e-01
R4395 n1_7364_20336 n1_9150_20336 1.020571e+01
R4396 n1_9150_20336 n1_9333_20336 1.045714e+00
R4397 n1_9333_20336 n1_9521_20336 1.074286e+00
R4398 n1_9521_20336 n1_9614_20336 5.314286e-01
R4399 n1_11400_20336 n1_11583_20336 1.045714e+00
R4400 n1_11583_20336 n1_11771_20336 1.074286e+00
R4401 n1_11771_20336 n1_11864_20336 5.314286e-01
R4402 n1_11864_20336 n1_13650_20336 1.020571e+01
R4403 n1_13650_20336 n1_13833_20336 1.045714e+00
R4404 n1_13833_20336 n1_14021_20336 1.074286e+00
R4405 n1_14021_20336 n1_14114_20336 5.314286e-01
R4406 n1_14114_20336 n1_15900_20336 1.020571e+01
R4407 n1_15900_20336 n1_16083_20336 1.045714e+00
R4408 n1_16083_20336 n1_16271_20336 1.074286e+00
R4409 n1_16271_20336 n1_16364_20336 5.314286e-01
R4410 n1_16364_20336 n1_18150_20336 1.020571e+01
R4411 n1_18150_20336 n1_18333_20336 1.045714e+00
R4412 n1_18333_20336 n1_18521_20336 1.074286e+00
R4413 n1_18521_20336 n1_18614_20336 5.314286e-01
R4414 n1_18614_20336 n1_20583_20336 1.125143e+01
R4415 n1_20583_20336 n1_20771_20336 1.074286e+00
R4416 n1_333_20519 n1_521_20519 1.074286e+00
R4417 n1_521_20519 n1_2400_20519 1.073714e+01
R4418 n1_2400_20519 n1_2583_20519 1.045714e+00
R4419 n1_2583_20519 n1_2771_20519 1.074286e+00
R4420 n1_2771_20519 n1_2864_20519 5.314286e-01
R4421 n1_2864_20519 n1_4650_20519 1.020571e+01
R4422 n1_4650_20519 n1_4833_20519 1.045714e+00
R4423 n1_4833_20519 n1_5021_20519 1.074286e+00
R4424 n1_5021_20519 n1_5114_20519 5.314286e-01
R4425 n1_5114_20519 n1_6900_20519 1.020571e+01
R4426 n1_6900_20519 n1_7083_20519 1.045714e+00
R4427 n1_7083_20519 n1_7271_20519 1.074286e+00
R4428 n1_7271_20519 n1_7364_20519 5.314286e-01
R4429 n1_7364_20519 n1_9150_20519 1.020571e+01
R4430 n1_9150_20519 n1_9333_20519 1.045714e+00
R4431 n1_9333_20519 n1_9521_20519 1.074286e+00
R4432 n1_9521_20519 n1_9614_20519 5.314286e-01
R4433 n1_11400_20519 n1_11583_20519 1.045714e+00
R4434 n1_11583_20519 n1_11771_20519 1.074286e+00
R4435 n1_11771_20519 n1_11864_20519 5.314286e-01
R4436 n1_11864_20519 n1_13650_20519 1.020571e+01
R4437 n1_13650_20519 n1_13833_20519 1.045714e+00
R4438 n1_13833_20519 n1_14021_20519 1.074286e+00
R4439 n1_14021_20519 n1_14114_20519 5.314286e-01
R4440 n1_14114_20519 n1_15900_20519 1.020571e+01
R4441 n1_15900_20519 n1_16083_20519 1.045714e+00
R4442 n1_16083_20519 n1_16271_20519 1.074286e+00
R4443 n1_16271_20519 n1_16364_20519 5.314286e-01
R4444 n1_16364_20519 n1_18150_20519 1.020571e+01
R4445 n1_18150_20519 n1_18333_20519 1.045714e+00
R4446 n1_18333_20519 n1_18521_20519 1.074286e+00
R4447 n1_18521_20519 n1_18614_20519 5.314286e-01
R4448 n1_18614_20519 n1_20583_20519 1.125143e+01
R4449 n1_20583_20519 n1_20771_20519 1.074286e+00
R4450 n1_333_20552 n1_521_20552 1.074286e+00
R4451 n1_521_20552 n1_2400_20552 1.073714e+01
R4452 n1_2400_20552 n1_2583_20552 1.045714e+00
R4453 n1_2583_20552 n1_2771_20552 1.074286e+00
R4454 n1_2771_20552 n1_2864_20552 5.314286e-01
R4455 n1_2864_20552 n1_4650_20552 1.020571e+01
R4456 n1_4650_20552 n1_4833_20552 1.045714e+00
R4457 n1_4833_20552 n1_5021_20552 1.074286e+00
R4458 n1_5021_20552 n1_5114_20552 5.314286e-01
R4459 n1_5114_20552 n1_6900_20552 1.020571e+01
R4460 n1_6900_20552 n1_7083_20552 1.045714e+00
R4461 n1_7083_20552 n1_7271_20552 1.074286e+00
R4462 n1_7271_20552 n1_7364_20552 5.314286e-01
R4463 n1_7364_20552 n1_9150_20552 1.020571e+01
R4464 n1_9150_20552 n1_9333_20552 1.045714e+00
R4465 n1_9333_20552 n1_9521_20552 1.074286e+00
R4466 n1_9521_20552 n1_9614_20552 5.314286e-01
R4467 n1_11400_20552 n1_11583_20552 1.045714e+00
R4468 n1_11583_20552 n1_11771_20552 1.074286e+00
R4469 n1_11771_20552 n1_11864_20552 5.314286e-01
R4470 n1_11864_20552 n1_13650_20552 1.020571e+01
R4471 n1_13650_20552 n1_13833_20552 1.045714e+00
R4472 n1_13833_20552 n1_14021_20552 1.074286e+00
R4473 n1_14021_20552 n1_14114_20552 5.314286e-01
R4474 n1_14114_20552 n1_15900_20552 1.020571e+01
R4475 n1_15900_20552 n1_16083_20552 1.045714e+00
R4476 n1_16083_20552 n1_16271_20552 1.074286e+00
R4477 n1_16271_20552 n1_16364_20552 5.314286e-01
R4478 n1_16364_20552 n1_18150_20552 1.020571e+01
R4479 n1_18150_20552 n1_18333_20552 1.045714e+00
R4480 n1_18333_20552 n1_18521_20552 1.074286e+00
R4481 n1_18521_20552 n1_18614_20552 5.314286e-01
R4482 n1_18614_20552 n1_20583_20552 1.125143e+01
R4483 n1_20583_20552 n1_20771_20552 1.074286e+00
R4484 n1_333_20735 n1_380_20735 2.685714e-01
R4485 n1_380_20735 n1_2400_20735 1.154286e+01
R4486 n1_2400_20735 n1_2583_20735 1.045714e+00
R4487 n1_2583_20735 n1_2630_20735 2.685714e-01
R4488 n1_2630_20735 n1_2864_20735 1.337143e+00
R4489 n1_2864_20735 n1_4650_20735 1.020571e+01
R4490 n1_4650_20735 n1_4833_20735 1.045714e+00
R4491 n1_4833_20735 n1_4880_20735 2.685714e-01
R4492 n1_4880_20735 n1_5114_20735 1.337143e+00
R4493 n1_5114_20735 n1_6900_20735 1.020571e+01
R4494 n1_6900_20735 n1_7083_20735 1.045714e+00
R4495 n1_7083_20735 n1_7130_20735 2.685714e-01
R4496 n1_7130_20735 n1_7364_20735 1.337143e+00
R4497 n1_7364_20735 n1_9150_20735 1.020571e+01
R4498 n1_9150_20735 n1_9333_20735 1.045714e+00
R4499 n1_9333_20735 n1_9380_20735 2.685714e-01
R4500 n1_9380_20735 n1_9614_20735 1.337143e+00
R4501 n1_11400_20735 n1_11583_20735 1.045714e+00
R4502 n1_11583_20735 n1_11630_20735 2.685714e-01
R4503 n1_11630_20735 n1_11864_20735 1.337143e+00
R4504 n1_11864_20735 n1_13650_20735 1.020571e+01
R4505 n1_13650_20735 n1_13833_20735 1.045714e+00
R4506 n1_13833_20735 n1_13880_20735 2.685714e-01
R4507 n1_13880_20735 n1_14114_20735 1.337143e+00
R4508 n1_14114_20735 n1_15900_20735 1.020571e+01
R4509 n1_15900_20735 n1_16083_20735 1.045714e+00
R4510 n1_16083_20735 n1_16130_20735 2.685714e-01
R4511 n1_16130_20735 n1_16364_20735 1.337143e+00
R4512 n1_16364_20735 n1_18150_20735 1.020571e+01
R4513 n1_18150_20735 n1_18333_20735 1.045714e+00
R4514 n1_18333_20735 n1_18380_20735 2.685714e-01
R4515 n1_18380_20735 n1_18614_20735 1.337143e+00
R4516 n1_18614_20735 n1_20583_20735 1.125143e+01
R4517 n1_20583_20735 n1_20630_20735 2.685714e-01
R4518 n1_333_20768 n1_380_20768 2.685714e-01
R4519 n1_380_20768 n1_521_20768 8.057143e-01
R4520 n1_521_20768 n1_2400_20768 1.073714e+01
R4521 n1_2400_20768 n1_2583_20768 1.045714e+00
R4522 n1_2583_20768 n1_2630_20768 2.685714e-01
R4523 n1_2630_20768 n1_2771_20768 8.057143e-01
R4524 n1_2771_20768 n1_2864_20768 5.314286e-01
R4525 n1_2864_20768 n1_4650_20768 1.020571e+01
R4526 n1_4650_20768 n1_4833_20768 1.045714e+00
R4527 n1_4833_20768 n1_4880_20768 2.685714e-01
R4528 n1_4880_20768 n1_5021_20768 8.057143e-01
R4529 n1_5021_20768 n1_5114_20768 5.314286e-01
R4530 n1_5114_20768 n1_6900_20768 1.020571e+01
R4531 n1_6900_20768 n1_7083_20768 1.045714e+00
R4532 n1_7083_20768 n1_7130_20768 2.685714e-01
R4533 n1_7130_20768 n1_7271_20768 8.057143e-01
R4534 n1_7271_20768 n1_7364_20768 5.314286e-01
R4535 n1_7364_20768 n1_9150_20768 1.020571e+01
R4536 n1_9150_20768 n1_9333_20768 1.045714e+00
R4537 n1_9333_20768 n1_9380_20768 2.685714e-01
R4538 n1_9380_20768 n1_9521_20768 8.057143e-01
R4539 n1_9521_20768 n1_9614_20768 5.314286e-01
R4540 n1_11400_20768 n1_11583_20768 1.045714e+00
R4541 n1_11583_20768 n1_11630_20768 2.685714e-01
R4542 n1_11630_20768 n1_11771_20768 8.057143e-01
R4543 n1_11771_20768 n1_11864_20768 5.314286e-01
R4544 n1_11864_20768 n1_13650_20768 1.020571e+01
R4545 n1_13650_20768 n1_13833_20768 1.045714e+00
R4546 n1_13833_20768 n1_13880_20768 2.685714e-01
R4547 n1_13880_20768 n1_14021_20768 8.057143e-01
R4548 n1_14021_20768 n1_14114_20768 5.314286e-01
R4549 n1_14114_20768 n1_15900_20768 1.020571e+01
R4550 n1_15900_20768 n1_16083_20768 1.045714e+00
R4551 n1_16083_20768 n1_16130_20768 2.685714e-01
R4552 n1_16130_20768 n1_16271_20768 8.057143e-01
R4553 n1_16271_20768 n1_16364_20768 5.314286e-01
R4554 n1_16364_20768 n1_18150_20768 1.020571e+01
R4555 n1_18150_20768 n1_18333_20768 1.045714e+00
R4556 n1_18333_20768 n1_18380_20768 2.685714e-01
R4557 n1_18380_20768 n1_18521_20768 8.057143e-01
R4558 n1_18521_20768 n1_18614_20768 5.314286e-01
R4559 n1_18614_20768 n1_20583_20768 1.125143e+01
R4560 n1_20583_20768 n1_20630_20768 2.685714e-01
R4561 n1_333_13774 n1_521_13774 1.342857e-01
R4562 n1_333_4486 n1_521_4486 1.342857e-01
R4563 n1_333_18116 n1_521_18116 4.700000e-01
R4564 n1_333_19196 n1_521_19196 4.700000e-01
R4565 n1_333_19412 n1_521_19412 4.700000e-01
R4566 n1_521_215 n1_2400_215 1.073714e+01
R4567 n1_2400_215 n1_2583_215 1.045714e+00
R4568 n1_2583_215 n1_2771_215 1.074286e+00
R4569 n1_2771_215 n1_2864_215 5.314286e-01
R4570 n1_2864_215 n1_4650_215 1.020571e+01
R4571 n1_4650_215 n1_4833_215 1.045714e+00
R4572 n1_4833_215 n1_5021_215 1.074286e+00
R4573 n1_5021_215 n1_5114_215 5.314286e-01
R4574 n1_5114_215 n1_6900_215 1.020571e+01
R4575 n1_6900_215 n1_7083_215 1.045714e+00
R4576 n1_7083_215 n1_7271_215 1.074286e+00
R4577 n1_7271_215 n1_7364_215 5.314286e-01
R4578 n1_7364_215 n1_9150_215 1.020571e+01
R4579 n1_9150_215 n1_9333_215 1.045714e+00
R4580 n1_9333_215 n1_9521_215 1.074286e+00
R4581 n1_9521_215 n1_9614_215 5.314286e-01
R4582 n1_521_248 n1_2400_248 1.073714e+01
R4583 n1_2400_248 n1_2583_248 1.045714e+00
R4584 n1_2583_248 n1_2771_248 1.074286e+00
R4585 n1_2771_248 n1_2864_248 5.314286e-01
R4586 n1_2864_248 n1_4650_248 1.020571e+01
R4587 n1_4650_248 n1_4833_248 1.045714e+00
R4588 n1_4833_248 n1_5021_248 1.074286e+00
R4589 n1_5021_248 n1_5114_248 5.314286e-01
R4590 n1_5114_248 n1_6900_248 1.020571e+01
R4591 n1_6900_248 n1_7083_248 1.045714e+00
R4592 n1_7083_248 n1_7271_248 1.074286e+00
R4593 n1_7271_248 n1_7364_248 5.314286e-01
R4594 n1_7364_248 n1_9150_248 1.020571e+01
R4595 n1_9150_248 n1_9333_248 1.045714e+00
R4596 n1_9333_248 n1_9521_248 1.074286e+00
R4597 n1_9521_248 n1_9614_248 5.314286e-01
R4598 n1_521_20951 n1_2400_20951 1.073714e+01
R4599 n1_2400_20951 n1_2583_20951 1.045714e+00
R4600 n1_2583_20951 n1_2771_20951 1.074286e+00
R4601 n1_2771_20951 n1_2864_20951 5.314286e-01
R4602 n1_2864_20951 n1_4650_20951 1.020571e+01
R4603 n1_4650_20951 n1_4833_20951 1.045714e+00
R4604 n1_4833_20951 n1_5021_20951 1.074286e+00
R4605 n1_5021_20951 n1_5114_20951 5.314286e-01
R4606 n1_5114_20951 n1_6900_20951 1.020571e+01
R4607 n1_6900_20951 n1_7083_20951 1.045714e+00
R4608 n1_7083_20951 n1_7271_20951 1.074286e+00
R4609 n1_7271_20951 n1_7364_20951 5.314286e-01
R4610 n1_7364_20951 n1_9150_20951 1.020571e+01
R4611 n1_9150_20951 n1_9333_20951 1.045714e+00
R4612 n1_9333_20951 n1_9521_20951 1.074286e+00
R4613 n1_9521_20951 n1_9614_20951 5.314286e-01
R4614 n1_11400_20951 n1_11583_20951 1.045714e+00
R4615 n1_11583_20951 n1_11771_20951 1.074286e+00
R4616 n1_11771_20951 n1_11864_20951 5.314286e-01
R4617 n1_11864_20951 n1_13650_20951 1.020571e+01
R4618 n1_13650_20951 n1_13833_20951 1.045714e+00
R4619 n1_13833_20951 n1_14021_20951 1.074286e+00
R4620 n1_14021_20951 n1_14114_20951 5.314286e-01
R4621 n1_14114_20951 n1_15900_20951 1.020571e+01
R4622 n1_15900_20951 n1_16083_20951 1.045714e+00
R4623 n1_16083_20951 n1_16271_20951 1.074286e+00
R4624 n1_16271_20951 n1_16364_20951 5.314286e-01
R4625 n1_16364_20951 n1_18150_20951 1.020571e+01
R4626 n1_18150_20951 n1_18333_20951 1.045714e+00
R4627 n1_18333_20951 n1_18521_20951 1.074286e+00
R4628 n1_18521_20951 n1_18614_20951 5.314286e-01
R4629 n1_18614_20951 n1_20583_20951 1.125143e+01
R4630 n1_521_20984 n1_2400_20984 1.073714e+01
R4631 n1_2400_20984 n1_2583_20984 1.045714e+00
R4632 n1_2583_20984 n1_2771_20984 1.074286e+00
R4633 n1_2771_20984 n1_2864_20984 5.314286e-01
R4634 n1_2864_20984 n1_4650_20984 1.020571e+01
R4635 n1_4650_20984 n1_4833_20984 1.045714e+00
R4636 n1_4833_20984 n1_5021_20984 1.074286e+00
R4637 n1_5021_20984 n1_5114_20984 5.314286e-01
R4638 n1_5114_20984 n1_6900_20984 1.020571e+01
R4639 n1_6900_20984 n1_7083_20984 1.045714e+00
R4640 n1_7083_20984 n1_7271_20984 1.074286e+00
R4641 n1_7271_20984 n1_7364_20984 5.314286e-01
R4642 n1_7364_20984 n1_9150_20984 1.020571e+01
R4643 n1_9150_20984 n1_9333_20984 1.045714e+00
R4644 n1_9333_20984 n1_9521_20984 1.074286e+00
R4645 n1_9521_20984 n1_9614_20984 5.314286e-01
R4646 n1_11400_20984 n1_11583_20984 1.045714e+00
R4647 n1_11583_20984 n1_11771_20984 1.074286e+00
R4648 n1_11771_20984 n1_11864_20984 5.314286e-01
R4649 n1_11864_20984 n1_13650_20984 1.020571e+01
R4650 n1_13650_20984 n1_13833_20984 1.045714e+00
R4651 n1_13833_20984 n1_14021_20984 1.074286e+00
R4652 n1_14021_20984 n1_14114_20984 5.314286e-01
R4653 n1_14114_20984 n1_15900_20984 1.020571e+01
R4654 n1_15900_20984 n1_16083_20984 1.045714e+00
R4655 n1_16083_20984 n1_16271_20984 1.074286e+00
R4656 n1_16271_20984 n1_16364_20984 5.314286e-01
R4657 n1_16364_20984 n1_18150_20984 1.020571e+01
R4658 n1_18150_20984 n1_18333_20984 1.045714e+00
R4659 n1_18333_20984 n1_18521_20984 1.074286e+00
R4660 n1_18521_20984 n1_18614_20984 5.314286e-01
R4661 n1_18614_20984 n1_20583_20984 1.125143e+01
R4662 n1_2583_5446 n1_2771_5446 4.700000e-01
R4663 n1_2771_5446 n1_4833_5446 5.155000e+00
R4664 n1_4833_5446 n1_5021_5446 4.700000e-01
R4665 n1_2583_6549 n1_2771_6549 1.342857e-01
R4666 n1_2771_6549 n1_4833_6549 1.472857e+00
R4667 n1_4833_6549 n1_5021_6549 1.342857e-01
R4668 n1_2583_8902 n1_2771_8902 4.700000e-01
R4669 n1_2771_8902 n1_4833_8902 5.155000e+00
R4670 n1_4833_8902 n1_5021_8902 4.700000e-01
R4671 n1_5021_8902 n1_7083_8902 5.155000e+00
R4672 n1_7083_8902 n1_7271_8902 4.700000e-01
R4673 n1_2583_9982 n1_2771_9982 4.700000e-01
R4674 n1_2771_9982 n1_4833_9982 5.155000e+00
R4675 n1_4833_9982 n1_5021_9982 4.700000e-01
R4676 n1_5021_9982 n1_7083_9982 5.155000e+00
R4677 n1_7083_9982 n1_7271_9982 4.700000e-01
R4678 n1_2583_7822 n1_2771_7822 4.700000e-01
R4679 n1_2771_7822 n1_4833_7822 5.155000e+00
R4680 n1_4833_7822 n1_5021_7822 4.700000e-01
R4681 n1_5021_7822 n1_7083_7822 5.155000e+00
R4682 n1_7083_7822 n1_7271_7822 4.700000e-01
R4683 n1_2583_3428 n1_2771_3428 4.700000e-01
R4684 n1_2583_11182 n1_2771_11182 1.342857e-01
R4685 n1_2583_13558 n1_2771_13558 1.342857e-01
R4686 n1_2583_14660 n1_2771_14660 4.700000e-01
R4687 n1_2583_9022 n1_2771_9022 1.342857e-01
R4688 n1_2583_15524 n1_2771_15524 4.700000e-01
R4689 n1_2583_4508 n1_2771_4508 4.700000e-01
R4690 n1_2583_5588 n1_2771_5588 4.700000e-01
R4691 n1_2583_7964 n1_2771_7964 4.700000e-01
R4692 n1_2583_10124 n1_2771_10124 4.700000e-01
R4693 n1_2583_12284 n1_2771_12284 4.700000e-01
R4694 n1_2583_9044 n1_2771_9044 4.700000e-01
R4695 n1_2583_11204 n1_2771_11204 4.700000e-01
R4696 n1_2583_16798 n1_2771_16798 1.342857e-01
R4697 n1_2583_17684 n1_2771_17684 4.700000e-01
R4698 n1_2583_6646 n1_2771_6646 1.342857e-01
R4699 n1_2583_17036 n1_2771_17036 4.700000e-01
R4700 n1_2583_4076 n1_2771_4076 4.700000e-01
R4701 n1_2583_4270 n1_2771_4270 1.342857e-01
R4702 n1_2583_16582 n1_2771_16582 1.342857e-01
R4703 n1_2583_13990 n1_2630_13990 3.357143e-02
R4704 n1_2630_13990 n1_2771_13990 1.007143e-01
R4705 n1_2583_12262 n1_2771_12262 1.342857e-01
R4706 n1_2583_13796 n1_2771_13796 4.700000e-01
R4707 n1_2583_15740 n1_2771_15740 4.700000e-01
R4708 n1_2583_13580 n1_2771_13580 4.700000e-01
R4709 n1_2583_16820 n1_2771_16820 4.700000e-01
R4710 n1_2583_14206 n1_2771_14206 1.342857e-01
R4711 n1_2583_17662 n1_2771_17662 1.342857e-01
R4712 n1_4833_15524 n1_5021_15524 4.700000e-01
R4713 n1_4833_5588 n1_5021_5588 4.700000e-01
R4714 n1_4833_15740 n1_5021_15740 4.700000e-01
R4715 n1_4833_6646 n1_5021_6646 1.342857e-01
R4716 n1_4833_7964 n1_5021_7964 4.700000e-01
R4717 n1_4833_9044 n1_5021_9044 4.700000e-01
R4718 n1_4833_10124 n1_5021_10124 4.700000e-01
R4719 n1_4833_11204 n1_5021_11204 4.700000e-01
R4720 n1_4833_12284 n1_5021_12284 4.700000e-01
R4721 n1_4833_13580 n1_5021_13580 4.700000e-01
R4722 n1_4833_13990 n1_4880_13990 3.357143e-02
R4723 n1_4833_14206 n1_5021_14206 1.342857e-01
R4724 n1_4650_2132 n1_4833_2132 4.575000e-01
R4725 n1_4833_2132 n1_5021_2132 4.700000e-01
R4726 n1_4833_17036 n1_5021_17036 4.700000e-01
R4727 n1_4833_17684 n1_5021_17684 4.700000e-01
R4728 n1_4833_4292 n1_5021_4292 4.700000e-01
R4729 n1_4833_4508 n1_5021_4508 4.700000e-01
R4730 n1_4650_513 n1_4833_513 4.575000e-01
R4731 n1_4833_513 n1_4880_513 1.175000e-01
R4732 n1_4880_513 n1_5021_513 3.525000e-01
R4733 n1_5021_513 n1_5114_513 2.325000e-01
R4734 n1_4650_945 n1_4833_945 4.575000e-01
R4735 n1_4833_945 n1_5021_945 4.700000e-01
R4736 n1_5021_945 n1_5114_945 2.325000e-01
R4737 n1_4833_4486 n1_5021_4486 1.342857e-01
R4738 n1_4833_16172 n1_4880_16172 1.175000e-01
R4739 n1_4880_16172 n1_5021_16172 3.525000e-01
R4740 n1_4833_18548 n1_4880_18548 1.175000e-01
R4741 n1_4880_18548 n1_5021_18548 3.525000e-01
R4742 n1_5021_18548 n1_5114_18548 2.325000e-01
R4743 n1_4833_9022 n1_5021_9022 1.342857e-01
R4744 n1_4833_11182 n1_5021_11182 1.342857e-01
R4745 n1_4833_1916 n1_5021_1916 4.700000e-01
R4746 n1_5021_1916 n1_5114_1916 2.325000e-01
R4747 n1_4833_2564 n1_5021_2564 4.700000e-01
R4748 n1_5021_2564 n1_5114_2564 2.325000e-01
R4749 n1_4833_2996 n1_5021_2996 4.700000e-01
R4750 n1_4833_3212 n1_5021_3212 4.700000e-01
R4751 n1_4833_3644 n1_5021_3644 4.700000e-01
R4752 n1_4833_17468 n1_5021_17468 4.700000e-01
R4753 n1_4833_18764 n1_5021_18764 4.700000e-01
R4754 n1_5021_18764 n1_5114_18764 2.325000e-01
R4755 n1_4833_18980 n1_5021_18980 4.700000e-01
R4756 n1_5021_18980 n1_5114_18980 2.325000e-01
R4757 n1_4833_19196 n1_5021_19196 4.700000e-01
R4758 n1_5021_19196 n1_5114_19196 2.325000e-01
R4759 n1_5021_19628 n1_5114_19628 2.325000e-01
R4760 n1_7083_7964 n1_7271_7964 4.700000e-01
R4761 n1_7083_13580 n1_7271_13580 4.700000e-01
R4762 n1_7083_9044 n1_7271_9044 4.700000e-01
R4763 n1_7083_10124 n1_7271_10124 4.700000e-01
R4764 n1_7083_11204 n1_7271_11204 4.700000e-01
R4765 n1_7083_12284 n1_7271_12284 4.700000e-01
R4766 n1_6900_383 n1_7083_383 1.307143e-01
R4767 n1_7083_383 n1_7271_383 1.342857e-01
R4768 n1_7271_383 n1_7364_383 6.642857e-02
R4769 n1_7364_383 n1_9150_383 1.275714e+00
R4770 n1_9150_383 n1_9333_383 1.307143e-01
R4771 n1_9333_383 n1_9521_383 1.342857e-01
R4772 n1_9521_383 n1_9614_383 6.642857e-02
R4773 n1_6900_18548 n1_7083_18548 4.575000e-01
R4774 n1_7083_18548 n1_7130_18548 1.175000e-01
R4775 n1_7130_18548 n1_7271_18548 3.525000e-01
R4776 n1_7083_2996 n1_7271_2996 4.700000e-01
R4777 n1_6900_19196 n1_7083_19196 4.575000e-01
R4778 n1_7083_19196 n1_7271_19196 4.700000e-01
R4779 n1_6900_1916 n1_7083_1916 4.575000e-01
R4780 n1_7083_1916 n1_7271_1916 4.700000e-01
R4781 n1_7271_1916 n1_7364_1916 2.325000e-01
R4782 n1_6900_2564 n1_7083_2564 4.575000e-01
R4783 n1_7083_2564 n1_7271_2564 4.700000e-01
R4784 n1_7271_2564 n1_7364_2564 2.325000e-01
R4785 n1_7083_3644 n1_7271_3644 4.700000e-01
R4786 n1_7083_4292 n1_7271_4292 4.700000e-01
R4787 n1_7083_4724 n1_7271_4724 4.700000e-01
R4788 n1_7083_5372 n1_7271_5372 4.700000e-01
R4789 n1_7083_5588 n1_7271_5588 4.700000e-01
R4790 n1_7083_15740 n1_7271_15740 4.700000e-01
R4791 n1_7083_15956 n1_7271_15956 4.700000e-01
R4792 n1_7083_16172 n1_7130_16172 1.175000e-01
R4793 n1_7130_16172 n1_7271_16172 3.525000e-01
R4794 n1_7083_17468 n1_7271_17468 4.700000e-01
R4795 n1_6900_18764 n1_7083_18764 4.575000e-01
R4796 n1_7083_18764 n1_7271_18764 4.700000e-01
R4797 n1_7271_18764 n1_7364_18764 2.325000e-01
R4798 n1_7083_6646 n1_7271_6646 1.342857e-01
R4799 n1_7083_5566 n1_7271_5566 1.342857e-01
R4800 n1_7083_17230 n1_7271_17230 1.342857e-01
R4801 n1_7083_18526 n1_7130_18526 3.357143e-02
R4802 n1_7130_18526 n1_7271_18526 1.007143e-01
R4803 n1_7271_18526 n1_7364_18526 6.642857e-02
R4804 n1_7083_2974 n1_7271_2974 1.342857e-01
R4805 n1_7083_19390 n1_7271_19390 1.342857e-01
R4806 n1_7271_19390 n1_7364_19390 6.642857e-02
R4807 n1_7083_14553 n1_7271_14553 4.700000e-01
R4808 n1_9333_3644 n1_9521_3644 4.700000e-01
R4809 n1_9333_4724 n1_9521_4724 4.700000e-01
R4810 n1_9150_1894 n1_9333_1894 1.307143e-01
R4811 n1_9333_1894 n1_9521_1894 1.342857e-01
R4812 n1_9333_5372 n1_9521_5372 4.700000e-01
R4813 n1_9333_14012 n1_9380_14012 1.175000e-01
R4814 n1_9380_14012 n1_9521_14012 3.525000e-01
R4815 n1_9333_15956 n1_9521_15956 4.700000e-01
R4816 n1_9150_2564 n1_9333_2564 4.575000e-01
R4817 n1_9333_2564 n1_9521_2564 4.700000e-01
R4818 n1_9521_2564 n1_9614_2564 2.325000e-01
R4819 n1_9333_2996 n1_9521_2996 4.700000e-01
R4820 n1_9333_4292 n1_9521_4292 4.700000e-01
R4821 n1_9333_5588 n1_9521_5588 4.700000e-01
R4822 n1_9333_6668 n1_9521_6668 4.700000e-01
R4823 n1_9333_7100 n1_9521_7100 4.700000e-01
R4824 n1_9333_7316 n1_9521_7316 4.700000e-01
R4825 n1_9333_7532 n1_9521_7532 4.700000e-01
R4826 n1_9333_13796 n1_9521_13796 4.700000e-01
R4827 n1_9333_14228 n1_9521_14228 4.700000e-01
R4828 n1_9333_14660 n1_9521_14660 4.700000e-01
R4829 n1_9333_15740 n1_9521_15740 4.700000e-01
R4830 n1_9333_16172 n1_9380_16172 1.175000e-01
R4831 n1_9380_16172 n1_9521_16172 3.525000e-01
R4832 n1_9333_17468 n1_9521_17468 4.700000e-01
R4833 n1_9150_18548 n1_9333_18548 4.575000e-01
R4834 n1_9333_18548 n1_9380_18548 1.175000e-01
R4835 n1_9380_18548 n1_9521_18548 3.525000e-01
R4836 n1_9521_18548 n1_9614_18548 2.325000e-01
R4837 n1_9150_18764 n1_9333_18764 4.575000e-01
R4838 n1_9333_18764 n1_9521_18764 4.700000e-01
R4839 n1_9521_18764 n1_9614_18764 2.325000e-01
R4840 n1_9150_19412 n1_9333_19412 4.575000e-01
R4841 n1_9333_19412 n1_9521_19412 4.700000e-01
R4842 n1_9521_19412 n1_9614_19412 2.325000e-01
R4843 n1_9333_17230 n1_9521_17230 1.342857e-01
R4844 n1_9333_5350 n1_9521_5350 1.342857e-01
R4845 n1_9333_13990 n1_9380_13990 3.357143e-02
R4846 n1_9380_13990 n1_9521_13990 1.007143e-01
R4847 n1_9333_1916 n1_9521_1916 4.700000e-01
R4848 n1_9521_1916 n1_9614_1916 2.325000e-01
R4849 n1_9333_15934 n1_9521_15934 1.342857e-01
R4850 n1_11400_215 n1_11583_215 1.045714e+00
R4851 n1_11583_215 n1_11771_215 1.074286e+00
R4852 n1_11771_215 n1_11864_215 5.314286e-01
R4853 n1_11864_215 n1_13650_215 1.020571e+01
R4854 n1_13650_215 n1_13833_215 1.045714e+00
R4855 n1_13833_215 n1_14021_215 1.074286e+00
R4856 n1_14021_215 n1_14114_215 5.314286e-01
R4857 n1_14114_215 n1_15900_215 1.020571e+01
R4858 n1_15900_215 n1_16083_215 1.045714e+00
R4859 n1_16083_215 n1_16271_215 1.074286e+00
R4860 n1_16271_215 n1_16364_215 5.314286e-01
R4861 n1_16364_215 n1_18150_215 1.020571e+01
R4862 n1_18150_215 n1_18333_215 1.045714e+00
R4863 n1_18333_215 n1_18521_215 1.074286e+00
R4864 n1_18521_215 n1_18614_215 5.314286e-01
R4865 n1_18614_215 n1_20583_215 1.125143e+01
R4866 n1_11400_248 n1_11583_248 1.045714e+00
R4867 n1_11583_248 n1_11771_248 1.074286e+00
R4868 n1_11771_248 n1_11864_248 5.314286e-01
R4869 n1_11864_248 n1_13650_248 1.020571e+01
R4870 n1_13650_248 n1_13833_248 1.045714e+00
R4871 n1_13833_248 n1_14021_248 1.074286e+00
R4872 n1_14021_248 n1_14114_248 5.314286e-01
R4873 n1_14114_248 n1_15900_248 1.020571e+01
R4874 n1_15900_248 n1_16083_248 1.045714e+00
R4875 n1_16083_248 n1_16271_248 1.074286e+00
R4876 n1_16271_248 n1_16364_248 5.314286e-01
R4877 n1_16364_248 n1_18150_248 1.020571e+01
R4878 n1_18150_248 n1_18333_248 1.045714e+00
R4879 n1_18333_248 n1_18521_248 1.074286e+00
R4880 n1_18521_248 n1_18614_248 5.314286e-01
R4881 n1_18614_248 n1_20583_248 1.125143e+01
R4882 n1_11400_431 n1_11583_431 1.045714e+00
R4883 n1_11583_431 n1_11630_431 2.685714e-01
R4884 n1_11630_431 n1_11771_431 8.057143e-01
R4885 n1_11771_431 n1_11864_431 5.314286e-01
R4886 n1_11864_431 n1_13650_431 1.020571e+01
R4887 n1_13650_431 n1_13833_431 1.045714e+00
R4888 n1_13833_431 n1_13880_431 2.685714e-01
R4889 n1_13880_431 n1_14021_431 8.057143e-01
R4890 n1_14021_431 n1_14114_431 5.314286e-01
R4891 n1_14114_431 n1_15900_431 1.020571e+01
R4892 n1_15900_431 n1_16083_431 1.045714e+00
R4893 n1_16083_431 n1_16130_431 2.685714e-01
R4894 n1_16130_431 n1_16271_431 8.057143e-01
R4895 n1_16271_431 n1_16364_431 5.314286e-01
R4896 n1_16364_431 n1_18150_431 1.020571e+01
R4897 n1_18150_431 n1_18333_431 1.045714e+00
R4898 n1_18333_431 n1_18380_431 2.685714e-01
R4899 n1_18380_431 n1_18521_431 8.057143e-01
R4900 n1_18521_431 n1_18614_431 5.314286e-01
R4901 n1_18614_431 n1_20583_431 1.125143e+01
R4902 n1_20583_431 n1_20630_431 2.685714e-01
R4903 n1_11400_464 n1_11583_464 1.045714e+00
R4904 n1_11583_464 n1_11630_464 2.685714e-01
R4905 n1_11630_464 n1_11864_464 1.337143e+00
R4906 n1_11864_464 n1_13650_464 1.020571e+01
R4907 n1_13650_464 n1_13833_464 1.045714e+00
R4908 n1_13833_464 n1_13880_464 2.685714e-01
R4909 n1_13880_464 n1_14114_464 1.337143e+00
R4910 n1_14114_464 n1_15900_464 1.020571e+01
R4911 n1_15900_464 n1_16083_464 1.045714e+00
R4912 n1_16083_464 n1_16130_464 2.685714e-01
R4913 n1_16130_464 n1_16364_464 1.337143e+00
R4914 n1_16364_464 n1_18150_464 1.020571e+01
R4915 n1_18150_464 n1_18333_464 1.045714e+00
R4916 n1_18333_464 n1_18380_464 2.685714e-01
R4917 n1_18380_464 n1_18614_464 1.337143e+00
R4918 n1_18614_464 n1_20583_464 1.125143e+01
R4919 n1_20583_464 n1_20630_464 2.685714e-01
R4920 n1_11400_647 n1_11583_647 1.045714e+00
R4921 n1_11583_647 n1_11771_647 1.074286e+00
R4922 n1_11771_647 n1_11864_647 5.314286e-01
R4923 n1_11864_647 n1_13650_647 1.020571e+01
R4924 n1_13650_647 n1_13833_647 1.045714e+00
R4925 n1_13833_647 n1_14021_647 1.074286e+00
R4926 n1_14021_647 n1_14114_647 5.314286e-01
R4927 n1_14114_647 n1_15900_647 1.020571e+01
R4928 n1_15900_647 n1_16083_647 1.045714e+00
R4929 n1_16083_647 n1_16271_647 1.074286e+00
R4930 n1_16271_647 n1_16364_647 5.314286e-01
R4931 n1_16364_647 n1_18150_647 1.020571e+01
R4932 n1_18150_647 n1_18333_647 1.045714e+00
R4933 n1_18333_647 n1_18521_647 1.074286e+00
R4934 n1_18521_647 n1_18614_647 5.314286e-01
R4935 n1_18614_647 n1_20583_647 1.125143e+01
R4936 n1_20583_647 n1_20771_647 1.074286e+00
R4937 n1_11400_680 n1_11583_680 1.045714e+00
R4938 n1_11583_680 n1_11771_680 1.074286e+00
R4939 n1_11771_680 n1_11864_680 5.314286e-01
R4940 n1_11864_680 n1_13650_680 1.020571e+01
R4941 n1_13650_680 n1_13833_680 1.045714e+00
R4942 n1_13833_680 n1_14021_680 1.074286e+00
R4943 n1_14021_680 n1_14114_680 5.314286e-01
R4944 n1_14114_680 n1_15900_680 1.020571e+01
R4945 n1_15900_680 n1_16083_680 1.045714e+00
R4946 n1_16083_680 n1_16271_680 1.074286e+00
R4947 n1_16271_680 n1_16364_680 5.314286e-01
R4948 n1_16364_680 n1_18150_680 1.020571e+01
R4949 n1_18150_680 n1_18333_680 1.045714e+00
R4950 n1_18333_680 n1_18521_680 1.074286e+00
R4951 n1_18521_680 n1_18614_680 5.314286e-01
R4952 n1_18614_680 n1_20583_680 1.125143e+01
R4953 n1_20583_680 n1_20771_680 1.074286e+00
R4954 n1_11400_863 n1_11583_863 1.045714e+00
R4955 n1_11583_863 n1_11771_863 1.074286e+00
R4956 n1_11771_863 n1_11864_863 5.314286e-01
R4957 n1_11864_863 n1_13650_863 1.020571e+01
R4958 n1_13650_863 n1_13833_863 1.045714e+00
R4959 n1_13833_863 n1_14021_863 1.074286e+00
R4960 n1_14021_863 n1_14114_863 5.314286e-01
R4961 n1_14114_863 n1_15900_863 1.020571e+01
R4962 n1_15900_863 n1_16083_863 1.045714e+00
R4963 n1_16083_863 n1_16271_863 1.074286e+00
R4964 n1_16271_863 n1_16364_863 5.314286e-01
R4965 n1_16364_863 n1_18150_863 1.020571e+01
R4966 n1_18150_863 n1_18333_863 1.045714e+00
R4967 n1_18333_863 n1_18521_863 1.074286e+00
R4968 n1_18521_863 n1_18614_863 5.314286e-01
R4969 n1_18614_863 n1_20583_863 1.125143e+01
R4970 n1_20583_863 n1_20771_863 1.074286e+00
R4971 n1_11400_896 n1_11583_896 1.045714e+00
R4972 n1_11583_896 n1_11771_896 1.074286e+00
R4973 n1_11771_896 n1_11864_896 5.314286e-01
R4974 n1_11864_896 n1_13650_896 1.020571e+01
R4975 n1_13650_896 n1_13833_896 1.045714e+00
R4976 n1_13833_896 n1_14021_896 1.074286e+00
R4977 n1_14021_896 n1_14114_896 5.314286e-01
R4978 n1_14114_896 n1_15900_896 1.020571e+01
R4979 n1_15900_896 n1_16083_896 1.045714e+00
R4980 n1_16083_896 n1_16271_896 1.074286e+00
R4981 n1_16271_896 n1_16364_896 5.314286e-01
R4982 n1_16364_896 n1_18150_896 1.020571e+01
R4983 n1_18150_896 n1_18333_896 1.045714e+00
R4984 n1_18333_896 n1_18521_896 1.074286e+00
R4985 n1_18521_896 n1_18614_896 5.314286e-01
R4986 n1_18614_896 n1_20583_896 1.125143e+01
R4987 n1_20583_896 n1_20771_896 1.074286e+00
R4988 n1_11400_1079 n1_11583_1079 1.045714e+00
R4989 n1_11583_1079 n1_11771_1079 1.074286e+00
R4990 n1_11771_1079 n1_11864_1079 5.314286e-01
R4991 n1_11864_1079 n1_13650_1079 1.020571e+01
R4992 n1_13650_1079 n1_13833_1079 1.045714e+00
R4993 n1_13833_1079 n1_14021_1079 1.074286e+00
R4994 n1_14021_1079 n1_14114_1079 5.314286e-01
R4995 n1_14114_1079 n1_15900_1079 1.020571e+01
R4996 n1_15900_1079 n1_16083_1079 1.045714e+00
R4997 n1_16083_1079 n1_16271_1079 1.074286e+00
R4998 n1_16271_1079 n1_16364_1079 5.314286e-01
R4999 n1_16364_1079 n1_18150_1079 1.020571e+01
R5000 n1_18150_1079 n1_18333_1079 1.045714e+00
R5001 n1_18333_1079 n1_18521_1079 1.074286e+00
R5002 n1_18521_1079 n1_18614_1079 5.314286e-01
R5003 n1_18614_1079 n1_20583_1079 1.125143e+01
R5004 n1_20583_1079 n1_20771_1079 1.074286e+00
R5005 n1_11400_18548 n1_11583_18548 4.575000e-01
R5006 n1_11583_18548 n1_11630_18548 1.175000e-01
R5007 n1_11630_18548 n1_11771_18548 3.525000e-01
R5008 n1_11583_2760 n1_11630_2760 3.357143e-02
R5009 n1_11630_2760 n1_11771_2760 1.007143e-01
R5010 n1_11583_5566 n1_11771_5566 1.342857e-01
R5011 n1_11583_6646 n1_11771_6646 1.342857e-01
R5012 n1_11583_14012 n1_11630_14012 1.175000e-01
R5013 n1_11630_14012 n1_11771_14012 3.525000e-01
R5014 n1_11583_14220 n1_11771_14220 2.425806e-01
R5015 n1_11583_14660 n1_11771_14660 4.700000e-01
R5016 n1_11583_15740 n1_11771_15740 4.700000e-01
R5017 n1_11583_15956 n1_11771_15956 4.700000e-01
R5018 n1_11583_16172 n1_11630_16172 1.175000e-01
R5019 n1_11630_16172 n1_11771_16172 3.525000e-01
R5020 n1_11583_17468 n1_11771_17468 4.700000e-01
R5021 n1_11400_19412 n1_11583_19412 4.575000e-01
R5022 n1_11583_19412 n1_11771_19412 4.700000e-01
R5023 n1_11400_1894 n1_11583_1894 1.307143e-01
R5024 n1_11583_1894 n1_11771_1894 1.342857e-01
R5025 n1_11771_1894 n1_11864_1894 6.642857e-02
R5026 n1_11583_2974 n1_11771_2974 1.342857e-01
R5027 n1_11583_3622 n1_11771_3622 1.342857e-01
R5028 n1_11583_4270 n1_11771_4270 1.342857e-01
R5029 n1_11583_4702 n1_11771_4702 1.342857e-01
R5030 n1_11583_5350 n1_11771_5350 1.342857e-01
R5031 n1_11583_7294 n1_11630_7294 3.357143e-02
R5032 n1_11630_7294 n1_11771_7294 1.007143e-01
R5033 n1_11583_7510 n1_11771_7510 1.342857e-01
R5034 n1_11583_17244 n1_11771_17244 2.425806e-01
R5035 n1_11400_18764 n1_11583_18764 4.575000e-01
R5036 n1_11583_18764 n1_11771_18764 4.700000e-01
R5037 n1_11771_18764 n1_11864_18764 2.325000e-01
R5038 n1_11583_7078 n1_11771_7078 1.342857e-01
R5039 n1_11400_383 n1_11583_383 1.307143e-01
R5040 n1_11583_383 n1_11771_383 1.342857e-01
R5041 n1_11771_383 n1_11864_383 6.642857e-02
R5042 n1_11864_383 n1_13650_383 1.275714e+00
R5043 n1_13650_383 n1_13833_383 1.307143e-01
R5044 n1_13833_383 n1_14021_383 1.342857e-01
R5045 n1_14021_383 n1_14114_383 6.642857e-02
R5046 n1_14114_383 n1_15900_383 1.275714e+00
R5047 n1_15900_383 n1_16083_383 1.307143e-01
R5048 n1_16083_383 n1_16271_383 1.342857e-01
R5049 n1_16271_383 n1_16364_383 6.642857e-02
R5050 n1_16364_383 n1_18150_383 1.275714e+00
R5051 n1_18150_383 n1_18333_383 1.307143e-01
R5052 n1_18333_383 n1_18521_383 1.342857e-01
R5053 n1_18521_383 n1_18614_383 6.642857e-02
R5054 n1_18614_383 n1_20583_383 1.406429e+00
R5055 n1_11400_2543 n1_11583_2543 1.307143e-01
R5056 n1_11583_2543 n1_11771_2543 1.342857e-01
R5057 n1_11771_2543 n1_11864_2543 6.642857e-02
R5058 n1_11864_2543 n1_13650_2543 1.275714e+00
R5059 n1_13650_2543 n1_13833_2543 1.307143e-01
R5060 n1_13833_2543 n1_14021_2543 1.342857e-01
R5061 n1_14021_2543 n1_14114_2543 6.642857e-02
R5062 n1_14114_2543 n1_15900_2543 1.275714e+00
R5063 n1_15900_2543 n1_16083_2543 1.307143e-01
R5064 n1_16083_2543 n1_16271_2543 1.342857e-01
R5065 n1_16271_2543 n1_16364_2543 6.642857e-02
R5066 n1_16364_2543 n1_18150_2543 1.275714e+00
R5067 n1_18150_2543 n1_18333_2543 1.307143e-01
R5068 n1_18333_2543 n1_18521_2543 1.342857e-01
R5069 n1_18521_2543 n1_18614_2543 6.642857e-02
R5070 n1_18614_2543 n1_20583_2543 1.406429e+00
R5071 n1_20583_2543 n1_20771_2543 1.342857e-01
R5072 n1_11400_18527 n1_11583_18527 1.307143e-01
R5073 n1_11583_18527 n1_11630_18527 3.357143e-02
R5074 n1_11630_18527 n1_11771_18527 1.007143e-01
R5075 n1_11771_18527 n1_11864_18527 6.642857e-02
R5076 n1_11864_18527 n1_13650_18527 1.275714e+00
R5077 n1_13650_18527 n1_13833_18527 1.307143e-01
R5078 n1_13833_18527 n1_13880_18527 3.357143e-02
R5079 n1_13880_18527 n1_14021_18527 1.007143e-01
R5080 n1_14021_18527 n1_14114_18527 6.642857e-02
R5081 n1_14114_18527 n1_15900_18527 1.275714e+00
R5082 n1_15900_18527 n1_16083_18527 1.307143e-01
R5083 n1_16083_18527 n1_16130_18527 3.357143e-02
R5084 n1_16130_18527 n1_16271_18527 1.007143e-01
R5085 n1_16271_18527 n1_16364_18527 6.642857e-02
R5086 n1_16364_18527 n1_18150_18527 1.275714e+00
R5087 n1_18150_18527 n1_18333_18527 1.307143e-01
R5088 n1_18333_18527 n1_18380_18527 3.357143e-02
R5089 n1_18380_18527 n1_18521_18527 1.007143e-01
R5090 n1_18521_18527 n1_18614_18527 6.642857e-02
R5091 n1_18614_18527 n1_20583_18527 1.406429e+00
R5092 n1_20583_18527 n1_20630_18527 3.357143e-02
R5093 n1_20630_18527 n1_20771_18527 1.007143e-01
R5094 n1_11400_20687 n1_11583_20687 1.307143e-01
R5095 n1_11583_20687 n1_11630_20687 3.357143e-02
R5096 n1_11630_20687 n1_11771_20687 1.007143e-01
R5097 n1_11771_20687 n1_11864_20687 6.642857e-02
R5098 n1_11864_20687 n1_13650_20687 1.275714e+00
R5099 n1_13650_20687 n1_13833_20687 1.307143e-01
R5100 n1_13833_20687 n1_13880_20687 3.357143e-02
R5101 n1_13880_20687 n1_14021_20687 1.007143e-01
R5102 n1_14021_20687 n1_14114_20687 6.642857e-02
R5103 n1_14114_20687 n1_15900_20687 1.275714e+00
R5104 n1_15900_20687 n1_16083_20687 1.307143e-01
R5105 n1_16083_20687 n1_16130_20687 3.357143e-02
R5106 n1_16130_20687 n1_16271_20687 1.007143e-01
R5107 n1_16271_20687 n1_16364_20687 6.642857e-02
R5108 n1_16364_20687 n1_18150_20687 1.275714e+00
R5109 n1_18150_20687 n1_18333_20687 1.307143e-01
R5110 n1_18333_20687 n1_18380_20687 3.357143e-02
R5111 n1_18380_20687 n1_18521_20687 1.007143e-01
R5112 n1_18521_20687 n1_18614_20687 6.642857e-02
R5113 n1_18614_20687 n1_20583_20687 1.406429e+00
R5114 n1_20583_20687 n1_20630_20687 3.357143e-02
R5115 n1_20630_20687 n1_20771_20687 1.007143e-01
R5116 n1_11583_6862 n1_11771_6862 1.342857e-01
R5117 n1_11583_13774 n1_11771_13774 1.342857e-01
R5118 n1_11583_2542 n1_11771_2542 1.342857e-01
R5119 n1_11771_2542 n1_11864_2542 6.642857e-02
R5120 n1_11583_15948 n1_11771_15948 2.425806e-01
R5121 n1_11583_16604 n1_11771_16604 4.700000e-01
R5122 n1_11583_17684 n1_11771_17684 4.700000e-01
R5123 n1_11583_18332 n1_11771_18332 4.700000e-01
R5124 n1_11583_19404 n1_11771_19404 2.425806e-01
R5125 n1_11771_19404 n1_11864_19404 1.200000e-01
R5126 n1_11583_5782 n1_11771_5782 1.342857e-01
R5127 n1_11583_6430 n1_11771_6430 1.342857e-01
R5128 n1_13833_2877 n1_14021_2877 1.342857e-01
R5129 n1_14021_2877 n1_16083_2877 1.472857e+00
R5130 n1_16083_2877 n1_16271_2877 1.342857e-01
R5131 n1_13650_2445 n1_13833_2445 1.307143e-01
R5132 n1_13833_2445 n1_14021_2445 1.342857e-01
R5133 n1_14021_2445 n1_14114_2445 6.642857e-02
R5134 n1_14114_2445 n1_15900_2445 1.275714e+00
R5135 n1_15900_2445 n1_16083_2445 1.307143e-01
R5136 n1_16083_2445 n1_16271_2445 1.342857e-01
R5137 n1_16271_2445 n1_16364_2445 6.642857e-02
R5138 n1_13833_7845 n1_14021_7845 1.342857e-01
R5139 n1_14021_7845 n1_16083_7845 1.472857e+00
R5140 n1_16083_7845 n1_16271_7845 1.342857e-01
R5141 n1_16271_7845 n1_18333_7845 1.472857e+00
R5142 n1_18333_7845 n1_18521_7845 1.342857e-01
R5143 n1_13833_8925 n1_14021_8925 1.342857e-01
R5144 n1_14021_8925 n1_16083_8925 1.472857e+00
R5145 n1_16083_8925 n1_16271_8925 1.342857e-01
R5146 n1_16271_8925 n1_18333_8925 1.472857e+00
R5147 n1_18333_8925 n1_18521_8925 1.342857e-01
R5148 n1_13833_10005 n1_14021_10005 1.342857e-01
R5149 n1_14021_10005 n1_16083_10005 1.472857e+00
R5150 n1_16083_10005 n1_16271_10005 1.342857e-01
R5151 n1_16271_10005 n1_18333_10005 1.472857e+00
R5152 n1_18333_10005 n1_18521_10005 1.342857e-01
R5153 n1_13833_6430 n1_14021_6430 1.342857e-01
R5154 n1_13833_5782 n1_14021_5782 1.342857e-01
R5155 n1_13833_8806 n1_14021_8806 1.342857e-01
R5156 n1_13833_9886 n1_14021_9886 1.342857e-01
R5157 n1_13833_10988 n1_14021_10988 4.700000e-01
R5158 n1_13833_12068 n1_14021_12068 4.700000e-01
R5159 n1_13833_9022 n1_14021_9022 1.342857e-01
R5160 n1_13833_10102 n1_14021_10102 1.342857e-01
R5161 n1_13833_11204 n1_14021_11204 4.700000e-01
R5162 n1_13833_12284 n1_14021_12284 4.700000e-01
R5163 n1_13833_17684 n1_14021_17684 4.700000e-01
R5164 n1_13833_5134 n1_14021_5134 1.342857e-01
R5165 n1_13833_14220 n1_14021_14220 2.425806e-01
R5166 n1_13833_14868 n1_14021_14868 2.425806e-01
R5167 n1_13833_16604 n1_14021_16604 4.700000e-01
R5168 n1_13833_18324 n1_14021_18324 2.425806e-01
R5169 n1_13650_19412 n1_13833_19412 4.575000e-01
R5170 n1_13833_19412 n1_14021_19412 4.700000e-01
R5171 n1_13650_2542 n1_13833_2542 1.307143e-01
R5172 n1_13833_2542 n1_14021_2542 1.342857e-01
R5173 n1_14021_2542 n1_14114_2542 6.642857e-02
R5174 n1_13833_2974 n1_14021_2974 1.342857e-01
R5175 n1_13833_3622 n1_14021_3622 1.342857e-01
R5176 n1_13833_15524 n1_14021_15524 4.700000e-01
R5177 n1_13833_15956 n1_14021_15956 4.700000e-01
R5178 n1_13650_18764 n1_13833_18764 4.575000e-01
R5179 n1_13833_18764 n1_14021_18764 4.700000e-01
R5180 n1_14021_18764 n1_14114_18764 2.325000e-01
R5181 n1_13833_4270 n1_14021_4270 1.342857e-01
R5182 n1_13833_4702 n1_14021_4702 1.342857e-01
R5183 n1_13833_7942 n1_14021_7942 1.342857e-01
R5184 n1_13650_1894 n1_13833_1894 1.307143e-01
R5185 n1_13833_1894 n1_14021_1894 1.342857e-01
R5186 n1_14021_1894 n1_14114_1894 6.642857e-02
R5187 n1_13833_18332 n1_14021_18332 4.700000e-01
R5188 n1_13833_4054 n1_14021_4054 1.342857e-01
R5189 n1_13833_18094 n1_14021_18094 1.342857e-01
R5190 n1_13833_14652 n1_14021_14652 2.425806e-01
R5191 n1_13833_19404 n1_14021_19404 2.425806e-01
R5192 n1_14021_19404 n1_14114_19404 1.200000e-01
R5193 n1_13833_6646 n1_14021_6646 1.342857e-01
R5194 n1_13833_5350 n1_14021_5350 1.342857e-01
R5195 n1_16083_5253 n1_16271_5253 1.342857e-01
R5196 n1_16271_5253 n1_18333_5253 1.472857e+00
R5197 n1_18333_5253 n1_18521_5253 1.342857e-01
R5198 n1_16083_6333 n1_16271_6333 1.342857e-01
R5199 n1_16271_6333 n1_18333_6333 1.472857e+00
R5200 n1_18333_6333 n1_18521_6333 1.342857e-01
R5201 n1_18521_6333 n1_20583_6333 1.472857e+00
R5202 n1_16083_6430 n1_16271_6430 1.342857e-01
R5203 n1_16083_11204 n1_16271_11204 4.700000e-01
R5204 n1_16083_7942 n1_16271_7942 1.342857e-01
R5205 n1_16083_9022 n1_16271_9022 1.342857e-01
R5206 n1_16083_10102 n1_16271_10102 1.342857e-01
R5207 n1_16083_12284 n1_16271_12284 4.700000e-01
R5208 n1_16083_14652 n1_16271_14652 2.425806e-01
R5209 n1_16083_4702 n1_16271_4702 1.342857e-01
R5210 n1_15900_18764 n1_16083_18764 4.575000e-01
R5211 n1_16083_18764 n1_16271_18764 4.700000e-01
R5212 n1_15900_19412 n1_16083_19412 4.575000e-01
R5213 n1_16083_19412 n1_16271_19412 4.700000e-01
R5214 n1_15900_1894 n1_16083_1894 1.307143e-01
R5215 n1_16083_1894 n1_16271_1894 1.342857e-01
R5216 n1_16271_1894 n1_16364_1894 6.642857e-02
R5217 n1_16083_3406 n1_16271_3406 1.342857e-01
R5218 n1_16083_4486 n1_16271_4486 1.342857e-01
R5219 n1_16083_5566 n1_16271_5566 1.342857e-01
R5220 n1_16083_16604 n1_16271_16604 4.700000e-01
R5221 n1_16083_17684 n1_16271_17684 4.700000e-01
R5222 n1_16083_18332 n1_16271_18332 4.700000e-01
R5223 n1_16083_15740 n1_16271_15740 4.700000e-01
R5224 n1_15900_2542 n1_16083_2542 1.307143e-01
R5225 n1_16083_2542 n1_16271_2542 1.342857e-01
R5226 n1_16271_2542 n1_16364_2542 6.642857e-02
R5227 n1_16083_2974 n1_16271_2974 1.342857e-01
R5228 n1_16083_12276 n1_16271_12276 2.425806e-01
R5229 n1_16083_15300 n1_16271_15300 2.425806e-01
R5230 n1_16083_5350 n1_16271_5350 1.342857e-01
R5231 n1_16083_16798 n1_16271_16798 1.342857e-01
R5232 n1_16083_4919 n1_16130_4919 3.357143e-02
R5233 n1_16130_4919 n1_16271_4919 1.007143e-01
R5234 n1_16083_5134 n1_16271_5134 1.342857e-01
R5235 n1_16083_17676 n1_16271_17676 2.425806e-01
R5236 n1_16083_19196 n1_16271_19196 4.700000e-01
R5237 n1_16271_19196 n1_16364_19196 2.325000e-01
R5238 n1_16083_13788 n1_16271_13788 2.425806e-01
R5239 n1_16083_11196 n1_16271_11196 2.425806e-01
R5240 n1_16083_16820 n1_16271_16820 4.700000e-01
R5241 n1_18333_4920 n1_18380_4920 3.357143e-02
R5242 n1_18380_4920 n1_18521_4920 1.007143e-01
R5243 n1_18333_5134 n1_18521_5134 1.342857e-01
R5244 n1_18333_6430 n1_18521_6430 1.342857e-01
R5245 n1_18333_14652 n1_18521_14652 2.425806e-01
R5246 n1_18333_5566 n1_18521_5566 1.342857e-01
R5247 n1_18333_7942 n1_18521_7942 1.342857e-01
R5248 n1_18333_9022 n1_18521_9022 1.342857e-01
R5249 n1_18333_10102 n1_18521_10102 1.342857e-01
R5250 n1_18333_11196 n1_18521_11196 2.425806e-01
R5251 n1_18333_12284 n1_18521_12284 4.700000e-01
R5252 n1_18333_15740 n1_18521_15740 4.700000e-01
R5253 n1_18333_16820 n1_18521_16820 4.700000e-01
R5254 n1_18150_1894 n1_18333_1894 1.307143e-01
R5255 n1_18333_1894 n1_18521_1894 1.342857e-01
R5256 n1_18150_2542 n1_18333_2542 1.307143e-01
R5257 n1_18333_2542 n1_18521_2542 1.342857e-01
R5258 n1_18333_3406 n1_18521_3406 1.342857e-01
R5259 n1_18333_4702 n1_18521_4702 1.342857e-01
R5260 n1_18333_13796 n1_18521_13796 4.700000e-01
R5261 n1_18333_4486 n1_18521_4486 1.342857e-01
R5262 n1_18333_17230 n1_18521_17230 1.342857e-01
R5263 n1_18333_5350 n1_18521_5350 1.342857e-01
R5264 n1_18333_16812 n1_18521_16812 2.425806e-01
R5265 n1_18333_2110 n1_18521_2110 1.342857e-01
R5266 n1_18521_2110 n1_18614_2110 6.642857e-02
R5267 n1_18333_13788 n1_18521_13788 2.425806e-01
R5268 n1_18333_14660 n1_18521_14660 4.700000e-01
R5269 n1_18333_17900 n1_18521_17900 4.700000e-01
R5270 n1_18333_15308 n1_18521_15308 4.700000e-01
R5271 n1_20583_15308 n1_20771_15308 4.700000e-01
R5272 n1_20583_5782 n1_20771_5782 1.342857e-01
R5273 n1_20583_16798 n1_20771_16798 1.342857e-01
v33 _X_n2_15005_16221 0 0
rr5e n2_8255_17346 _X_n2_8255_17346 2.500000e-01
rr202 n3_18380_13971 _X_n3_18380_13971 2.500000e-01
v1f9 _X_n3_20630_11721 0 1.8
v1af _X_n3_9380_7221 0 1.8
rr192 n3_9380_11721 _X_n3_9380_11721 2.500000e-01
v35 _X_n2_15005_15096 0 0
v1 _X_n2_20630_12846 0 0
rr204 n3_16130_13971 _X_n3_16130_13971 2.500000e-01
rr194 n3_380_471 _X_n3_380_471 2.500000e-01
rr14a n2_4880_8346 _X_n2_4880_8346 2.500000e-01
v37 _X_n2_12755_20721 0 0
v3 _X_n2_19505_12846 0 0
rr6a n2_6005_18471 _X_n2_6005_18471 2.500000e-01
rr206 n3_20630_16221 _X_n3_20630_16221 2.500000e-01
rr196 n3_2630_471 _X_n3_2630_471 2.500000e-01
rr14c n2_6005_8346 _X_n2_6005_8346 2.500000e-01
v39 _X_n2_12755_19596 0 0
v1bb _X_n3_380_7221 0 1.8
v5 _X_n2_18380_12846 0 0
v41 _X_n2_12755_15096 0 0
rr6c n2_6005_17346 _X_n2_6005_17346 2.500000e-01
rr208 n3_18380_16221 _X_n3_18380_16221 2.500000e-01
rr198 n3_2630_2721 _X_n3_2630_2721 2.500000e-01
rr14e n2_7130_8346 _X_n2_7130_8346 2.500000e-01
rr210 n3_18380_18471 _X_n3_18380_18471 2.500000e-01
v1bd _X_n3_2630_7221 0 1.8
v7 _X_n2_17255_12846 0 0
v43 _X_n2_12755_13971 0 0
rr6e n2_6005_16221 _X_n2_6005_16221 2.500000e-01
rr212 n3_16130_20721 _X_n3_16130_20721 2.500000e-01
v1bf _X_n3_4880_7221 0 1.8
v9 _X_n2_16130_12846 0 0
v45 _X_n2_12755_12846 0 0
rr214 n3_16130_18471 _X_n3_16130_18471 2.500000e-01
rr15a n2_380_3846 _X_n2_380_3846 2.500000e-01
v47 _X_n2_10505_20721 0 0
rr7a n2_380_17346 _X_n2_380_17346 2.500000e-01
rr216 n3_16130_16221 _X_n3_16130_16221 2.500000e-01
rr15c n2_1505_3846 _X_n2_1505_3846 2.500000e-01
rra n2_15005_12846 _X_n2_15005_12846 2.500000e-01
v49 _X_n2_10505_19596 0 0
v1cb _X_n3_11630_4971 0 1.8
v51 _X_n2_10505_15096 0 0
rr7c n2_1505_17346 _X_n2_1505_17346 2.500000e-01
rr218 n3_13880_20721 _X_n3_13880_20721 2.500000e-01
rr15e n2_2630_3846 _X_n2_2630_3846 2.500000e-01
rrc n2_13880_12846 _X_n2_13880_12846 2.500000e-01
rr220 n3_11630_20721 _X_n3_11630_20721 2.500000e-01
v1cd _X_n3_11630_7221 0 1.8
v53 _X_n2_10505_13971 0 0
rr7e n2_2630_17346 _X_n2_2630_17346 2.500000e-01
rre n2_20630_15096 _X_n2_20630_15096 2.500000e-01
rr222 n3_11630_18471 _X_n3_11630_18471 2.500000e-01
v1cf _X_n3_13880_471 0 1.8
v101 _X_n2_15005_10596 0 0
v55 _X_n2_10505_12846 0 0
rr224 n3_11630_16221 _X_n3_11630_16221 2.500000e-01
rr16a n3_7130_20721 _X_n3_7130_20721 2.500000e-01
v103 _X_n2_13880_10596 0 0
v57 _X_n2_10505_11721 0 0
rr8a n2_4880_15096 _X_n2_4880_15096 2.500000e-01
rr226 n3_11630_13971 _X_n3_11630_13971 2.500000e-01
rr16c n3_7130_18471 _X_n3_7130_18471 2.500000e-01
v105 _X_n2_12755_10596 0 0
v59 _X_n2_8255_20721 0 0
v1db _X_n3_20630_471 0 1.8
v61 _X_n2_8255_16221 0 0
rr8c n2_6005_15096 _X_n2_6005_15096 2.500000e-01
rr228 n3_11630_11721 _X_n3_11630_11721 2.500000e-01
rr16e n3_7130_16221 _X_n3_7130_16221 2.500000e-01
v107 _X_n2_11630_10596 0 0
v1dd _X_n3_20630_2721 0 1.8
v63 _X_n2_8255_15096 0 0
rr8e n2_380_12846 _X_n2_380_12846 2.500000e-01
v109 _X_n2_1505_471 0 0
v1df _X_n3_18380_2721 0 1.8
v111 _X_n2_3755_3846 0 0
v1b _X_n2_19505_17346 0 0
v65 _X_n2_8255_13971 0 0
rr17a n3_2630_18471 _X_n3_2630_18471 2.500000e-01
v113 _X_n2_6005_471 0 0
v1d _X_n2_18380_17346 0 0
v67 _X_n2_6005_20721 0 0
rr9a n2_7130_12846 _X_n2_7130_12846 2.500000e-01
rr17c n3_380_16221 _X_n3_380_16221 2.500000e-01
v115 _X_n2_6005_1596 0 0
v1f _X_n2_20630_19596 0 0
v69 _X_n2_6005_19596 0 0
v1eb _X_n3_16130_7221 0 1.8
v71 _X_n2_3755_20721 0 0
rr9c n2_8255_12846 _X_n2_8255_12846 2.500000e-01
rr17e n3_2630_16221 _X_n3_2630_16221 2.500000e-01
v117 _X_n2_6005_2721 0 0
v1ed _X_n3_13880_7221 0 1.8
v73 _X_n2_3755_19596 0 0
rr9e n2_380_10596 _X_n2_380_10596 2.500000e-01
v119 _X_n2_6005_3846 0 0
v1ef _X_n3_20630_9471 0 1.8
v121 _X_n2_8255_1596 0 0
v2b _X_n2_15005_20721 0 0
v75 _X_n2_3755_18471 0 0
rr18a n3_380_11721 _X_n3_380_11721 2.500000e-01
v123 _X_n2_8255_2721 0 0
v2d _X_n2_15005_19596 0 0
v77 _X_n2_1505_20721 0 0
rr18c n3_2630_11721 _X_n3_2630_11721 2.500000e-01
v125 _X_n2_8255_3846 0 0
v2f _X_n2_15005_18471 0 0
v79 _X_n2_380_19596 0 0
v1fb _X_n3_18380_11721 0 1.8
* vias from: 2 to 2
v81 _X_n2_3755_17346 0 0
rr18e n3_4880_11721 _X_n3_4880_11721 2.500000e-01
v127 _X_n2_8255_4971 0 0
v1fd _X_n3_16130_11721 0 1.8
v83 _X_n2_380_15096 0 0
v129 _X_n2_8255_6096 0 0
v1ff _X_n3_13880_11721 0 1.8
v131 _X_n2_10505_1596 0 0
v3b _X_n2_12755_18471 0 0
v85 _X_n2_1505_15096 0 0
rr20a n3_20630_18471 _X_n3_20630_18471 2.500000e-01
rr19a n3_4880_471 _X_n3_4880_471 2.500000e-01
v133 _X_n2_10505_2721 0 0
v3d _X_n2_12755_17346 0 0
v87 _X_n2_2630_15096 0 0
rr20c n3_20630_20721 _X_n3_20630_20721 2.500000e-01
rr19c n3_4880_2721 _X_n3_4880_2721 2.500000e-01
v135 _X_n2_10505_3846 0 0
v3f _X_n2_12755_16221 0 0
v89 _X_n2_3755_15096 0 0
vb _X_n2_15005_12846 0 0
v91 _X_n2_1505_12846 0 0
rr20e n3_18380_20721 _X_n3_18380_20721 2.500000e-01
rr19e n3_4880_4971 _X_n3_4880_4971 2.500000e-01
v137 _X_n2_10505_4971 0 0
vd _X_n2_13880_12846 0 0
v93 _X_n2_2630_12846 0 0
v139 _X_n2_10505_6096 0 0
v141 _X_n2_10505_10596 0 0
vf _X_n2_20630_15096 0 0
v4b _X_n2_10505_18471 0 0
v95 _X_n2_3755_12846 0 0
rr21a n3_13880_18471 _X_n3_13880_18471 2.500000e-01
v143 _X_n2_380_8346 0 0
v4d _X_n2_10505_17346 0 0
v97 _X_n2_4880_12846 0 0
rr21c n3_13880_16221 _X_n3_13880_16221 2.500000e-01
v145 _X_n2_1505_8346 0 0
* layer: M6,GND net: 2
R5274 n2_241_633 n2_241_666 2.095238e-02
R5275 n2_241_666 n2_241_849 1.161905e-01
R5276 n2_241_849 n2_241_882 2.095238e-02
R5277 n2_241_882 n2_241_1065 1.161905e-01
R5278 n2_241_1065 n2_241_1098 2.095238e-02
R5279 n2_241_1098 n2_241_1281 1.161905e-01
R5280 n2_241_1281 n2_241_1314 2.095238e-02
R5281 n2_241_1314 n2_241_1497 1.161905e-01
R5282 n2_241_1497 n2_241_1530 2.095238e-02
R5283 n2_241_1530 n2_241_1549 1.206349e-02
R5284 n2_241_1645 n2_241_1713 4.317460e-02
R5285 n2_241_1713 n2_241_1746 2.095238e-02
R5286 n2_241_1746 n2_241_1929 1.161905e-01
R5287 n2_241_1929 n2_241_1962 2.095238e-02
R5288 n2_241_1962 n2_241_2145 1.161905e-01
R5289 n2_241_2145 n2_241_2178 2.095238e-02
R5290 n2_241_2178 n2_241_2361 1.161905e-01
R5291 n2_241_2361 n2_241_2394 2.095238e-02
R5292 n2_241_2394 n2_241_2577 1.161905e-01
R5293 n2_241_2577 n2_241_2610 2.095238e-02
R5294 n2_241_2610 n2_241_2793 1.161905e-01
R5295 n2_241_2793 n2_241_2826 2.095238e-02
R5296 n2_241_2826 n2_241_3009 1.161905e-01
R5297 n2_241_3009 n2_241_3042 2.095238e-02
R5298 n2_241_3042 n2_241_3225 1.161905e-01
R5299 n2_241_3225 n2_241_3258 2.095238e-02
R5300 n2_241_3258 n2_241_3441 1.161905e-01
R5301 n2_241_3441 n2_241_3474 2.095238e-02
R5302 n2_241_3474 n2_241_3657 1.161905e-01
R5303 n2_241_3657 n2_241_3690 2.095238e-02
R5304 n2_241_3690 n2_241_3799 6.920635e-02
R5305 n2_241_3873 n2_241_3895 1.396825e-02
R5306 n2_241_3895 n2_241_3906 6.984127e-03
R5307 n2_241_3906 n2_241_4089 1.161905e-01
R5308 n2_241_4089 n2_241_4122 2.095238e-02
R5309 n2_241_4122 n2_241_4305 1.161905e-01
R5310 n2_241_4305 n2_241_4338 2.095238e-02
R5311 n2_241_4338 n2_241_4375 2.349206e-02
R5312 n2_241_4375 n2_241_4521 9.269841e-02
R5313 n2_241_4521 n2_241_4554 2.095238e-02
R5314 n2_241_4554 n2_241_4737 1.161905e-01
R5315 n2_241_4737 n2_241_4770 2.095238e-02
R5316 n2_241_4770 n2_241_4953 1.161905e-01
R5317 n2_241_4953 n2_241_4986 2.095238e-02
R5318 n2_241_4986 n2_241_5169 1.161905e-01
R5319 n2_241_5169 n2_241_5202 2.095238e-02
R5320 n2_241_5202 n2_241_5385 1.161905e-01
R5321 n2_241_5385 n2_241_5418 2.095238e-02
R5322 n2_241_5418 n2_241_5601 1.161905e-01
R5323 n2_241_5601 n2_241_5634 2.095238e-02
R5324 n2_241_5634 n2_241_5817 1.161905e-01
R5325 n2_241_5817 n2_241_5850 2.095238e-02
R5326 n2_241_5850 n2_241_6033 1.161905e-01
R5327 n2_241_6033 n2_241_6049 1.015873e-02
R5328 n2_241_6049 n2_241_6066 1.079365e-02
R5329 n2_241_6145 n2_241_6249 6.603175e-02
R5330 n2_241_6249 n2_241_6282 2.095238e-02
R5331 n2_241_6282 n2_241_6465 1.161905e-01
R5332 n2_241_6465 n2_241_6498 2.095238e-02
R5333 n2_241_6498 n2_241_6681 1.161905e-01
R5334 n2_241_6681 n2_241_6714 2.095238e-02
R5335 n2_241_6714 n2_241_6897 1.161905e-01
R5336 n2_241_6897 n2_241_6930 2.095238e-02
R5337 n2_241_6930 n2_241_7113 1.161905e-01
R5338 n2_241_7113 n2_241_7146 2.095238e-02
R5339 n2_241_7146 n2_241_7329 1.161905e-01
R5340 n2_241_7329 n2_241_7362 2.095238e-02
R5341 n2_241_7362 n2_241_7545 1.161905e-01
R5342 n2_241_7545 n2_241_7578 2.095238e-02
R5343 n2_241_7578 n2_241_7761 1.161905e-01
R5344 n2_241_7761 n2_241_7794 2.095238e-02
R5345 n2_241_7794 n2_241_7977 1.161905e-01
R5346 n2_241_7977 n2_241_8010 2.095238e-02
R5347 n2_241_8010 n2_241_8193 1.161905e-01
R5348 n2_241_8193 n2_241_8226 2.095238e-02
R5349 n2_241_8226 n2_241_8299 4.634921e-02
R5350 n2_241_8395 n2_241_8409 8.888889e-03
R5351 n2_241_8409 n2_241_8442 2.095238e-02
R5352 n2_241_8442 n2_241_8625 1.161905e-01
R5353 n2_241_8625 n2_241_8658 2.095238e-02
R5354 n2_241_8658 n2_241_8841 1.161905e-01
R5355 n2_241_8841 n2_241_8874 2.095238e-02
R5356 n2_241_8874 n2_241_9057 1.161905e-01
R5357 n2_241_9057 n2_241_9090 2.095238e-02
R5358 n2_241_9090 n2_241_9273 1.161905e-01
R5359 n2_241_9273 n2_241_9306 2.095238e-02
R5360 n2_241_9306 n2_241_9489 1.161905e-01
R5361 n2_241_9489 n2_241_9522 2.095238e-02
R5362 n2_241_9522 n2_241_9705 1.161905e-01
R5363 n2_241_9705 n2_241_9738 2.095238e-02
R5364 n2_241_9738 n2_241_9921 1.161905e-01
R5365 n2_241_9921 n2_241_9954 2.095238e-02
R5366 n2_241_9954 n2_241_10137 1.161905e-01
R5367 n2_241_10137 n2_241_10170 2.095238e-02
R5368 n2_241_10170 n2_241_10353 1.161905e-01
R5369 n2_241_10353 n2_241_10386 2.095238e-02
R5370 n2_241_10386 n2_241_10549 1.034921e-01
R5371 n2_241_10549 n2_241_10569 1.269841e-02
R5372 n2_241_10645 n2_241_10785 8.888889e-02
R5373 n2_241_10785 n2_241_10818 2.095238e-02
R5374 n2_241_10818 n2_241_11001 1.161905e-01
R5375 n2_241_11001 n2_241_11034 2.095238e-02
R5376 n2_241_11034 n2_241_11217 1.161905e-01
R5377 n2_241_11217 n2_241_11250 2.095238e-02
R5378 n2_241_11250 n2_241_11433 1.161905e-01
R5379 n2_241_11433 n2_241_11466 2.095238e-02
R5380 n2_241_11466 n2_241_11649 1.161905e-01
R5381 n2_241_11649 n2_241_11682 2.095238e-02
R5382 n2_241_11682 n2_241_11865 1.161905e-01
R5383 n2_241_11865 n2_241_11898 2.095238e-02
R5384 n2_241_11898 n2_241_12081 1.161905e-01
R5385 n2_241_12081 n2_241_12114 2.095238e-02
R5386 n2_241_12114 n2_241_12297 1.161905e-01
R5387 n2_241_12297 n2_241_12330 2.095238e-02
R5388 n2_241_12330 n2_241_12513 1.161905e-01
R5389 n2_241_12513 n2_241_12546 2.095238e-02
R5390 n2_241_12546 n2_241_12729 1.161905e-01
R5391 n2_241_12729 n2_241_12762 2.095238e-02
R5392 n2_241_12762 n2_241_12799 2.349206e-02
R5393 n2_241_12895 n2_241_12945 3.174603e-02
R5394 n2_241_12945 n2_241_12978 2.095238e-02
R5395 n2_241_12978 n2_241_13161 1.161905e-01
R5396 n2_241_13161 n2_241_13194 2.095238e-02
R5397 n2_241_13194 n2_241_13377 1.161905e-01
R5398 n2_241_13377 n2_241_13410 2.095238e-02
R5399 n2_241_13410 n2_241_13593 1.161905e-01
R5400 n2_241_13593 n2_241_13626 2.095238e-02
R5401 n2_241_13626 n2_241_13663 2.349206e-02
R5402 n2_241_13663 n2_241_13809 9.269841e-02
R5403 n2_241_13809 n2_241_13842 2.095238e-02
R5404 n2_241_13842 n2_241_14025 1.161905e-01
R5405 n2_241_14025 n2_241_14058 2.095238e-02
R5406 n2_241_14058 n2_241_14241 1.161905e-01
R5407 n2_241_14241 n2_241_14274 2.095238e-02
R5408 n2_241_14274 n2_241_14457 1.161905e-01
R5409 n2_241_14457 n2_241_14490 2.095238e-02
R5410 n2_241_14490 n2_241_14673 1.161905e-01
R5411 n2_241_14673 n2_241_14706 2.095238e-02
R5412 n2_241_14706 n2_241_14889 1.161905e-01
R5413 n2_241_14889 n2_241_14922 2.095238e-02
R5414 n2_241_14922 n2_241_15049 8.063492e-02
R5415 n2_241_15138 n2_241_15145 4.444444e-03
R5416 n2_241_15145 n2_241_15321 1.117460e-01
R5417 n2_241_15321 n2_241_15354 2.095238e-02
R5418 n2_241_15354 n2_241_15537 1.161905e-01
R5419 n2_241_15537 n2_241_15570 2.095238e-02
R5420 n2_241_15570 n2_241_15753 1.161905e-01
R5421 n2_241_15753 n2_241_15786 2.095238e-02
R5422 n2_241_15786 n2_241_15969 1.161905e-01
R5423 n2_241_15969 n2_241_16002 2.095238e-02
R5424 n2_241_16002 n2_241_16185 1.161905e-01
R5425 n2_241_16185 n2_241_16218 2.095238e-02
R5426 n2_241_16218 n2_241_16401 1.161905e-01
R5427 n2_241_16401 n2_241_16434 2.095238e-02
R5428 n2_241_16434 n2_241_16617 1.161905e-01
R5429 n2_241_16617 n2_241_16650 2.095238e-02
R5430 n2_241_16650 n2_241_16833 1.161905e-01
R5431 n2_241_16833 n2_241_16866 2.095238e-02
R5432 n2_241_16866 n2_241_17049 1.161905e-01
R5433 n2_241_17049 n2_241_17082 2.095238e-02
R5434 n2_241_17082 n2_241_17265 1.161905e-01
R5435 n2_241_17265 n2_241_17298 2.095238e-02
R5436 n2_241_17298 n2_241_17299 6.349206e-04
R5437 n2_241_17395 n2_241_17481 5.460317e-02
R5438 n2_241_17481 n2_241_17514 2.095238e-02
R5439 n2_241_17514 n2_241_17697 1.161905e-01
R5440 n2_241_17697 n2_241_17730 2.095238e-02
R5441 n2_241_17730 n2_241_17913 1.161905e-01
R5442 n2_241_17913 n2_241_17946 2.095238e-02
R5443 n2_241_17946 n2_241_17960 8.888889e-03
R5444 n2_241_17960 n2_241_18129 1.073016e-01
R5445 n2_241_18129 n2_241_18162 2.095238e-02
R5446 n2_241_18162 n2_241_18345 1.161905e-01
R5447 n2_241_18345 n2_241_18378 2.095238e-02
R5448 n2_241_18378 n2_241_18561 1.161905e-01
R5449 n2_241_18561 n2_241_18594 2.095238e-02
R5450 n2_241_18594 n2_241_18777 1.161905e-01
R5451 n2_241_18777 n2_241_18810 2.095238e-02
R5452 n2_241_18810 n2_241_18993 1.161905e-01
R5453 n2_241_18993 n2_241_19026 2.095238e-02
R5454 n2_241_19026 n2_241_19040 8.888889e-03
R5455 n2_241_19040 n2_241_19209 1.073016e-01
R5456 n2_241_19209 n2_241_19242 2.095238e-02
R5457 n2_241_19242 n2_241_19256 8.888889e-03
R5458 n2_241_19256 n2_241_19425 1.073016e-01
R5459 n2_241_19425 n2_241_19458 2.095238e-02
R5460 n2_241_19458 n2_241_19472 8.888889e-03
R5461 n2_241_19472 n2_241_19549 4.888889e-02
R5462 n2_241_19641 n2_241_19645 2.539683e-03
R5463 n2_241_19645 n2_241_19674 1.841270e-02
R5464 n2_241_19674 n2_241_19857 1.161905e-01
R5465 n2_241_19857 n2_241_19890 2.095238e-02
R5466 n2_241_19890 n2_241_20073 1.161905e-01
R5467 n2_241_20073 n2_241_20106 2.095238e-02
R5468 n2_241_20106 n2_241_20289 1.161905e-01
R5469 n2_241_20289 n2_241_20322 2.095238e-02
R5470 n2_241_20322 n2_241_20505 1.161905e-01
R5471 n2_241_20505 n2_241_20538 2.095238e-02
R5472 n2_241_1549 n2_380_1549 8.825397e-02
R5473 n2_380_1549 n2_429_1549 3.111111e-02
R5474 n2_241_1645 n2_380_1645 8.825397e-02
R5475 n2_380_1645 n2_429_1645 3.111111e-02
R5476 n2_241_3799 n2_380_3799 8.825397e-02
R5477 n2_380_3799 n2_429_3799 3.111111e-02
R5478 n2_241_3895 n2_380_3895 8.825397e-02
R5479 n2_380_3895 n2_429_3895 3.111111e-02
R5480 n2_241_6049 n2_380_6049 8.825397e-02
R5481 n2_380_6049 n2_429_6049 3.111111e-02
R5482 n2_241_6145 n2_380_6145 8.825397e-02
R5483 n2_380_6145 n2_429_6145 3.111111e-02
R5484 n2_241_8299 n2_380_8299 8.825397e-02
R5485 n2_380_8299 n2_429_8299 3.111111e-02
R5486 n2_241_8395 n2_380_8395 8.825397e-02
R5487 n2_380_8395 n2_429_8395 3.111111e-02
R5488 n2_241_10549 n2_380_10549 8.825397e-02
R5489 n2_380_10549 n2_429_10549 3.111111e-02
R5490 n2_241_10645 n2_380_10645 8.825397e-02
R5491 n2_380_10645 n2_429_10645 3.111111e-02
R5492 n2_241_12799 n2_380_12799 8.825397e-02
R5493 n2_380_12799 n2_429_12799 3.111111e-02
R5494 n2_241_12895 n2_380_12895 8.825397e-02
R5495 n2_380_12895 n2_429_12895 3.111111e-02
R5496 n2_241_15049 n2_380_15049 8.825397e-02
R5497 n2_380_15049 n2_429_15049 3.111111e-02
R5498 n2_241_15145 n2_380_15145 8.825397e-02
R5499 n2_380_15145 n2_429_15145 3.111111e-02
R5500 n2_241_17299 n2_380_17299 8.825397e-02
R5501 n2_380_17299 n2_429_17299 3.111111e-02
R5502 n2_241_17395 n2_380_17395 8.825397e-02
R5503 n2_380_17395 n2_429_17395 3.111111e-02
R5504 n2_241_19549 n2_380_19549 8.825397e-02
R5505 n2_380_19549 n2_429_19549 3.111111e-02
R5506 n2_241_19645 n2_380_19645 8.825397e-02
R5507 n2_380_19645 n2_429_19645 3.111111e-02
R5508 n2_429_633 n2_429_666 2.095238e-02
R5509 n2_429_666 n2_429_849 1.161905e-01
R5510 n2_429_849 n2_429_882 2.095238e-02
R5511 n2_429_882 n2_429_1065 1.161905e-01
R5512 n2_429_1065 n2_429_1098 2.095238e-02
R5513 n2_429_1098 n2_429_1281 1.161905e-01
R5514 n2_429_1281 n2_429_1314 2.095238e-02
R5515 n2_429_1314 n2_429_1497 1.161905e-01
R5516 n2_429_1497 n2_429_1530 2.095238e-02
R5517 n2_429_1530 n2_429_1549 1.206349e-02
R5518 n2_429_1549 n2_429_1645 6.095238e-02
R5519 n2_429_1645 n2_429_1713 4.317460e-02
R5520 n2_429_1713 n2_429_1746 2.095238e-02
R5521 n2_429_1746 n2_429_1929 1.161905e-01
R5522 n2_429_1929 n2_429_1962 2.095238e-02
R5523 n2_429_1962 n2_429_2145 1.161905e-01
R5524 n2_429_2145 n2_429_2178 2.095238e-02
R5525 n2_429_2178 n2_429_2361 1.161905e-01
R5526 n2_429_2361 n2_429_2394 2.095238e-02
R5527 n2_429_2394 n2_429_2577 1.161905e-01
R5528 n2_429_2577 n2_429_2610 2.095238e-02
R5529 n2_429_2826 n2_429_3009 1.161905e-01
R5530 n2_429_3009 n2_429_3042 2.095238e-02
R5531 n2_429_3042 n2_429_3225 1.161905e-01
R5532 n2_429_3225 n2_429_3258 2.095238e-02
R5533 n2_429_3258 n2_429_3441 1.161905e-01
R5534 n2_429_3441 n2_429_3474 2.095238e-02
R5535 n2_429_3474 n2_429_3657 1.161905e-01
R5536 n2_429_3657 n2_429_3690 2.095238e-02
R5537 n2_429_3690 n2_429_3799 6.920635e-02
R5538 n2_429_3799 n2_429_3873 4.698413e-02
R5539 n2_429_3873 n2_429_3895 1.396825e-02
R5540 n2_429_3895 n2_429_3906 6.984127e-03
R5541 n2_429_3906 n2_429_4089 1.161905e-01
R5542 n2_429_4089 n2_429_4122 2.095238e-02
R5543 n2_429_4122 n2_429_4305 1.161905e-01
R5544 n2_429_4305 n2_429_4338 2.095238e-02
R5545 n2_429_4338 n2_429_4375 2.349206e-02
R5546 n2_429_4375 n2_429_4521 9.269841e-02
R5547 n2_429_4521 n2_429_4554 2.095238e-02
R5548 n2_429_4554 n2_429_4737 1.161905e-01
R5549 n2_429_4737 n2_429_4770 2.095238e-02
R5550 n2_429_5169 n2_429_5202 2.095238e-02
R5551 n2_429_5202 n2_429_5385 1.161905e-01
R5552 n2_429_5385 n2_429_5418 2.095238e-02
R5553 n2_429_5418 n2_429_5601 1.161905e-01
R5554 n2_429_5601 n2_429_5634 2.095238e-02
R5555 n2_429_5634 n2_429_5817 1.161905e-01
R5556 n2_429_5817 n2_429_5850 2.095238e-02
R5557 n2_429_5850 n2_429_6033 1.161905e-01
R5558 n2_429_6033 n2_429_6049 1.015873e-02
R5559 n2_429_6049 n2_429_6066 1.079365e-02
R5560 n2_429_6066 n2_429_6145 5.015873e-02
R5561 n2_429_6145 n2_429_6249 6.603175e-02
R5562 n2_429_6249 n2_429_6282 2.095238e-02
R5563 n2_429_6282 n2_429_6465 1.161905e-01
R5564 n2_429_6465 n2_429_6498 2.095238e-02
R5565 n2_429_6498 n2_429_6681 1.161905e-01
R5566 n2_429_6681 n2_429_6714 2.095238e-02
R5567 n2_429_6714 n2_429_6897 1.161905e-01
R5568 n2_429_6897 n2_429_6930 2.095238e-02
R5569 n2_429_6930 n2_429_7113 1.161905e-01
R5570 n2_429_7329 n2_429_7362 2.095238e-02
R5571 n2_429_7362 n2_429_7545 1.161905e-01
R5572 n2_429_7545 n2_429_7578 2.095238e-02
R5573 n2_429_7578 n2_429_7761 1.161905e-01
R5574 n2_429_7761 n2_429_7794 2.095238e-02
R5575 n2_429_7794 n2_429_7977 1.161905e-01
R5576 n2_429_7977 n2_429_8010 2.095238e-02
R5577 n2_429_8010 n2_429_8193 1.161905e-01
R5578 n2_429_8193 n2_429_8226 2.095238e-02
R5579 n2_429_8226 n2_429_8299 4.634921e-02
R5580 n2_429_8299 n2_429_8395 6.095238e-02
R5581 n2_429_8395 n2_429_8409 8.888889e-03
R5582 n2_429_8409 n2_429_8442 2.095238e-02
R5583 n2_429_8442 n2_429_8625 1.161905e-01
R5584 n2_429_8625 n2_429_8658 2.095238e-02
R5585 n2_429_8658 n2_429_8841 1.161905e-01
R5586 n2_429_8841 n2_429_8874 2.095238e-02
R5587 n2_429_8874 n2_429_9057 1.161905e-01
R5588 n2_429_9057 n2_429_9090 2.095238e-02
R5589 n2_429_9090 n2_429_9273 1.161905e-01
R5590 n2_429_9273 n2_429_9306 2.095238e-02
R5591 n2_429_9705 n2_429_9738 2.095238e-02
R5592 n2_429_9738 n2_429_9921 1.161905e-01
R5593 n2_429_9921 n2_429_9954 2.095238e-02
R5594 n2_429_9954 n2_429_10137 1.161905e-01
R5595 n2_429_10137 n2_429_10170 2.095238e-02
R5596 n2_429_10170 n2_429_10353 1.161905e-01
R5597 n2_429_10353 n2_429_10386 2.095238e-02
R5598 n2_429_10386 n2_429_10549 1.034921e-01
R5599 n2_429_10549 n2_429_10569 1.269841e-02
R5600 n2_429_10569 n2_429_10602 2.095238e-02
R5601 n2_429_10602 n2_429_10645 2.730159e-02
R5602 n2_429_10645 n2_429_10785 8.888889e-02
R5603 n2_429_10785 n2_429_10818 2.095238e-02
R5604 n2_429_10818 n2_429_11001 1.161905e-01
R5605 n2_429_11001 n2_429_11034 2.095238e-02
R5606 n2_429_11034 n2_429_11217 1.161905e-01
R5607 n2_429_11217 n2_429_11250 2.095238e-02
R5608 n2_429_11250 n2_429_11433 1.161905e-01
R5609 n2_429_11433 n2_429_11466 2.095238e-02
R5610 n2_429_11865 n2_429_11898 2.095238e-02
R5611 n2_429_11898 n2_429_12081 1.161905e-01
R5612 n2_429_12081 n2_429_12114 2.095238e-02
R5613 n2_429_12114 n2_429_12297 1.161905e-01
R5614 n2_429_12297 n2_429_12330 2.095238e-02
R5615 n2_429_12330 n2_429_12513 1.161905e-01
R5616 n2_429_12513 n2_429_12546 2.095238e-02
R5617 n2_429_12546 n2_429_12729 1.161905e-01
R5618 n2_429_12729 n2_429_12762 2.095238e-02
R5619 n2_429_12762 n2_429_12799 2.349206e-02
R5620 n2_429_12799 n2_429_12895 6.095238e-02
R5621 n2_429_12895 n2_429_12945 3.174603e-02
R5622 n2_429_12945 n2_429_12978 2.095238e-02
R5623 n2_429_12978 n2_429_13161 1.161905e-01
R5624 n2_429_13161 n2_429_13194 2.095238e-02
R5625 n2_429_13194 n2_429_13377 1.161905e-01
R5626 n2_429_13377 n2_429_13410 2.095238e-02
R5627 n2_429_13410 n2_429_13593 1.161905e-01
R5628 n2_429_13593 n2_429_13626 2.095238e-02
R5629 n2_429_13626 n2_429_13663 2.349206e-02
R5630 n2_429_13663 n2_429_13809 9.269841e-02
R5631 n2_429_13809 n2_429_13842 2.095238e-02
R5632 n2_429_14241 n2_429_14274 2.095238e-02
R5633 n2_429_14274 n2_429_14457 1.161905e-01
R5634 n2_429_14457 n2_429_14490 2.095238e-02
R5635 n2_429_14490 n2_429_14673 1.161905e-01
R5636 n2_429_14673 n2_429_14706 2.095238e-02
R5637 n2_429_14706 n2_429_14889 1.161905e-01
R5638 n2_429_14889 n2_429_14922 2.095238e-02
R5639 n2_429_14922 n2_429_15049 8.063492e-02
R5640 n2_429_15049 n2_429_15105 3.555556e-02
R5641 n2_429_15105 n2_429_15138 2.095238e-02
R5642 n2_429_15138 n2_429_15145 4.444444e-03
R5643 n2_429_15145 n2_429_15321 1.117460e-01
R5644 n2_429_15321 n2_429_15354 2.095238e-02
R5645 n2_429_15354 n2_429_15537 1.161905e-01
R5646 n2_429_15537 n2_429_15570 2.095238e-02
R5647 n2_429_15570 n2_429_15753 1.161905e-01
R5648 n2_429_15753 n2_429_15786 2.095238e-02
R5649 n2_429_15786 n2_429_15969 1.161905e-01
R5650 n2_429_15969 n2_429_16002 2.095238e-02
R5651 n2_429_16401 n2_429_16434 2.095238e-02
R5652 n2_429_16434 n2_429_16617 1.161905e-01
R5653 n2_429_16617 n2_429_16650 2.095238e-02
R5654 n2_429_16650 n2_429_16833 1.161905e-01
R5655 n2_429_16833 n2_429_16866 2.095238e-02
R5656 n2_429_16866 n2_429_17049 1.161905e-01
R5657 n2_429_17049 n2_429_17082 2.095238e-02
R5658 n2_429_17082 n2_429_17265 1.161905e-01
R5659 n2_429_17265 n2_429_17298 2.095238e-02
R5660 n2_429_17298 n2_429_17299 6.349206e-04
R5661 n2_429_17299 n2_429_17395 6.095238e-02
R5662 n2_429_17395 n2_429_17481 5.460317e-02
R5663 n2_429_17481 n2_429_17514 2.095238e-02
R5664 n2_429_17514 n2_429_17697 1.161905e-01
R5665 n2_429_17697 n2_429_17730 2.095238e-02
R5666 n2_429_17730 n2_429_17913 1.161905e-01
R5667 n2_429_17913 n2_429_17946 2.095238e-02
R5668 n2_429_17946 n2_429_17960 8.888889e-03
R5669 n2_429_17960 n2_429_18129 1.073016e-01
R5670 n2_429_18129 n2_429_18162 2.095238e-02
R5671 n2_429_18162 n2_429_18345 1.161905e-01
R5672 n2_429_18594 n2_429_18777 1.161905e-01
R5673 n2_429_18777 n2_429_18810 2.095238e-02
R5674 n2_429_18810 n2_429_18993 1.161905e-01
R5675 n2_429_18993 n2_429_19026 2.095238e-02
R5676 n2_429_19026 n2_429_19040 8.888889e-03
R5677 n2_429_19040 n2_429_19209 1.073016e-01
R5678 n2_429_19209 n2_429_19242 2.095238e-02
R5679 n2_429_19242 n2_429_19256 8.888889e-03
R5680 n2_429_19256 n2_429_19425 1.073016e-01
R5681 n2_429_19425 n2_429_19458 2.095238e-02
R5682 n2_429_19458 n2_429_19472 8.888889e-03
R5683 n2_429_19472 n2_429_19549 4.888889e-02
R5684 n2_429_19549 n2_429_19641 5.841270e-02
R5685 n2_429_19641 n2_429_19645 2.539683e-03
R5686 n2_429_19645 n2_429_19674 1.841270e-02
R5687 n2_429_19674 n2_429_19857 1.161905e-01
R5688 n2_429_19857 n2_429_19890 2.095238e-02
R5689 n2_429_19890 n2_429_20073 1.161905e-01
R5690 n2_429_20073 n2_429_20106 2.095238e-02
R5691 n2_429_20106 n2_429_20289 1.161905e-01
R5692 n2_429_20289 n2_429_20322 2.095238e-02
R5693 n2_429_20322 n2_429_20505 1.161905e-01
R5694 n2_429_20505 n2_429_20538 2.095238e-02
R5695 n2_1366_201 n2_1366_234 2.095238e-02
R5696 n2_1366_234 n2_1366_417 1.161905e-01
R5697 n2_1366_417 n2_1366_424 4.444444e-03
R5698 n2_1366_424 n2_1366_450 1.650794e-02
R5699 n2_1366_520 n2_1366_633 7.174603e-02
R5700 n2_1366_633 n2_1366_666 2.095238e-02
R5701 n2_1366_666 n2_1366_849 1.161905e-01
R5702 n2_1366_849 n2_1366_882 2.095238e-02
R5703 n2_1366_882 n2_1366_1065 1.161905e-01
R5704 n2_1366_1065 n2_1366_1098 2.095238e-02
R5705 n2_1366_1098 n2_1366_1281 1.161905e-01
R5706 n2_1366_1281 n2_1366_1314 2.095238e-02
R5707 n2_1366_1314 n2_1366_1497 1.161905e-01
R5708 n2_1366_1497 n2_1366_1530 2.095238e-02
R5709 n2_1366_1530 n2_1366_1713 1.161905e-01
R5710 n2_1366_1713 n2_1366_1746 2.095238e-02
R5711 n2_1366_1746 n2_1366_1760 8.888889e-03
R5712 n2_1366_1760 n2_1366_1929 1.073016e-01
R5713 n2_1366_1929 n2_1366_1962 2.095238e-02
R5714 n2_1366_1962 n2_1366_2145 1.161905e-01
R5715 n2_1366_2145 n2_1366_2178 2.095238e-02
R5716 n2_1366_2178 n2_1366_2361 1.161905e-01
R5717 n2_1366_2361 n2_1366_2394 2.095238e-02
R5718 n2_1366_2394 n2_1366_2577 1.161905e-01
R5719 n2_1366_2577 n2_1366_2610 2.095238e-02
R5720 n2_1366_2610 n2_1366_2793 1.161905e-01
R5721 n2_1366_2793 n2_1366_2826 2.095238e-02
R5722 n2_1366_2826 n2_1366_3009 1.161905e-01
R5723 n2_1366_3009 n2_1366_3042 2.095238e-02
R5724 n2_1366_3042 n2_1366_3225 1.161905e-01
R5725 n2_1366_3225 n2_1366_3258 2.095238e-02
R5726 n2_1366_3258 n2_1366_3272 8.888889e-03
R5727 n2_1366_3272 n2_1366_3441 1.073016e-01
R5728 n2_1366_3441 n2_1366_3474 2.095238e-02
R5729 n2_1366_3474 n2_1366_3657 1.161905e-01
R5730 n2_1366_3657 n2_1366_3690 2.095238e-02
R5731 n2_1366_3690 n2_1366_3704 8.888889e-03
R5732 n2_1366_3704 n2_1366_3799 6.031746e-02
R5733 n2_1366_3873 n2_1366_3895 1.396825e-02
R5734 n2_1366_3895 n2_1366_3906 6.984127e-03
R5735 n2_1366_3906 n2_1366_3920 8.888889e-03
R5736 n2_1366_3920 n2_1366_4089 1.073016e-01
R5737 n2_1366_4089 n2_1366_4122 2.095238e-02
R5738 n2_1366_4122 n2_1366_4159 2.349206e-02
R5739 n2_1366_4159 n2_1366_4305 9.269841e-02
R5740 n2_1366_4305 n2_1366_4338 2.095238e-02
R5741 n2_1366_4338 n2_1366_4352 8.888889e-03
R5742 n2_1366_4352 n2_1366_4375 1.460317e-02
R5743 n2_1366_4375 n2_1366_4521 9.269841e-02
R5744 n2_1366_4521 n2_1366_4554 2.095238e-02
R5745 n2_1366_4554 n2_1366_4737 1.161905e-01
R5746 n2_1366_4737 n2_1366_4770 2.095238e-02
R5747 n2_1366_4770 n2_1366_4953 1.161905e-01
R5748 n2_1366_4953 n2_1366_4986 2.095238e-02
R5749 n2_1366_4986 n2_1366_5169 1.161905e-01
R5750 n2_1366_5169 n2_1366_5202 2.095238e-02
R5751 n2_1366_5202 n2_1366_5385 1.161905e-01
R5752 n2_1366_5385 n2_1366_5418 2.095238e-02
R5753 n2_1366_5418 n2_1366_5432 8.888889e-03
R5754 n2_1366_5432 n2_1366_5601 1.073016e-01
R5755 n2_1366_5601 n2_1366_5634 2.095238e-02
R5756 n2_1366_5634 n2_1366_5817 1.161905e-01
R5757 n2_1366_5817 n2_1366_5850 2.095238e-02
R5758 n2_1366_5850 n2_1366_6033 1.161905e-01
R5759 n2_1366_6033 n2_1366_6049 1.015873e-02
R5760 n2_1366_6049 n2_1366_6066 1.079365e-02
R5761 n2_1366_6145 n2_1366_6249 6.603175e-02
R5762 n2_1366_6249 n2_1366_6282 2.095238e-02
R5763 n2_1366_6282 n2_1366_6465 1.161905e-01
R5764 n2_1366_6465 n2_1366_6498 2.095238e-02
R5765 n2_1366_6498 n2_1366_6535 2.349206e-02
R5766 n2_1366_6535 n2_1366_6681 9.269841e-02
R5767 n2_1366_6681 n2_1366_6714 2.095238e-02
R5768 n2_1366_6714 n2_1366_6897 1.161905e-01
R5769 n2_1366_6897 n2_1366_6930 2.095238e-02
R5770 n2_1366_6930 n2_1366_7113 1.161905e-01
R5771 n2_1366_7113 n2_1366_7146 2.095238e-02
R5772 n2_1366_7146 n2_1366_7329 1.161905e-01
R5773 n2_1366_7329 n2_1366_7362 2.095238e-02
R5774 n2_1366_7362 n2_1366_7545 1.161905e-01
R5775 n2_1366_7545 n2_1366_7578 2.095238e-02
R5776 n2_1366_7578 n2_1366_7761 1.161905e-01
R5777 n2_1366_7761 n2_1366_7794 2.095238e-02
R5778 n2_1366_7794 n2_1366_7808 8.888889e-03
R5779 n2_1366_7808 n2_1366_7977 1.073016e-01
R5780 n2_1366_7977 n2_1366_8010 2.095238e-02
R5781 n2_1366_8010 n2_1366_8193 1.161905e-01
R5782 n2_1366_8193 n2_1366_8226 2.095238e-02
R5783 n2_1366_8226 n2_1366_8299 4.634921e-02
R5784 n2_1366_8395 n2_1366_8409 8.888889e-03
R5785 n2_1366_8409 n2_1366_8442 2.095238e-02
R5786 n2_1366_8442 n2_1366_8625 1.161905e-01
R5787 n2_1366_8625 n2_1366_8658 2.095238e-02
R5788 n2_1366_8658 n2_1366_8841 1.161905e-01
R5789 n2_1366_8841 n2_1366_8874 2.095238e-02
R5790 n2_1366_8874 n2_1366_8888 8.888889e-03
R5791 n2_1366_8888 n2_1366_8911 1.460317e-02
R5792 n2_1366_8911 n2_1366_9057 9.269841e-02
R5793 n2_1366_9057 n2_1366_9090 2.095238e-02
R5794 n2_1366_9090 n2_1366_9273 1.161905e-01
R5795 n2_1366_9273 n2_1366_9306 2.095238e-02
R5796 n2_1366_9306 n2_1366_9489 1.161905e-01
R5797 n2_1366_9489 n2_1366_9522 2.095238e-02
R5798 n2_1366_9522 n2_1366_9705 1.161905e-01
R5799 n2_1366_9705 n2_1366_9738 2.095238e-02
R5800 n2_1366_9738 n2_1366_9921 1.161905e-01
R5801 n2_1366_9921 n2_1366_9954 2.095238e-02
R5802 n2_1366_9954 n2_1366_9968 8.888889e-03
R5803 n2_1366_9968 n2_1366_10137 1.073016e-01
R5804 n2_1366_10137 n2_1366_10170 2.095238e-02
R5805 n2_1366_10170 n2_1366_10353 1.161905e-01
R5806 n2_1366_10353 n2_1366_10386 2.095238e-02
R5807 n2_1366_10386 n2_1366_10549 1.034921e-01
R5808 n2_1366_10549 n2_1366_10569 1.269841e-02
R5809 n2_1366_10645 n2_1366_10785 8.888889e-02
R5810 n2_1366_10785 n2_1366_10818 2.095238e-02
R5811 n2_1366_10818 n2_1366_11001 1.161905e-01
R5812 n2_1366_11001 n2_1366_11034 2.095238e-02
R5813 n2_1366_11034 n2_1366_11048 8.888889e-03
R5814 n2_1366_11048 n2_1366_11071 1.460317e-02
R5815 n2_1366_11071 n2_1366_11217 9.269841e-02
R5816 n2_1366_11217 n2_1366_11250 2.095238e-02
R5817 n2_1366_11250 n2_1366_11433 1.161905e-01
R5818 n2_1366_11433 n2_1366_11466 2.095238e-02
R5819 n2_1366_11466 n2_1366_11649 1.161905e-01
R5820 n2_1366_11649 n2_1366_11682 2.095238e-02
R5821 n2_1366_11682 n2_1366_11865 1.161905e-01
R5822 n2_1366_11865 n2_1366_11898 2.095238e-02
R5823 n2_1366_11898 n2_1366_12081 1.161905e-01
R5824 n2_1366_12081 n2_1366_12114 2.095238e-02
R5825 n2_1366_12114 n2_1366_12128 8.888889e-03
R5826 n2_1366_12128 n2_1366_12297 1.073016e-01
R5827 n2_1366_12297 n2_1366_12330 2.095238e-02
R5828 n2_1366_12330 n2_1366_12513 1.161905e-01
R5829 n2_1366_12513 n2_1366_12546 2.095238e-02
R5830 n2_1366_12546 n2_1366_12729 1.161905e-01
R5831 n2_1366_12729 n2_1366_12762 2.095238e-02
R5832 n2_1366_12762 n2_1366_12799 2.349206e-02
R5833 n2_1366_12895 n2_1366_12945 3.174603e-02
R5834 n2_1366_12945 n2_1366_12978 2.095238e-02
R5835 n2_1366_12978 n2_1366_13161 1.161905e-01
R5836 n2_1366_13161 n2_1366_13194 2.095238e-02
R5837 n2_1366_13194 n2_1366_13377 1.161905e-01
R5838 n2_1366_13377 n2_1366_13410 2.095238e-02
R5839 n2_1366_13410 n2_1366_13447 2.349206e-02
R5840 n2_1366_13447 n2_1366_13593 9.269841e-02
R5841 n2_1366_13593 n2_1366_13626 2.095238e-02
R5842 n2_1366_13626 n2_1366_13663 2.349206e-02
R5843 n2_1366_13663 n2_1366_13809 9.269841e-02
R5844 n2_1366_13809 n2_1366_13842 2.095238e-02
R5845 n2_1366_13842 n2_1366_14025 1.161905e-01
R5846 n2_1366_14025 n2_1366_14058 2.095238e-02
R5847 n2_1366_14058 n2_1366_14241 1.161905e-01
R5848 n2_1366_14241 n2_1366_14274 2.095238e-02
R5849 n2_1366_14274 n2_1366_14457 1.161905e-01
R5850 n2_1366_14457 n2_1366_14490 2.095238e-02
R5851 n2_1366_14490 n2_1366_14504 8.888889e-03
R5852 n2_1366_14504 n2_1366_14673 1.073016e-01
R5853 n2_1366_14673 n2_1366_14706 2.095238e-02
R5854 n2_1366_14706 n2_1366_14889 1.161905e-01
R5855 n2_1366_14889 n2_1366_14922 2.095238e-02
R5856 n2_1366_14922 n2_1366_15049 8.063492e-02
R5857 n2_1366_15138 n2_1366_15145 4.444444e-03
R5858 n2_1366_15145 n2_1366_15321 1.117460e-01
R5859 n2_1366_15321 n2_1366_15354 2.095238e-02
R5860 n2_1366_15354 n2_1366_15368 8.888889e-03
R5861 n2_1366_15368 n2_1366_15537 1.073016e-01
R5862 n2_1366_15537 n2_1366_15570 2.095238e-02
R5863 n2_1366_15570 n2_1366_15753 1.161905e-01
R5864 n2_1366_15753 n2_1366_15786 2.095238e-02
R5865 n2_1366_15786 n2_1366_15969 1.161905e-01
R5866 n2_1366_15969 n2_1366_16002 2.095238e-02
R5867 n2_1366_16002 n2_1366_16185 1.161905e-01
R5868 n2_1366_16185 n2_1366_16218 2.095238e-02
R5869 n2_1366_16218 n2_1366_16401 1.161905e-01
R5870 n2_1366_16401 n2_1366_16434 2.095238e-02
R5871 n2_1366_16434 n2_1366_16471 2.349206e-02
R5872 n2_1366_16471 n2_1366_16617 9.269841e-02
R5873 n2_1366_16617 n2_1366_16650 2.095238e-02
R5874 n2_1366_16650 n2_1366_16687 2.349206e-02
R5875 n2_1366_16687 n2_1366_16833 9.269841e-02
R5876 n2_1366_16833 n2_1366_16866 2.095238e-02
R5877 n2_1366_16866 n2_1366_16880 8.888889e-03
R5878 n2_1366_16880 n2_1366_17049 1.073016e-01
R5879 n2_1366_17049 n2_1366_17082 2.095238e-02
R5880 n2_1366_17082 n2_1366_17265 1.161905e-01
R5881 n2_1366_17265 n2_1366_17298 2.095238e-02
R5882 n2_1366_17298 n2_1366_17299 6.349206e-04
R5883 n2_1366_17395 n2_1366_17481 5.460317e-02
R5884 n2_1366_17481 n2_1366_17514 2.095238e-02
R5885 n2_1366_17514 n2_1366_17528 8.888889e-03
R5886 n2_1366_17528 n2_1366_17697 1.073016e-01
R5887 n2_1366_17697 n2_1366_17730 2.095238e-02
R5888 n2_1366_17730 n2_1366_17913 1.161905e-01
R5889 n2_1366_17913 n2_1366_17946 2.095238e-02
R5890 n2_1366_17946 n2_1366_17960 8.888889e-03
R5891 n2_1366_17960 n2_1366_18129 1.073016e-01
R5892 n2_1366_18129 n2_1366_18162 2.095238e-02
R5893 n2_1366_18162 n2_1366_18345 1.161905e-01
R5894 n2_1366_18345 n2_1366_18378 2.095238e-02
R5895 n2_1366_18378 n2_1366_18561 1.161905e-01
R5896 n2_1366_18561 n2_1366_18594 2.095238e-02
R5897 n2_1366_18594 n2_1366_18777 1.161905e-01
R5898 n2_1366_18777 n2_1366_18810 2.095238e-02
R5899 n2_1366_18810 n2_1366_18993 1.161905e-01
R5900 n2_1366_18993 n2_1366_19026 2.095238e-02
R5901 n2_1366_19026 n2_1366_19040 8.888889e-03
R5902 n2_1366_19040 n2_1366_19209 1.073016e-01
R5903 n2_1366_19209 n2_1366_19242 2.095238e-02
R5904 n2_1366_19242 n2_1366_19256 8.888889e-03
R5905 n2_1366_19256 n2_1366_19425 1.073016e-01
R5906 n2_1366_19425 n2_1366_19458 2.095238e-02
R5907 n2_1366_19458 n2_1366_19472 8.888889e-03
R5908 n2_1366_19472 n2_1366_19641 1.073016e-01
R5909 n2_1366_19641 n2_1366_19674 2.095238e-02
R5910 n2_1366_19674 n2_1366_19857 1.161905e-01
R5911 n2_1366_19857 n2_1366_19890 2.095238e-02
R5912 n2_1366_19890 n2_1366_20073 1.161905e-01
R5913 n2_1366_20073 n2_1366_20106 2.095238e-02
R5914 n2_1366_20106 n2_1366_20289 1.161905e-01
R5915 n2_1366_20289 n2_1366_20322 2.095238e-02
R5916 n2_1366_20322 n2_1366_20505 1.161905e-01
R5917 n2_1366_20505 n2_1366_20538 2.095238e-02
R5918 n2_1366_20538 n2_1366_20674 8.634921e-02
R5919 n2_1366_20754 n2_1366_20770 1.015873e-02
R5920 n2_1366_20770 n2_1366_20937 1.060317e-01
R5921 n2_1366_20937 n2_1366_20970 2.095238e-02
R5922 n2_1366_3799 n2_1505_3799 8.825397e-02
R5923 n2_1505_3799 n2_1554_3799 3.111111e-02
R5924 n2_1366_3895 n2_1505_3895 8.825397e-02
R5925 n2_1505_3895 n2_1554_3895 3.111111e-02
R5926 n2_1366_6049 n2_1505_6049 8.825397e-02
R5927 n2_1505_6049 n2_1554_6049 3.111111e-02
R5928 n2_1366_6145 n2_1505_6145 8.825397e-02
R5929 n2_1505_6145 n2_1554_6145 3.111111e-02
R5930 n2_1366_8299 n2_1505_8299 8.825397e-02
R5931 n2_1505_8299 n2_1554_8299 3.111111e-02
R5932 n2_1366_8395 n2_1505_8395 8.825397e-02
R5933 n2_1505_8395 n2_1554_8395 3.111111e-02
R5934 n2_1366_10549 n2_1505_10549 8.825397e-02
R5935 n2_1505_10549 n2_1554_10549 3.111111e-02
R5936 n2_1366_10645 n2_1505_10645 8.825397e-02
R5937 n2_1505_10645 n2_1554_10645 3.111111e-02
R5938 n2_1366_12799 n2_1505_12799 8.825397e-02
R5939 n2_1505_12799 n2_1554_12799 3.111111e-02
R5940 n2_1366_12895 n2_1505_12895 8.825397e-02
R5941 n2_1505_12895 n2_1554_12895 3.111111e-02
R5942 n2_1366_15049 n2_1505_15049 8.825397e-02
R5943 n2_1505_15049 n2_1554_15049 3.111111e-02
R5944 n2_1366_15145 n2_1505_15145 8.825397e-02
R5945 n2_1505_15145 n2_1554_15145 3.111111e-02
R5946 n2_1366_17299 n2_1505_17299 8.825397e-02
R5947 n2_1505_17299 n2_1554_17299 3.111111e-02
R5948 n2_1366_17395 n2_1505_17395 8.825397e-02
R5949 n2_1505_17395 n2_1554_17395 3.111111e-02
R5950 n2_1366_424 n2_1458_424 5.841270e-02
R5951 n2_1458_424 n2_1505_424 2.984127e-02
R5952 n2_1505_424 n2_1554_424 3.111111e-02
R5953 n2_1554_424 n2_1646_424 5.841270e-02
R5954 n2_1366_520 n2_1458_520 5.841270e-02
R5955 n2_1458_520 n2_1505_520 2.984127e-02
R5956 n2_1505_520 n2_1554_520 3.111111e-02
R5957 n2_1554_520 n2_1646_520 5.841270e-02
R5958 n2_1366_20674 n2_1458_20674 5.841270e-02
R5959 n2_1458_20674 n2_1505_20674 2.984127e-02
R5960 n2_1505_20674 n2_1554_20674 3.111111e-02
R5961 n2_1554_20674 n2_1646_20674 5.841270e-02
R5962 n2_1366_20770 n2_1458_20770 5.841270e-02
R5963 n2_1458_20770 n2_1505_20770 2.984127e-02
R5964 n2_1505_20770 n2_1554_20770 3.111111e-02
R5965 n2_1554_20770 n2_1646_20770 5.841270e-02
R5966 n2_1458_201 n2_1458_234 2.095238e-02
R5967 n2_1458_234 n2_1458_417 1.161905e-01
R5968 n2_1458_417 n2_1458_424 4.444444e-03
R5969 n2_1458_424 n2_1458_450 1.650794e-02
R5970 n2_1458_450 n2_1458_520 4.444444e-02
R5971 n2_1458_520 n2_1458_633 7.174603e-02
R5972 n2_1458_633 n2_1458_666 2.095238e-02
R5973 n2_1458_666 n2_1458_849 1.161905e-01
R5974 n2_1458_849 n2_1458_882 2.095238e-02
R5975 n2_1458_882 n2_1458_1065 1.161905e-01
R5976 n2_1458_1065 n2_1458_1098 2.095238e-02
R5977 n2_1458_1098 n2_1458_1281 1.161905e-01
R5978 n2_1458_1281 n2_1458_1314 2.095238e-02
R5979 n2_1458_1314 n2_1458_1497 1.161905e-01
R5980 n2_1458_19857 n2_1458_19890 2.095238e-02
R5981 n2_1458_19890 n2_1458_20073 1.161905e-01
R5982 n2_1458_20073 n2_1458_20106 2.095238e-02
R5983 n2_1458_20106 n2_1458_20289 1.161905e-01
R5984 n2_1458_20289 n2_1458_20322 2.095238e-02
R5985 n2_1458_20322 n2_1458_20505 1.161905e-01
R5986 n2_1458_20505 n2_1458_20538 2.095238e-02
R5987 n2_1458_20538 n2_1458_20674 8.634921e-02
R5988 n2_1458_20674 n2_1458_20721 2.984127e-02
R5989 n2_1458_20721 n2_1458_20754 2.095238e-02
R5990 n2_1458_20754 n2_1458_20770 1.015873e-02
R5991 n2_1458_20770 n2_1458_20937 1.060317e-01
R5992 n2_1458_20937 n2_1458_20970 2.095238e-02
R5993 n2_1554_201 n2_1554_234 2.095238e-02
R5994 n2_1554_234 n2_1554_417 1.161905e-01
R5995 n2_1554_417 n2_1554_424 4.444444e-03
R5996 n2_1554_424 n2_1554_450 1.650794e-02
R5997 n2_1554_450 n2_1554_520 4.444444e-02
R5998 n2_1554_520 n2_1554_633 7.174603e-02
R5999 n2_1554_633 n2_1554_666 2.095238e-02
R6000 n2_1554_666 n2_1554_849 1.161905e-01
R6001 n2_1554_849 n2_1554_882 2.095238e-02
R6002 n2_1554_882 n2_1554_1065 1.161905e-01
R6003 n2_1554_1065 n2_1554_1098 2.095238e-02
R6004 n2_1554_1098 n2_1554_1281 1.161905e-01
R6005 n2_1554_1281 n2_1554_1314 2.095238e-02
R6006 n2_1554_1314 n2_1554_1497 1.161905e-01
R6007 n2_1554_1713 n2_1554_1746 2.095238e-02
R6008 n2_1554_1746 n2_1554_1760 8.888889e-03
R6009 n2_1554_1760 n2_1554_1929 1.073016e-01
R6010 n2_1554_1929 n2_1554_1962 2.095238e-02
R6011 n2_1554_1962 n2_1554_2145 1.161905e-01
R6012 n2_1554_2145 n2_1554_2178 2.095238e-02
R6013 n2_1554_2178 n2_1554_2361 1.161905e-01
R6014 n2_1554_2361 n2_1554_2394 2.095238e-02
R6015 n2_1554_2394 n2_1554_2577 1.161905e-01
R6016 n2_1554_2577 n2_1554_2610 2.095238e-02
R6017 n2_1554_2826 n2_1554_3009 1.161905e-01
R6018 n2_1554_3009 n2_1554_3042 2.095238e-02
R6019 n2_1554_3042 n2_1554_3225 1.161905e-01
R6020 n2_1554_3225 n2_1554_3258 2.095238e-02
R6021 n2_1554_3258 n2_1554_3272 8.888889e-03
R6022 n2_1554_3272 n2_1554_3441 1.073016e-01
R6023 n2_1554_3441 n2_1554_3474 2.095238e-02
R6024 n2_1554_3474 n2_1554_3657 1.161905e-01
R6025 n2_1554_3657 n2_1554_3690 2.095238e-02
R6026 n2_1554_3690 n2_1554_3704 8.888889e-03
R6027 n2_1554_3704 n2_1554_3799 6.031746e-02
R6028 n2_1554_3799 n2_1554_3873 4.698413e-02
R6029 n2_1554_3873 n2_1554_3895 1.396825e-02
R6030 n2_1554_3895 n2_1554_3906 6.984127e-03
R6031 n2_1554_3906 n2_1554_3920 8.888889e-03
R6032 n2_1554_3920 n2_1554_4089 1.073016e-01
R6033 n2_1554_4089 n2_1554_4122 2.095238e-02
R6034 n2_1554_4122 n2_1554_4159 2.349206e-02
R6035 n2_1554_4159 n2_1554_4305 9.269841e-02
R6036 n2_1554_4305 n2_1554_4338 2.095238e-02
R6037 n2_1554_4338 n2_1554_4352 8.888889e-03
R6038 n2_1554_4352 n2_1554_4375 1.460317e-02
R6039 n2_1554_4375 n2_1554_4521 9.269841e-02
R6040 n2_1554_4521 n2_1554_4554 2.095238e-02
R6041 n2_1554_4554 n2_1554_4737 1.161905e-01
R6042 n2_1554_4737 n2_1554_4770 2.095238e-02
R6043 n2_1554_5169 n2_1554_5202 2.095238e-02
R6044 n2_1554_5202 n2_1554_5385 1.161905e-01
R6045 n2_1554_5385 n2_1554_5418 2.095238e-02
R6046 n2_1554_5418 n2_1554_5432 8.888889e-03
R6047 n2_1554_5432 n2_1554_5534 6.476190e-02
R6048 n2_1554_5534 n2_1554_5601 4.253968e-02
R6049 n2_1554_5601 n2_1554_5634 2.095238e-02
R6050 n2_1554_5634 n2_1554_5817 1.161905e-01
R6051 n2_1554_5817 n2_1554_5850 2.095238e-02
R6052 n2_1554_5850 n2_1554_6033 1.161905e-01
R6053 n2_1554_6033 n2_1554_6049 1.015873e-02
R6054 n2_1554_6049 n2_1554_6066 1.079365e-02
R6055 n2_1554_6066 n2_1554_6145 5.015873e-02
R6056 n2_1554_6145 n2_1554_6249 6.603175e-02
R6057 n2_1554_6249 n2_1554_6282 2.095238e-02
R6058 n2_1554_6282 n2_1554_6465 1.161905e-01
R6059 n2_1554_6465 n2_1554_6498 2.095238e-02
R6060 n2_1554_6498 n2_1554_6535 2.349206e-02
R6061 n2_1554_6535 n2_1554_6681 9.269841e-02
R6062 n2_1554_6681 n2_1554_6714 2.095238e-02
R6063 n2_1554_6714 n2_1554_6897 1.161905e-01
R6064 n2_1554_6897 n2_1554_6930 2.095238e-02
R6065 n2_1554_6930 n2_1554_7113 1.161905e-01
R6066 n2_1554_7329 n2_1554_7362 2.095238e-02
R6067 n2_1554_7362 n2_1554_7545 1.161905e-01
R6068 n2_1554_7545 n2_1554_7578 2.095238e-02
R6069 n2_1554_7578 n2_1554_7761 1.161905e-01
R6070 n2_1554_7761 n2_1554_7794 2.095238e-02
R6071 n2_1554_7794 n2_1554_7808 8.888889e-03
R6072 n2_1554_7808 n2_1554_7977 1.073016e-01
R6073 n2_1554_7977 n2_1554_8010 2.095238e-02
R6074 n2_1554_8010 n2_1554_8193 1.161905e-01
R6075 n2_1554_8193 n2_1554_8226 2.095238e-02
R6076 n2_1554_8226 n2_1554_8299 4.634921e-02
R6077 n2_1554_8299 n2_1554_8395 6.095238e-02
R6078 n2_1554_8395 n2_1554_8409 8.888889e-03
R6079 n2_1554_8409 n2_1554_8442 2.095238e-02
R6080 n2_1554_8442 n2_1554_8625 1.161905e-01
R6081 n2_1554_8625 n2_1554_8658 2.095238e-02
R6082 n2_1554_8658 n2_1554_8841 1.161905e-01
R6083 n2_1554_8841 n2_1554_8874 2.095238e-02
R6084 n2_1554_8874 n2_1554_8888 8.888889e-03
R6085 n2_1554_8888 n2_1554_8911 1.460317e-02
R6086 n2_1554_8911 n2_1554_9057 9.269841e-02
R6087 n2_1554_9057 n2_1554_9090 2.095238e-02
R6088 n2_1554_9090 n2_1554_9273 1.161905e-01
R6089 n2_1554_9273 n2_1554_9306 2.095238e-02
R6090 n2_1554_9705 n2_1554_9738 2.095238e-02
R6091 n2_1554_9738 n2_1554_9921 1.161905e-01
R6092 n2_1554_9921 n2_1554_9954 2.095238e-02
R6093 n2_1554_9954 n2_1554_9968 8.888889e-03
R6094 n2_1554_9968 n2_1554_10137 1.073016e-01
R6095 n2_1554_10137 n2_1554_10170 2.095238e-02
R6096 n2_1554_10170 n2_1554_10353 1.161905e-01
R6097 n2_1554_10353 n2_1554_10386 2.095238e-02
R6098 n2_1554_10386 n2_1554_10549 1.034921e-01
R6099 n2_1554_10549 n2_1554_10569 1.269841e-02
R6100 n2_1554_10569 n2_1554_10602 2.095238e-02
R6101 n2_1554_10602 n2_1554_10645 2.730159e-02
R6102 n2_1554_10645 n2_1554_10785 8.888889e-02
R6103 n2_1554_10785 n2_1554_10818 2.095238e-02
R6104 n2_1554_10818 n2_1554_11001 1.161905e-01
R6105 n2_1554_11001 n2_1554_11034 2.095238e-02
R6106 n2_1554_11034 n2_1554_11048 8.888889e-03
R6107 n2_1554_11048 n2_1554_11071 1.460317e-02
R6108 n2_1554_11071 n2_1554_11217 9.269841e-02
R6109 n2_1554_11217 n2_1554_11250 2.095238e-02
R6110 n2_1554_11250 n2_1554_11433 1.161905e-01
R6111 n2_1554_11433 n2_1554_11466 2.095238e-02
R6112 n2_1554_11865 n2_1554_11898 2.095238e-02
R6113 n2_1554_11898 n2_1554_12081 1.161905e-01
R6114 n2_1554_12081 n2_1554_12114 2.095238e-02
R6115 n2_1554_12114 n2_1554_12128 8.888889e-03
R6116 n2_1554_12128 n2_1554_12297 1.073016e-01
R6117 n2_1554_12297 n2_1554_12330 2.095238e-02
R6118 n2_1554_12330 n2_1554_12513 1.161905e-01
R6119 n2_1554_12513 n2_1554_12546 2.095238e-02
R6120 n2_1554_12546 n2_1554_12729 1.161905e-01
R6121 n2_1554_12729 n2_1554_12762 2.095238e-02
R6122 n2_1554_12762 n2_1554_12799 2.349206e-02
R6123 n2_1554_12799 n2_1554_12895 6.095238e-02
R6124 n2_1554_12895 n2_1554_12945 3.174603e-02
R6125 n2_1554_12945 n2_1554_12978 2.095238e-02
R6126 n2_1554_12978 n2_1554_13161 1.161905e-01
R6127 n2_1554_13161 n2_1554_13194 2.095238e-02
R6128 n2_1554_13194 n2_1554_13377 1.161905e-01
R6129 n2_1554_13377 n2_1554_13410 2.095238e-02
R6130 n2_1554_13410 n2_1554_13447 2.349206e-02
R6131 n2_1554_13447 n2_1554_13593 9.269841e-02
R6132 n2_1554_13593 n2_1554_13626 2.095238e-02
R6133 n2_1554_13626 n2_1554_13663 2.349206e-02
R6134 n2_1554_13663 n2_1554_13809 9.269841e-02
R6135 n2_1554_13809 n2_1554_13842 2.095238e-02
R6136 n2_1554_14241 n2_1554_14274 2.095238e-02
R6137 n2_1554_14274 n2_1554_14457 1.161905e-01
R6138 n2_1554_14457 n2_1554_14490 2.095238e-02
R6139 n2_1554_14490 n2_1554_14504 8.888889e-03
R6140 n2_1554_14504 n2_1554_14673 1.073016e-01
R6141 n2_1554_14673 n2_1554_14706 2.095238e-02
R6142 n2_1554_14706 n2_1554_14889 1.161905e-01
R6143 n2_1554_14889 n2_1554_14922 2.095238e-02
R6144 n2_1554_14922 n2_1554_15049 8.063492e-02
R6145 n2_1554_15049 n2_1554_15105 3.555556e-02
R6146 n2_1554_15105 n2_1554_15138 2.095238e-02
R6147 n2_1554_15138 n2_1554_15145 4.444444e-03
R6148 n2_1554_15145 n2_1554_15321 1.117460e-01
R6149 n2_1554_15321 n2_1554_15354 2.095238e-02
R6150 n2_1554_15354 n2_1554_15368 8.888889e-03
R6151 n2_1554_15368 n2_1554_15537 1.073016e-01
R6152 n2_1554_15537 n2_1554_15570 2.095238e-02
R6153 n2_1554_15570 n2_1554_15753 1.161905e-01
R6154 n2_1554_15753 n2_1554_15786 2.095238e-02
R6155 n2_1554_15786 n2_1554_15969 1.161905e-01
R6156 n2_1554_15969 n2_1554_16002 2.095238e-02
R6157 n2_1554_16401 n2_1554_16434 2.095238e-02
R6158 n2_1554_16434 n2_1554_16471 2.349206e-02
R6159 n2_1554_16471 n2_1554_16617 9.269841e-02
R6160 n2_1554_16617 n2_1554_16650 2.095238e-02
R6161 n2_1554_16650 n2_1554_16687 2.349206e-02
R6162 n2_1554_16687 n2_1554_16833 9.269841e-02
R6163 n2_1554_16833 n2_1554_16866 2.095238e-02
R6164 n2_1554_16866 n2_1554_16880 8.888889e-03
R6165 n2_1554_16880 n2_1554_17049 1.073016e-01
R6166 n2_1554_17049 n2_1554_17082 2.095238e-02
R6167 n2_1554_17082 n2_1554_17265 1.161905e-01
R6168 n2_1554_17265 n2_1554_17298 2.095238e-02
R6169 n2_1554_17298 n2_1554_17299 6.349206e-04
R6170 n2_1554_17299 n2_1554_17395 6.095238e-02
R6171 n2_1554_17395 n2_1554_17481 5.460317e-02
R6172 n2_1554_17481 n2_1554_17514 2.095238e-02
R6173 n2_1554_17514 n2_1554_17528 8.888889e-03
R6174 n2_1554_17528 n2_1554_17697 1.073016e-01
R6175 n2_1554_17697 n2_1554_17730 2.095238e-02
R6176 n2_1554_17730 n2_1554_17913 1.161905e-01
R6177 n2_1554_17913 n2_1554_17946 2.095238e-02
R6178 n2_1554_17946 n2_1554_17960 8.888889e-03
R6179 n2_1554_17960 n2_1554_18129 1.073016e-01
R6180 n2_1554_18129 n2_1554_18162 2.095238e-02
R6181 n2_1554_18162 n2_1554_18345 1.161905e-01
R6182 n2_1554_18594 n2_1554_18777 1.161905e-01
R6183 n2_1554_18777 n2_1554_18810 2.095238e-02
R6184 n2_1554_18810 n2_1554_18993 1.161905e-01
R6185 n2_1554_18993 n2_1554_19026 2.095238e-02
R6186 n2_1554_19026 n2_1554_19040 8.888889e-03
R6187 n2_1554_19040 n2_1554_19209 1.073016e-01
R6188 n2_1554_19209 n2_1554_19242 2.095238e-02
R6189 n2_1554_19242 n2_1554_19256 8.888889e-03
R6190 n2_1554_19256 n2_1554_19425 1.073016e-01
R6191 n2_1554_19425 n2_1554_19458 2.095238e-02
R6192 n2_1554_19458 n2_1554_19472 8.888889e-03
R6193 n2_1554_19857 n2_1554_19890 2.095238e-02
R6194 n2_1554_19890 n2_1554_20073 1.161905e-01
R6195 n2_1554_20073 n2_1554_20106 2.095238e-02
R6196 n2_1554_20106 n2_1554_20289 1.161905e-01
R6197 n2_1554_20289 n2_1554_20322 2.095238e-02
R6198 n2_1554_20322 n2_1554_20505 1.161905e-01
R6199 n2_1554_20505 n2_1554_20538 2.095238e-02
R6200 n2_1554_20538 n2_1554_20674 8.634921e-02
R6201 n2_1554_20674 n2_1554_20721 2.984127e-02
R6202 n2_1554_20721 n2_1554_20754 2.095238e-02
R6203 n2_1554_20754 n2_1554_20770 1.015873e-02
R6204 n2_1554_20770 n2_1554_20937 1.060317e-01
R6205 n2_1554_20937 n2_1554_20970 2.095238e-02
R6206 n2_1646_201 n2_1646_234 2.095238e-02
R6207 n2_1646_234 n2_1646_417 1.161905e-01
R6208 n2_1646_417 n2_1646_424 4.444444e-03
R6209 n2_1646_424 n2_1646_450 1.650794e-02
R6210 n2_1646_520 n2_1646_633 7.174603e-02
R6211 n2_1646_633 n2_1646_666 2.095238e-02
R6212 n2_1646_666 n2_1646_849 1.161905e-01
R6213 n2_1646_849 n2_1646_882 2.095238e-02
R6214 n2_1646_882 n2_1646_1065 1.161905e-01
R6215 n2_1646_1065 n2_1646_1098 2.095238e-02
R6216 n2_1646_1098 n2_1646_1281 1.161905e-01
R6217 n2_1646_1281 n2_1646_1314 2.095238e-02
R6218 n2_1646_1314 n2_1646_1497 1.161905e-01
R6219 n2_1646_1497 n2_1646_1530 2.095238e-02
R6220 n2_1646_19641 n2_1646_19674 2.095238e-02
R6221 n2_1646_19674 n2_1646_19857 1.161905e-01
R6222 n2_1646_19857 n2_1646_19890 2.095238e-02
R6223 n2_1646_19890 n2_1646_20073 1.161905e-01
R6224 n2_1646_20073 n2_1646_20106 2.095238e-02
R6225 n2_1646_20106 n2_1646_20289 1.161905e-01
R6226 n2_1646_20289 n2_1646_20322 2.095238e-02
R6227 n2_1646_20322 n2_1646_20505 1.161905e-01
R6228 n2_1646_20505 n2_1646_20538 2.095238e-02
R6229 n2_1646_20538 n2_1646_20674 8.634921e-02
R6230 n2_1646_20754 n2_1646_20770 1.015873e-02
R6231 n2_1646_20770 n2_1646_20937 1.060317e-01
R6232 n2_1646_20937 n2_1646_20970 2.095238e-02
R6233 n2_2491_2793 n2_2491_2826 2.095238e-02
R6234 n2_2491_2826 n2_2491_3009 1.161905e-01
R6235 n2_2491_3009 n2_2491_3042 2.095238e-02
R6236 n2_2491_3042 n2_2491_3225 1.161905e-01
R6237 n2_2491_3225 n2_2491_3258 2.095238e-02
R6238 n2_2491_3258 n2_2491_3272 8.888889e-03
R6239 n2_2491_3272 n2_2491_3441 1.073016e-01
R6240 n2_2491_3441 n2_2491_3474 2.095238e-02
R6241 n2_2491_3474 n2_2491_3657 1.161905e-01
R6242 n2_2491_3657 n2_2491_3690 2.095238e-02
R6243 n2_2491_3690 n2_2491_3704 8.888889e-03
R6244 n2_2491_3704 n2_2491_3799 6.031746e-02
R6245 n2_2491_3873 n2_2491_3895 1.396825e-02
R6246 n2_2491_3895 n2_2491_3906 6.984127e-03
R6247 n2_2491_3906 n2_2491_3920 8.888889e-03
R6248 n2_2491_3920 n2_2491_4089 1.073016e-01
R6249 n2_2491_4089 n2_2491_4122 2.095238e-02
R6250 n2_2491_4122 n2_2491_4159 2.349206e-02
R6251 n2_2491_4159 n2_2491_4305 9.269841e-02
R6252 n2_2491_4305 n2_2491_4338 2.095238e-02
R6253 n2_2491_4338 n2_2491_4352 8.888889e-03
R6254 n2_2491_4352 n2_2491_4521 1.073016e-01
R6255 n2_2491_4521 n2_2491_4554 2.095238e-02
R6256 n2_2491_4554 n2_2491_4737 1.161905e-01
R6257 n2_2491_4737 n2_2491_4770 2.095238e-02
R6258 n2_2491_4770 n2_2491_4953 1.161905e-01
R6259 n2_2491_4953 n2_2491_4986 2.095238e-02
R6260 n2_2491_4986 n2_2491_5169 1.161905e-01
R6261 n2_2491_5169 n2_2491_5202 2.095238e-02
R6262 n2_2491_5202 n2_2491_5385 1.161905e-01
R6263 n2_2491_5385 n2_2491_5418 2.095238e-02
R6264 n2_2491_5418 n2_2491_5432 8.888889e-03
R6265 n2_2491_5432 n2_2491_5601 1.073016e-01
R6266 n2_2491_5601 n2_2491_5634 2.095238e-02
R6267 n2_2491_5634 n2_2491_5817 1.161905e-01
R6268 n2_2491_5817 n2_2491_5850 2.095238e-02
R6269 n2_2491_5850 n2_2491_6033 1.161905e-01
R6270 n2_2491_6033 n2_2491_6049 1.015873e-02
R6271 n2_2491_6049 n2_2491_6066 1.079365e-02
R6272 n2_2491_6145 n2_2491_6249 6.603175e-02
R6273 n2_2491_6249 n2_2491_6282 2.095238e-02
R6274 n2_2491_6282 n2_2491_6465 1.161905e-01
R6275 n2_2491_6465 n2_2491_6498 2.095238e-02
R6276 n2_2491_6498 n2_2491_6535 2.349206e-02
R6277 n2_2491_6535 n2_2491_6681 9.269841e-02
R6278 n2_2491_6681 n2_2491_6714 2.095238e-02
R6279 n2_2491_6714 n2_2491_6897 1.161905e-01
R6280 n2_2491_6897 n2_2491_6930 2.095238e-02
R6281 n2_2491_6930 n2_2491_7113 1.161905e-01
R6282 n2_2491_7113 n2_2491_7146 2.095238e-02
R6283 n2_2491_7146 n2_2491_7329 1.161905e-01
R6284 n2_2491_7329 n2_2491_7362 2.095238e-02
R6285 n2_2491_7362 n2_2491_7545 1.161905e-01
R6286 n2_2491_7545 n2_2491_7578 2.095238e-02
R6287 n2_2491_7578 n2_2491_7761 1.161905e-01
R6288 n2_2491_7761 n2_2491_7794 2.095238e-02
R6289 n2_2491_7794 n2_2491_7808 8.888889e-03
R6290 n2_2491_7808 n2_2491_7977 1.073016e-01
R6291 n2_2491_7977 n2_2491_8010 2.095238e-02
R6292 n2_2491_8010 n2_2491_8193 1.161905e-01
R6293 n2_2491_8193 n2_2491_8226 2.095238e-02
R6294 n2_2491_8226 n2_2491_8299 4.634921e-02
R6295 n2_2491_8395 n2_2491_8409 8.888889e-03
R6296 n2_2491_8409 n2_2491_8442 2.095238e-02
R6297 n2_2491_8442 n2_2491_8625 1.161905e-01
R6298 n2_2491_8625 n2_2491_8658 2.095238e-02
R6299 n2_2491_8658 n2_2491_8841 1.161905e-01
R6300 n2_2491_8841 n2_2491_8874 2.095238e-02
R6301 n2_2491_8874 n2_2491_8888 8.888889e-03
R6302 n2_2491_8888 n2_2491_8911 1.460317e-02
R6303 n2_2491_8911 n2_2491_9057 9.269841e-02
R6304 n2_2491_9057 n2_2491_9090 2.095238e-02
R6305 n2_2491_9090 n2_2491_9273 1.161905e-01
R6306 n2_2491_9273 n2_2491_9306 2.095238e-02
R6307 n2_2491_9306 n2_2491_9489 1.161905e-01
R6308 n2_2491_9489 n2_2491_9522 2.095238e-02
R6309 n2_2491_9522 n2_2491_9705 1.161905e-01
R6310 n2_2491_9705 n2_2491_9738 2.095238e-02
R6311 n2_2491_9738 n2_2491_9921 1.161905e-01
R6312 n2_2491_9921 n2_2491_9954 2.095238e-02
R6313 n2_2491_9954 n2_2491_9968 8.888889e-03
R6314 n2_2491_9968 n2_2491_10137 1.073016e-01
R6315 n2_2491_10137 n2_2491_10170 2.095238e-02
R6316 n2_2491_10170 n2_2491_10353 1.161905e-01
R6317 n2_2491_10353 n2_2491_10386 2.095238e-02
R6318 n2_2491_10386 n2_2491_10549 1.034921e-01
R6319 n2_2491_10549 n2_2491_10569 1.269841e-02
R6320 n2_2491_10645 n2_2491_10785 8.888889e-02
R6321 n2_2491_10785 n2_2491_10818 2.095238e-02
R6322 n2_2491_10818 n2_2491_11001 1.161905e-01
R6323 n2_2491_11001 n2_2491_11034 2.095238e-02
R6324 n2_2491_11034 n2_2491_11048 8.888889e-03
R6325 n2_2491_11048 n2_2491_11071 1.460317e-02
R6326 n2_2491_11071 n2_2491_11217 9.269841e-02
R6327 n2_2491_11217 n2_2491_11250 2.095238e-02
R6328 n2_2491_11250 n2_2491_11433 1.161905e-01
R6329 n2_2491_11433 n2_2491_11466 2.095238e-02
R6330 n2_2491_11466 n2_2491_11649 1.161905e-01
R6331 n2_2491_11649 n2_2491_11682 2.095238e-02
R6332 n2_2491_11682 n2_2491_11865 1.161905e-01
R6333 n2_2491_11865 n2_2491_11898 2.095238e-02
R6334 n2_2491_11898 n2_2491_12081 1.161905e-01
R6335 n2_2491_12081 n2_2491_12114 2.095238e-02
R6336 n2_2491_12114 n2_2491_12128 8.888889e-03
R6337 n2_2491_12128 n2_2491_12151 1.460317e-02
R6338 n2_2491_12151 n2_2491_12297 9.269841e-02
R6339 n2_2491_12297 n2_2491_12330 2.095238e-02
R6340 n2_2491_12330 n2_2491_12513 1.161905e-01
R6341 n2_2491_12513 n2_2491_12546 2.095238e-02
R6342 n2_2491_12546 n2_2491_12729 1.161905e-01
R6343 n2_2491_12729 n2_2491_12762 2.095238e-02
R6344 n2_2491_12762 n2_2491_12799 2.349206e-02
R6345 n2_2491_12895 n2_2491_12945 3.174603e-02
R6346 n2_2491_12945 n2_2491_12978 2.095238e-02
R6347 n2_2491_12978 n2_2491_13161 1.161905e-01
R6348 n2_2491_13161 n2_2491_13194 2.095238e-02
R6349 n2_2491_13194 n2_2491_13377 1.161905e-01
R6350 n2_2491_13377 n2_2491_13410 2.095238e-02
R6351 n2_2491_13410 n2_2491_13424 8.888889e-03
R6352 n2_2491_13424 n2_2491_13447 1.460317e-02
R6353 n2_2491_13447 n2_2491_13593 9.269841e-02
R6354 n2_2491_13593 n2_2491_13626 2.095238e-02
R6355 n2_2491_13626 n2_2491_13640 8.888889e-03
R6356 n2_2491_13640 n2_2491_13809 1.073016e-01
R6357 n2_2491_13809 n2_2491_13842 2.095238e-02
R6358 n2_2491_13842 n2_2491_13879 2.349206e-02
R6359 n2_2491_13879 n2_2491_14025 9.269841e-02
R6360 n2_2491_14025 n2_2491_14058 2.095238e-02
R6361 n2_2491_14058 n2_2491_14100 2.666667e-02
R6362 n2_2491_14100 n2_2491_14241 8.952381e-02
R6363 n2_2491_14241 n2_2491_14274 2.095238e-02
R6364 n2_2491_14274 n2_2491_14457 1.161905e-01
R6365 n2_2491_14457 n2_2491_14490 2.095238e-02
R6366 n2_2491_14490 n2_2491_14504 8.888889e-03
R6367 n2_2491_14504 n2_2491_14536 2.031746e-02
R6368 n2_2491_14536 n2_2491_14673 8.698413e-02
R6369 n2_2491_14673 n2_2491_14706 2.095238e-02
R6370 n2_2491_14706 n2_2491_14889 1.161905e-01
R6371 n2_2491_14889 n2_2491_14922 2.095238e-02
R6372 n2_2491_14922 n2_2491_15049 8.063492e-02
R6373 n2_2491_15138 n2_2491_15145 4.444444e-03
R6374 n2_2491_15145 n2_2491_15321 1.117460e-01
R6375 n2_2491_15321 n2_2491_15354 2.095238e-02
R6376 n2_2491_15354 n2_2491_15368 8.888889e-03
R6377 n2_2491_15368 n2_2491_15537 1.073016e-01
R6378 n2_2491_15537 n2_2491_15570 2.095238e-02
R6379 n2_2491_15570 n2_2491_15584 8.888889e-03
R6380 n2_2491_15584 n2_2491_15753 1.073016e-01
R6381 n2_2491_15753 n2_2491_15786 2.095238e-02
R6382 n2_2491_15786 n2_2491_15969 1.161905e-01
R6383 n2_2491_15969 n2_2491_16002 2.095238e-02
R6384 n2_2491_16002 n2_2491_16185 1.161905e-01
R6385 n2_2491_16185 n2_2491_16218 2.095238e-02
R6386 n2_2491_16218 n2_2491_16401 1.161905e-01
R6387 n2_2491_16401 n2_2491_16434 2.095238e-02
R6388 n2_2491_16434 n2_2491_16471 2.349206e-02
R6389 n2_2491_16471 n2_2491_16617 9.269841e-02
R6390 n2_2491_16617 n2_2491_16650 2.095238e-02
R6391 n2_2491_16650 n2_2491_16664 8.888889e-03
R6392 n2_2491_16664 n2_2491_16687 1.460317e-02
R6393 n2_2491_16687 n2_2491_16833 9.269841e-02
R6394 n2_2491_16833 n2_2491_16866 2.095238e-02
R6395 n2_2491_16866 n2_2491_16880 8.888889e-03
R6396 n2_2491_16880 n2_2491_17049 1.073016e-01
R6397 n2_2491_17049 n2_2491_17082 2.095238e-02
R6398 n2_2491_17082 n2_2491_17265 1.161905e-01
R6399 n2_2491_17265 n2_2491_17298 2.095238e-02
R6400 n2_2491_17298 n2_2491_17299 6.349206e-04
R6401 n2_2491_17395 n2_2491_17481 5.460317e-02
R6402 n2_2491_17481 n2_2491_17514 2.095238e-02
R6403 n2_2491_17514 n2_2491_17528 8.888889e-03
R6404 n2_2491_17528 n2_2491_17551 1.460317e-02
R6405 n2_2491_17551 n2_2491_17697 9.269841e-02
R6406 n2_2491_17697 n2_2491_17730 2.095238e-02
R6407 n2_2491_17730 n2_2491_17913 1.161905e-01
R6408 n2_2491_17913 n2_2491_17946 2.095238e-02
R6409 n2_2491_17946 n2_2491_17960 8.888889e-03
R6410 n2_2491_17960 n2_2491_18129 1.073016e-01
R6411 n2_2491_18129 n2_2491_18162 2.095238e-02
R6412 n2_2491_18162 n2_2491_18345 1.161905e-01
R6413 n2_2491_18345 n2_2491_18378 2.095238e-02
R6414 n2_2491_3799 n2_2630_3799 8.825397e-02
R6415 n2_2630_3799 n2_2679_3799 3.111111e-02
R6416 n2_2491_3895 n2_2630_3895 8.825397e-02
R6417 n2_2630_3895 n2_2679_3895 3.111111e-02
R6418 n2_2491_6049 n2_2630_6049 8.825397e-02
R6419 n2_2630_6049 n2_2679_6049 3.111111e-02
R6420 n2_2491_6145 n2_2630_6145 8.825397e-02
R6421 n2_2630_6145 n2_2679_6145 3.111111e-02
R6422 n2_2491_8299 n2_2630_8299 8.825397e-02
R6423 n2_2630_8299 n2_2679_8299 3.111111e-02
R6424 n2_2491_8395 n2_2630_8395 8.825397e-02
R6425 n2_2630_8395 n2_2679_8395 3.111111e-02
R6426 n2_2491_10549 n2_2630_10549 8.825397e-02
R6427 n2_2630_10549 n2_2679_10549 3.111111e-02
R6428 n2_2491_10645 n2_2630_10645 8.825397e-02
R6429 n2_2630_10645 n2_2679_10645 3.111111e-02
R6430 n2_2491_12799 n2_2630_12799 8.825397e-02
R6431 n2_2630_12799 n2_2679_12799 3.111111e-02
R6432 n2_2491_12895 n2_2630_12895 8.825397e-02
R6433 n2_2630_12895 n2_2679_12895 3.111111e-02
R6434 n2_2491_15049 n2_2630_15049 8.825397e-02
R6435 n2_2630_15049 n2_2679_15049 3.111111e-02
R6436 n2_2491_15145 n2_2630_15145 8.825397e-02
R6437 n2_2630_15145 n2_2679_15145 3.111111e-02
R6438 n2_2491_17299 n2_2630_17299 8.825397e-02
R6439 n2_2630_17299 n2_2679_17299 3.111111e-02
R6440 n2_2491_17395 n2_2630_17395 8.825397e-02
R6441 n2_2630_17395 n2_2679_17395 3.111111e-02
R6442 n2_2679_2826 n2_2679_3009 1.161905e-01
R6443 n2_2679_3009 n2_2679_3042 2.095238e-02
R6444 n2_2679_3042 n2_2679_3225 1.161905e-01
R6445 n2_2679_3225 n2_2679_3258 2.095238e-02
R6446 n2_2679_3258 n2_2679_3272 8.888889e-03
R6447 n2_2679_3272 n2_2679_3441 1.073016e-01
R6448 n2_2679_3441 n2_2679_3474 2.095238e-02
R6449 n2_2679_3474 n2_2679_3657 1.161905e-01
R6450 n2_2679_3657 n2_2679_3690 2.095238e-02
R6451 n2_2679_3690 n2_2679_3704 8.888889e-03
R6452 n2_2679_3704 n2_2679_3799 6.031746e-02
R6453 n2_2679_3799 n2_2679_3873 4.698413e-02
R6454 n2_2679_3873 n2_2679_3895 1.396825e-02
R6455 n2_2679_3895 n2_2679_3906 6.984127e-03
R6456 n2_2679_3906 n2_2679_3920 8.888889e-03
R6457 n2_2679_3920 n2_2679_4089 1.073016e-01
R6458 n2_2679_4089 n2_2679_4122 2.095238e-02
R6459 n2_2679_4122 n2_2679_4159 2.349206e-02
R6460 n2_2679_4159 n2_2679_4305 9.269841e-02
R6461 n2_2679_4305 n2_2679_4338 2.095238e-02
R6462 n2_2679_4338 n2_2679_4352 8.888889e-03
R6463 n2_2679_4352 n2_2679_4521 1.073016e-01
R6464 n2_2679_4521 n2_2679_4554 2.095238e-02
R6465 n2_2679_4554 n2_2679_4737 1.161905e-01
R6466 n2_2679_4737 n2_2679_4770 2.095238e-02
R6467 n2_2679_5169 n2_2679_5202 2.095238e-02
R6468 n2_2679_5202 n2_2679_5385 1.161905e-01
R6469 n2_2679_5385 n2_2679_5418 2.095238e-02
R6470 n2_2679_5418 n2_2679_5432 8.888889e-03
R6471 n2_2679_5432 n2_2679_5601 1.073016e-01
R6472 n2_2679_5601 n2_2679_5634 2.095238e-02
R6473 n2_2679_5634 n2_2679_5817 1.161905e-01
R6474 n2_2679_5817 n2_2679_5850 2.095238e-02
R6475 n2_2679_5850 n2_2679_6033 1.161905e-01
R6476 n2_2679_6033 n2_2679_6049 1.015873e-02
R6477 n2_2679_6049 n2_2679_6066 1.079365e-02
R6478 n2_2679_6066 n2_2679_6145 5.015873e-02
R6479 n2_2679_6145 n2_2679_6249 6.603175e-02
R6480 n2_2679_6249 n2_2679_6282 2.095238e-02
R6481 n2_2679_6282 n2_2679_6465 1.161905e-01
R6482 n2_2679_6465 n2_2679_6498 2.095238e-02
R6483 n2_2679_6498 n2_2679_6535 2.349206e-02
R6484 n2_2679_6535 n2_2679_6681 9.269841e-02
R6485 n2_2679_6681 n2_2679_6714 2.095238e-02
R6486 n2_2679_6714 n2_2679_6897 1.161905e-01
R6487 n2_2679_6897 n2_2679_6930 2.095238e-02
R6488 n2_2679_6930 n2_2679_7113 1.161905e-01
R6489 n2_2679_7329 n2_2679_7362 2.095238e-02
R6490 n2_2679_7362 n2_2679_7545 1.161905e-01
R6491 n2_2679_7545 n2_2679_7578 2.095238e-02
R6492 n2_2679_7578 n2_2679_7761 1.161905e-01
R6493 n2_2679_7761 n2_2679_7794 2.095238e-02
R6494 n2_2679_7794 n2_2679_7808 8.888889e-03
R6495 n2_2679_7808 n2_2679_7977 1.073016e-01
R6496 n2_2679_7977 n2_2679_8010 2.095238e-02
R6497 n2_2679_8010 n2_2679_8193 1.161905e-01
R6498 n2_2679_8193 n2_2679_8226 2.095238e-02
R6499 n2_2679_8226 n2_2679_8299 4.634921e-02
R6500 n2_2679_8299 n2_2679_8395 6.095238e-02
R6501 n2_2679_8395 n2_2679_8409 8.888889e-03
R6502 n2_2679_8409 n2_2679_8442 2.095238e-02
R6503 n2_2679_8442 n2_2679_8625 1.161905e-01
R6504 n2_2679_8625 n2_2679_8658 2.095238e-02
R6505 n2_2679_8658 n2_2679_8841 1.161905e-01
R6506 n2_2679_8841 n2_2679_8874 2.095238e-02
R6507 n2_2679_8874 n2_2679_8888 8.888889e-03
R6508 n2_2679_8888 n2_2679_8911 1.460317e-02
R6509 n2_2679_8911 n2_2679_9057 9.269841e-02
R6510 n2_2679_9057 n2_2679_9090 2.095238e-02
R6511 n2_2679_9090 n2_2679_9273 1.161905e-01
R6512 n2_2679_9273 n2_2679_9306 2.095238e-02
R6513 n2_2679_9705 n2_2679_9738 2.095238e-02
R6514 n2_2679_9738 n2_2679_9921 1.161905e-01
R6515 n2_2679_9921 n2_2679_9954 2.095238e-02
R6516 n2_2679_9954 n2_2679_9968 8.888889e-03
R6517 n2_2679_9968 n2_2679_10137 1.073016e-01
R6518 n2_2679_10137 n2_2679_10170 2.095238e-02
R6519 n2_2679_10170 n2_2679_10353 1.161905e-01
R6520 n2_2679_10353 n2_2679_10386 2.095238e-02
R6521 n2_2679_10386 n2_2679_10549 1.034921e-01
R6522 n2_2679_10549 n2_2679_10569 1.269841e-02
R6523 n2_2679_10569 n2_2679_10602 2.095238e-02
R6524 n2_2679_10602 n2_2679_10645 2.730159e-02
R6525 n2_2679_10645 n2_2679_10785 8.888889e-02
R6526 n2_2679_10785 n2_2679_10818 2.095238e-02
R6527 n2_2679_10818 n2_2679_11001 1.161905e-01
R6528 n2_2679_11001 n2_2679_11034 2.095238e-02
R6529 n2_2679_11034 n2_2679_11048 8.888889e-03
R6530 n2_2679_11048 n2_2679_11071 1.460317e-02
R6531 n2_2679_11071 n2_2679_11217 9.269841e-02
R6532 n2_2679_11217 n2_2679_11250 2.095238e-02
R6533 n2_2679_11250 n2_2679_11433 1.161905e-01
R6534 n2_2679_11433 n2_2679_11466 2.095238e-02
R6535 n2_2679_11865 n2_2679_11898 2.095238e-02
R6536 n2_2679_11898 n2_2679_12081 1.161905e-01
R6537 n2_2679_12081 n2_2679_12114 2.095238e-02
R6538 n2_2679_12114 n2_2679_12128 8.888889e-03
R6539 n2_2679_12128 n2_2679_12151 1.460317e-02
R6540 n2_2679_12151 n2_2679_12297 9.269841e-02
R6541 n2_2679_12297 n2_2679_12330 2.095238e-02
R6542 n2_2679_12330 n2_2679_12513 1.161905e-01
R6543 n2_2679_12513 n2_2679_12546 2.095238e-02
R6544 n2_2679_12546 n2_2679_12729 1.161905e-01
R6545 n2_2679_12729 n2_2679_12762 2.095238e-02
R6546 n2_2679_12762 n2_2679_12799 2.349206e-02
R6547 n2_2679_12799 n2_2679_12895 6.095238e-02
R6548 n2_2679_12895 n2_2679_12945 3.174603e-02
R6549 n2_2679_12945 n2_2679_12978 2.095238e-02
R6550 n2_2679_12978 n2_2679_13161 1.161905e-01
R6551 n2_2679_13161 n2_2679_13194 2.095238e-02
R6552 n2_2679_13194 n2_2679_13377 1.161905e-01
R6553 n2_2679_13377 n2_2679_13410 2.095238e-02
R6554 n2_2679_13410 n2_2679_13424 8.888889e-03
R6555 n2_2679_13424 n2_2679_13447 1.460317e-02
R6556 n2_2679_13447 n2_2679_13593 9.269841e-02
R6557 n2_2679_13593 n2_2679_13626 2.095238e-02
R6558 n2_2679_13626 n2_2679_13640 8.888889e-03
R6559 n2_2679_13640 n2_2679_13809 1.073016e-01
R6560 n2_2679_13809 n2_2679_13842 2.095238e-02
R6561 n2_2679_14100 n2_2679_14241 8.952381e-02
R6562 n2_2679_14241 n2_2679_14274 2.095238e-02
R6563 n2_2679_14274 n2_2679_14457 1.161905e-01
R6564 n2_2679_14457 n2_2679_14490 2.095238e-02
R6565 n2_2679_14490 n2_2679_14504 8.888889e-03
R6566 n2_2679_14504 n2_2679_14536 2.031746e-02
R6567 n2_2679_14536 n2_2679_14673 8.698413e-02
R6568 n2_2679_14673 n2_2679_14706 2.095238e-02
R6569 n2_2679_14706 n2_2679_14889 1.161905e-01
R6570 n2_2679_14889 n2_2679_14922 2.095238e-02
R6571 n2_2679_14922 n2_2679_15049 8.063492e-02
R6572 n2_2679_15049 n2_2679_15105 3.555556e-02
R6573 n2_2679_15105 n2_2679_15138 2.095238e-02
R6574 n2_2679_15138 n2_2679_15145 4.444444e-03
R6575 n2_2679_15145 n2_2679_15321 1.117460e-01
R6576 n2_2679_15321 n2_2679_15354 2.095238e-02
R6577 n2_2679_15354 n2_2679_15368 8.888889e-03
R6578 n2_2679_15368 n2_2679_15537 1.073016e-01
R6579 n2_2679_15537 n2_2679_15570 2.095238e-02
R6580 n2_2679_15570 n2_2679_15584 8.888889e-03
R6581 n2_2679_15584 n2_2679_15753 1.073016e-01
R6582 n2_2679_15753 n2_2679_15786 2.095238e-02
R6583 n2_2679_15786 n2_2679_15969 1.161905e-01
R6584 n2_2679_15969 n2_2679_16002 2.095238e-02
R6585 n2_2679_16401 n2_2679_16434 2.095238e-02
R6586 n2_2679_16434 n2_2679_16471 2.349206e-02
R6587 n2_2679_16471 n2_2679_16617 9.269841e-02
R6588 n2_2679_16617 n2_2679_16650 2.095238e-02
R6589 n2_2679_16650 n2_2679_16664 8.888889e-03
R6590 n2_2679_16664 n2_2679_16687 1.460317e-02
R6591 n2_2679_16687 n2_2679_16833 9.269841e-02
R6592 n2_2679_16833 n2_2679_16866 2.095238e-02
R6593 n2_2679_16866 n2_2679_16880 8.888889e-03
R6594 n2_2679_16880 n2_2679_17049 1.073016e-01
R6595 n2_2679_17049 n2_2679_17082 2.095238e-02
R6596 n2_2679_17082 n2_2679_17265 1.161905e-01
R6597 n2_2679_17265 n2_2679_17298 2.095238e-02
R6598 n2_2679_17298 n2_2679_17299 6.349206e-04
R6599 n2_2679_17299 n2_2679_17395 6.095238e-02
R6600 n2_2679_17395 n2_2679_17481 5.460317e-02
R6601 n2_2679_17481 n2_2679_17514 2.095238e-02
R6602 n2_2679_17514 n2_2679_17528 8.888889e-03
R6603 n2_2679_17528 n2_2679_17551 1.460317e-02
R6604 n2_2679_17551 n2_2679_17697 9.269841e-02
R6605 n2_2679_17697 n2_2679_17730 2.095238e-02
R6606 n2_2679_17730 n2_2679_17913 1.161905e-01
R6607 n2_2679_17913 n2_2679_17946 2.095238e-02
R6608 n2_2679_17946 n2_2679_17960 8.888889e-03
R6609 n2_2679_17960 n2_2679_18129 1.073016e-01
R6610 n2_2679_18129 n2_2679_18162 2.095238e-02
R6611 n2_2679_18162 n2_2679_18345 1.161905e-01
R6612 n2_3616_201 n2_3616_234 2.095238e-02
R6613 n2_3616_234 n2_3616_356 7.746032e-02
R6614 n2_3616_356 n2_3616_417 3.873016e-02
R6615 n2_3616_417 n2_3616_424 4.444444e-03
R6616 n2_3616_424 n2_3616_450 1.650794e-02
R6617 n2_3616_520 n2_3616_633 7.174603e-02
R6618 n2_3616_633 n2_3616_666 2.095238e-02
R6619 n2_3616_666 n2_3616_788 7.746032e-02
R6620 n2_3616_788 n2_3616_849 3.873016e-02
R6621 n2_3616_849 n2_3616_882 2.095238e-02
R6622 n2_3616_882 n2_3616_1065 1.161905e-01
R6623 n2_3616_1065 n2_3616_1098 2.095238e-02
R6624 n2_3616_1098 n2_3616_1281 1.161905e-01
R6625 n2_3616_1281 n2_3616_1314 2.095238e-02
R6626 n2_3616_1314 n2_3616_1497 1.161905e-01
R6627 n2_3616_1497 n2_3616_1530 2.095238e-02
R6628 n2_3616_1530 n2_3616_1549 1.206349e-02
R6629 n2_3616_1645 n2_3616_1652 4.444444e-03
R6630 n2_3616_1652 n2_3616_1713 3.873016e-02
R6631 n2_3616_1713 n2_3616_1746 2.095238e-02
R6632 n2_3616_1746 n2_3616_1929 1.161905e-01
R6633 n2_3616_1929 n2_3616_1962 2.095238e-02
R6634 n2_3616_1962 n2_3616_1976 8.888889e-03
R6635 n2_3616_1976 n2_3616_2145 1.073016e-01
R6636 n2_3616_2145 n2_3616_2178 2.095238e-02
R6637 n2_3616_2178 n2_3616_2361 1.161905e-01
R6638 n2_3616_2361 n2_3616_2394 2.095238e-02
R6639 n2_3616_2394 n2_3616_2577 1.161905e-01
R6640 n2_3616_2577 n2_3616_2610 2.095238e-02
R6641 n2_3616_2610 n2_3616_2674 4.063492e-02
R6642 n2_3616_2770 n2_3616_2793 1.460317e-02
R6643 n2_3616_2793 n2_3616_2826 2.095238e-02
R6644 n2_3616_2826 n2_3616_3009 1.161905e-01
R6645 n2_3616_3009 n2_3616_3042 2.095238e-02
R6646 n2_3616_3042 n2_3616_3225 1.161905e-01
R6647 n2_3616_3225 n2_3616_3258 2.095238e-02
R6648 n2_3616_3258 n2_3616_3441 1.161905e-01
R6649 n2_3616_3441 n2_3616_3474 2.095238e-02
R6650 n2_3616_3474 n2_3616_3657 1.161905e-01
R6651 n2_3616_3657 n2_3616_3690 2.095238e-02
R6652 n2_3616_3690 n2_3616_3704 8.888889e-03
R6653 n2_3616_3704 n2_3616_3799 6.031746e-02
R6654 n2_3616_3873 n2_3616_3895 1.396825e-02
R6655 n2_3616_3895 n2_3616_3906 6.984127e-03
R6656 n2_3616_3906 n2_3616_3920 8.888889e-03
R6657 n2_3616_3920 n2_3616_4089 1.073016e-01
R6658 n2_3616_4089 n2_3616_4122 2.095238e-02
R6659 n2_3616_4122 n2_3616_4136 8.888889e-03
R6660 n2_3616_4136 n2_3616_4159 1.460317e-02
R6661 n2_3616_4159 n2_3616_4305 9.269841e-02
R6662 n2_3616_4305 n2_3616_4338 2.095238e-02
R6663 n2_3616_4338 n2_3616_4352 8.888889e-03
R6664 n2_3616_4352 n2_3616_4375 1.460317e-02
R6665 n2_3616_4375 n2_3616_4521 9.269841e-02
R6666 n2_3616_4521 n2_3616_4554 2.095238e-02
R6667 n2_3616_4554 n2_3616_4737 1.161905e-01
R6668 n2_3616_4737 n2_3616_4770 2.095238e-02
R6669 n2_3616_4770 n2_3616_4953 1.161905e-01
R6670 n2_3616_4953 n2_3616_4986 2.095238e-02
R6671 n2_3616_4986 n2_3616_5169 1.161905e-01
R6672 n2_3616_5169 n2_3616_5202 2.095238e-02
R6673 n2_3616_5202 n2_3616_5385 1.161905e-01
R6674 n2_3616_5385 n2_3616_5418 2.095238e-02
R6675 n2_3616_5418 n2_3616_5432 8.888889e-03
R6676 n2_3616_5432 n2_3616_5601 1.073016e-01
R6677 n2_3616_5601 n2_3616_5634 2.095238e-02
R6678 n2_3616_5634 n2_3616_5817 1.161905e-01
R6679 n2_3616_5817 n2_3616_5850 2.095238e-02
R6680 n2_3616_5850 n2_3616_6033 1.161905e-01
R6681 n2_3616_6033 n2_3616_6049 1.015873e-02
R6682 n2_3616_6049 n2_3616_6066 1.079365e-02
R6683 n2_3616_6145 n2_3616_6249 6.603175e-02
R6684 n2_3616_6249 n2_3616_6282 2.095238e-02
R6685 n2_3616_6282 n2_3616_6465 1.161905e-01
R6686 n2_3616_6465 n2_3616_6498 2.095238e-02
R6687 n2_3616_6498 n2_3616_6535 2.349206e-02
R6688 n2_3616_6535 n2_3616_6681 9.269841e-02
R6689 n2_3616_6681 n2_3616_6714 2.095238e-02
R6690 n2_3616_6714 n2_3616_6897 1.161905e-01
R6691 n2_3616_6897 n2_3616_6930 2.095238e-02
R6692 n2_3616_6930 n2_3616_7113 1.161905e-01
R6693 n2_3616_7113 n2_3616_7146 2.095238e-02
R6694 n2_3616_7146 n2_3616_7329 1.161905e-01
R6695 n2_3616_7329 n2_3616_7362 2.095238e-02
R6696 n2_3616_7362 n2_3616_7545 1.161905e-01
R6697 n2_3616_7545 n2_3616_7578 2.095238e-02
R6698 n2_3616_7578 n2_3616_7761 1.161905e-01
R6699 n2_3616_7761 n2_3616_7794 2.095238e-02
R6700 n2_3616_7794 n2_3616_7808 8.888889e-03
R6701 n2_3616_7808 n2_3616_7977 1.073016e-01
R6702 n2_3616_7977 n2_3616_8010 2.095238e-02
R6703 n2_3616_8010 n2_3616_8193 1.161905e-01
R6704 n2_3616_8193 n2_3616_8226 2.095238e-02
R6705 n2_3616_8226 n2_3616_8299 4.634921e-02
R6706 n2_3616_8395 n2_3616_8409 8.888889e-03
R6707 n2_3616_8409 n2_3616_8442 2.095238e-02
R6708 n2_3616_8442 n2_3616_8625 1.161905e-01
R6709 n2_3616_8625 n2_3616_8658 2.095238e-02
R6710 n2_3616_8658 n2_3616_8841 1.161905e-01
R6711 n2_3616_8841 n2_3616_8874 2.095238e-02
R6712 n2_3616_8874 n2_3616_8888 8.888889e-03
R6713 n2_3616_8888 n2_3616_8911 1.460317e-02
R6714 n2_3616_8911 n2_3616_9057 9.269841e-02
R6715 n2_3616_9057 n2_3616_9090 2.095238e-02
R6716 n2_3616_9090 n2_3616_9273 1.161905e-01
R6717 n2_3616_9273 n2_3616_9306 2.095238e-02
R6718 n2_3616_9306 n2_3616_9489 1.161905e-01
R6719 n2_3616_9489 n2_3616_9522 2.095238e-02
R6720 n2_3616_9522 n2_3616_9705 1.161905e-01
R6721 n2_3616_9705 n2_3616_9738 2.095238e-02
R6722 n2_3616_9738 n2_3616_9921 1.161905e-01
R6723 n2_3616_9921 n2_3616_9954 2.095238e-02
R6724 n2_3616_9954 n2_3616_9968 8.888889e-03
R6725 n2_3616_9968 n2_3616_10137 1.073016e-01
R6726 n2_3616_10137 n2_3616_10170 2.095238e-02
R6727 n2_3616_10170 n2_3616_10353 1.161905e-01
R6728 n2_3616_10353 n2_3616_10386 2.095238e-02
R6729 n2_3616_10386 n2_3616_10549 1.034921e-01
R6730 n2_3616_10549 n2_3616_10569 1.269841e-02
R6731 n2_3616_10645 n2_3616_10785 8.888889e-02
R6732 n2_3616_10785 n2_3616_10818 2.095238e-02
R6733 n2_3616_10818 n2_3616_11001 1.161905e-01
R6734 n2_3616_11001 n2_3616_11034 2.095238e-02
R6735 n2_3616_11034 n2_3616_11048 8.888889e-03
R6736 n2_3616_11048 n2_3616_11217 1.073016e-01
R6737 n2_3616_11217 n2_3616_11250 2.095238e-02
R6738 n2_3616_11250 n2_3616_11433 1.161905e-01
R6739 n2_3616_11433 n2_3616_11466 2.095238e-02
R6740 n2_3616_11466 n2_3616_11649 1.161905e-01
R6741 n2_3616_11649 n2_3616_11682 2.095238e-02
R6742 n2_3616_11682 n2_3616_11865 1.161905e-01
R6743 n2_3616_11865 n2_3616_11898 2.095238e-02
R6744 n2_3616_11898 n2_3616_12081 1.161905e-01
R6745 n2_3616_12081 n2_3616_12114 2.095238e-02
R6746 n2_3616_12114 n2_3616_12128 8.888889e-03
R6747 n2_3616_12128 n2_3616_12151 1.460317e-02
R6748 n2_3616_12151 n2_3616_12297 9.269841e-02
R6749 n2_3616_12297 n2_3616_12330 2.095238e-02
R6750 n2_3616_12330 n2_3616_12513 1.161905e-01
R6751 n2_3616_12513 n2_3616_12546 2.095238e-02
R6752 n2_3616_12546 n2_3616_12729 1.161905e-01
R6753 n2_3616_12729 n2_3616_12762 2.095238e-02
R6754 n2_3616_12762 n2_3616_12799 2.349206e-02
R6755 n2_3616_12895 n2_3616_12945 3.174603e-02
R6756 n2_3616_12945 n2_3616_12978 2.095238e-02
R6757 n2_3616_12978 n2_3616_13161 1.161905e-01
R6758 n2_3616_13161 n2_3616_13194 2.095238e-02
R6759 n2_3616_13194 n2_3616_13377 1.161905e-01
R6760 n2_3616_13377 n2_3616_13410 2.095238e-02
R6761 n2_3616_13410 n2_3616_13424 8.888889e-03
R6762 n2_3616_13424 n2_3616_13593 1.073016e-01
R6763 n2_3616_13593 n2_3616_13626 2.095238e-02
R6764 n2_3616_13626 n2_3616_13640 8.888889e-03
R6765 n2_3616_13640 n2_3616_13809 1.073016e-01
R6766 n2_3616_13809 n2_3616_13842 2.095238e-02
R6767 n2_3616_13842 n2_3616_13879 2.349206e-02
R6768 n2_3616_13879 n2_3616_14025 9.269841e-02
R6769 n2_3616_14025 n2_3616_14058 2.095238e-02
R6770 n2_3616_14058 n2_3616_14100 2.666667e-02
R6771 n2_3616_14100 n2_3616_14241 8.952381e-02
R6772 n2_3616_14241 n2_3616_14274 2.095238e-02
R6773 n2_3616_14274 n2_3616_14457 1.161905e-01
R6774 n2_3616_14457 n2_3616_14490 2.095238e-02
R6775 n2_3616_14490 n2_3616_14536 2.920635e-02
R6776 n2_3616_14536 n2_3616_14673 8.698413e-02
R6777 n2_3616_14673 n2_3616_14706 2.095238e-02
R6778 n2_3616_14706 n2_3616_14889 1.161905e-01
R6779 n2_3616_14889 n2_3616_14922 2.095238e-02
R6780 n2_3616_14922 n2_3616_15049 8.063492e-02
R6781 n2_3616_15138 n2_3616_15145 4.444444e-03
R6782 n2_3616_15145 n2_3616_15321 1.117460e-01
R6783 n2_3616_15321 n2_3616_15354 2.095238e-02
R6784 n2_3616_15354 n2_3616_15368 8.888889e-03
R6785 n2_3616_15368 n2_3616_15537 1.073016e-01
R6786 n2_3616_15537 n2_3616_15570 2.095238e-02
R6787 n2_3616_15570 n2_3616_15584 8.888889e-03
R6788 n2_3616_15584 n2_3616_15753 1.073016e-01
R6789 n2_3616_15753 n2_3616_15786 2.095238e-02
R6790 n2_3616_15786 n2_3616_15969 1.161905e-01
R6791 n2_3616_15969 n2_3616_16002 2.095238e-02
R6792 n2_3616_16002 n2_3616_16185 1.161905e-01
R6793 n2_3616_16185 n2_3616_16218 2.095238e-02
R6794 n2_3616_16218 n2_3616_16401 1.161905e-01
R6795 n2_3616_16401 n2_3616_16434 2.095238e-02
R6796 n2_3616_16434 n2_3616_16471 2.349206e-02
R6797 n2_3616_16471 n2_3616_16617 9.269841e-02
R6798 n2_3616_16617 n2_3616_16650 2.095238e-02
R6799 n2_3616_16650 n2_3616_16664 8.888889e-03
R6800 n2_3616_16664 n2_3616_16833 1.073016e-01
R6801 n2_3616_16833 n2_3616_16866 2.095238e-02
R6802 n2_3616_16866 n2_3616_16880 8.888889e-03
R6803 n2_3616_16880 n2_3616_17049 1.073016e-01
R6804 n2_3616_17049 n2_3616_17082 2.095238e-02
R6805 n2_3616_17082 n2_3616_17265 1.161905e-01
R6806 n2_3616_17265 n2_3616_17298 2.095238e-02
R6807 n2_3616_17298 n2_3616_17299 6.349206e-04
R6808 n2_3616_17395 n2_3616_17481 5.460317e-02
R6809 n2_3616_17481 n2_3616_17514 2.095238e-02
R6810 n2_3616_17514 n2_3616_17528 8.888889e-03
R6811 n2_3616_17528 n2_3616_17551 1.460317e-02
R6812 n2_3616_17551 n2_3616_17697 9.269841e-02
R6813 n2_3616_17697 n2_3616_17730 2.095238e-02
R6814 n2_3616_17730 n2_3616_17913 1.161905e-01
R6815 n2_3616_17913 n2_3616_17946 2.095238e-02
R6816 n2_3616_17946 n2_3616_18129 1.161905e-01
R6817 n2_3616_18129 n2_3616_18162 2.095238e-02
R6818 n2_3616_18162 n2_3616_18345 1.161905e-01
R6819 n2_3616_18345 n2_3616_18378 2.095238e-02
R6820 n2_3616_18378 n2_3616_18424 2.920635e-02
R6821 n2_3616_18520 n2_3616_18561 2.603175e-02
R6822 n2_3616_18561 n2_3616_18594 2.095238e-02
R6823 n2_3616_18594 n2_3616_18777 1.161905e-01
R6824 n2_3616_18777 n2_3616_18810 2.095238e-02
R6825 n2_3616_18810 n2_3616_18993 1.161905e-01
R6826 n2_3616_18993 n2_3616_19026 2.095238e-02
R6827 n2_3616_19026 n2_3616_19209 1.161905e-01
R6828 n2_3616_19209 n2_3616_19242 2.095238e-02
R6829 n2_3616_19242 n2_3616_19425 1.161905e-01
R6830 n2_3616_19425 n2_3616_19458 2.095238e-02
R6831 n2_3616_19458 n2_3616_19549 5.777778e-02
R6832 n2_3616_19641 n2_3616_19645 2.539683e-03
R6833 n2_3616_19645 n2_3616_19674 1.841270e-02
R6834 n2_3616_19674 n2_3616_19857 1.161905e-01
R6835 n2_3616_19857 n2_3616_19890 2.095238e-02
R6836 n2_3616_19890 n2_3616_20073 1.161905e-01
R6837 n2_3616_20073 n2_3616_20106 2.095238e-02
R6838 n2_3616_20106 n2_3616_20289 1.161905e-01
R6839 n2_3616_20289 n2_3616_20322 2.095238e-02
R6840 n2_3616_20322 n2_3616_20505 1.161905e-01
R6841 n2_3616_20505 n2_3616_20538 2.095238e-02
R6842 n2_3616_20538 n2_3616_20674 8.634921e-02
R6843 n2_3616_20754 n2_3616_20770 1.015873e-02
R6844 n2_3616_20770 n2_3616_20937 1.060317e-01
R6845 n2_3616_20937 n2_3616_20970 2.095238e-02
R6846 n2_3616_3895 n2_3708_3895 5.841270e-02
R6847 n2_3708_3895 n2_3755_3895 2.984127e-02
R6848 n2_3755_3895 n2_3804_3895 3.111111e-02
R6849 n2_3616_6049 n2_3755_6049 8.825397e-02
R6850 n2_3755_6049 n2_3804_6049 3.111111e-02
R6851 n2_3616_6145 n2_3755_6145 8.825397e-02
R6852 n2_3755_6145 n2_3804_6145 3.111111e-02
R6853 n2_3616_8299 n2_3755_8299 8.825397e-02
R6854 n2_3755_8299 n2_3804_8299 3.111111e-02
R6855 n2_3616_8395 n2_3755_8395 8.825397e-02
R6856 n2_3755_8395 n2_3804_8395 3.111111e-02
R6857 n2_3616_10549 n2_3755_10549 8.825397e-02
R6858 n2_3755_10549 n2_3804_10549 3.111111e-02
R6859 n2_3616_10645 n2_3755_10645 8.825397e-02
R6860 n2_3755_10645 n2_3804_10645 3.111111e-02
R6861 n2_3616_12799 n2_3755_12799 8.825397e-02
R6862 n2_3755_12799 n2_3804_12799 3.111111e-02
R6863 n2_3616_12895 n2_3755_12895 8.825397e-02
R6864 n2_3755_12895 n2_3804_12895 3.111111e-02
R6865 n2_3616_15049 n2_3755_15049 8.825397e-02
R6866 n2_3755_15049 n2_3804_15049 3.111111e-02
R6867 n2_3616_15145 n2_3755_15145 8.825397e-02
R6868 n2_3755_15145 n2_3804_15145 3.111111e-02
R6869 n2_3616_17299 n2_3708_17299 5.841270e-02
R6870 n2_3708_17299 n2_3755_17299 2.984127e-02
R6871 n2_3755_17299 n2_3804_17299 3.111111e-02
R6872 n2_3616_424 n2_3708_424 5.841270e-02
R6873 n2_3708_424 n2_3755_424 2.984127e-02
R6874 n2_3755_424 n2_3804_424 3.111111e-02
R6875 n2_3804_424 n2_3896_424 5.841270e-02
R6876 n2_3616_520 n2_3708_520 5.841270e-02
R6877 n2_3708_520 n2_3755_520 2.984127e-02
R6878 n2_3755_520 n2_3804_520 3.111111e-02
R6879 n2_3804_520 n2_3896_520 5.841270e-02
R6880 n2_3616_1549 n2_3708_1549 5.841270e-02
R6881 n2_3708_1549 n2_3755_1549 2.984127e-02
R6882 n2_3755_1549 n2_3804_1549 3.111111e-02
R6883 n2_3804_1549 n2_3896_1549 5.841270e-02
R6884 n2_3616_1645 n2_3708_1645 5.841270e-02
R6885 n2_3708_1645 n2_3755_1645 2.984127e-02
R6886 n2_3755_1645 n2_3804_1645 3.111111e-02
R6887 n2_3804_1645 n2_3896_1645 5.841270e-02
R6888 n2_3616_2674 n2_3708_2674 5.841270e-02
R6889 n2_3708_2674 n2_3755_2674 2.984127e-02
R6890 n2_3755_2674 n2_3804_2674 3.111111e-02
R6891 n2_3804_2674 n2_3896_2674 5.841270e-02
R6892 n2_3616_2770 n2_3708_2770 5.841270e-02
R6893 n2_3708_2770 n2_3755_2770 2.984127e-02
R6894 n2_3755_2770 n2_3804_2770 3.111111e-02
R6895 n2_3804_2770 n2_3896_2770 5.841270e-02
R6896 n2_3616_3799 n2_3708_3799 5.841270e-02
R6897 n2_3708_3799 n2_3755_3799 2.984127e-02
R6898 n2_3755_3799 n2_3804_3799 3.111111e-02
R6899 n2_3804_3799 n2_3896_3799 5.841270e-02
R6900 n2_3616_17395 n2_3708_17395 5.841270e-02
R6901 n2_3708_17395 n2_3755_17395 2.984127e-02
R6902 n2_3755_17395 n2_3804_17395 3.111111e-02
R6903 n2_3804_17395 n2_3896_17395 5.841270e-02
R6904 n2_3616_18424 n2_3708_18424 5.841270e-02
R6905 n2_3708_18424 n2_3755_18424 2.984127e-02
R6906 n2_3755_18424 n2_3804_18424 3.111111e-02
R6907 n2_3804_18424 n2_3896_18424 5.841270e-02
R6908 n2_3616_18520 n2_3708_18520 5.841270e-02
R6909 n2_3708_18520 n2_3755_18520 2.984127e-02
R6910 n2_3755_18520 n2_3804_18520 3.111111e-02
R6911 n2_3804_18520 n2_3896_18520 5.841270e-02
R6912 n2_3616_19549 n2_3708_19549 5.841270e-02
R6913 n2_3708_19549 n2_3755_19549 2.984127e-02
R6914 n2_3755_19549 n2_3804_19549 3.111111e-02
R6915 n2_3804_19549 n2_3896_19549 5.841270e-02
R6916 n2_3616_19645 n2_3708_19645 5.841270e-02
R6917 n2_3708_19645 n2_3755_19645 2.984127e-02
R6918 n2_3755_19645 n2_3804_19645 3.111111e-02
R6919 n2_3804_19645 n2_3896_19645 5.841270e-02
R6920 n2_3616_20674 n2_3708_20674 5.841270e-02
R6921 n2_3708_20674 n2_3755_20674 2.984127e-02
R6922 n2_3755_20674 n2_3804_20674 3.111111e-02
R6923 n2_3804_20674 n2_3896_20674 5.841270e-02
R6924 n2_3616_20770 n2_3708_20770 5.841270e-02
R6925 n2_3708_20770 n2_3755_20770 2.984127e-02
R6926 n2_3755_20770 n2_3804_20770 3.111111e-02
R6927 n2_3804_20770 n2_3896_20770 5.841270e-02
R6928 n2_3708_201 n2_3708_234 2.095238e-02
R6929 n2_3708_234 n2_3708_356 7.746032e-02
R6930 n2_3708_356 n2_3708_417 3.873016e-02
R6931 n2_3708_417 n2_3708_424 4.444444e-03
R6932 n2_3708_424 n2_3708_450 1.650794e-02
R6933 n2_3708_450 n2_3708_520 4.444444e-02
R6934 n2_3708_520 n2_3708_633 7.174603e-02
R6935 n2_3708_633 n2_3708_666 2.095238e-02
R6936 n2_3708_666 n2_3708_788 7.746032e-02
R6937 n2_3708_788 n2_3708_849 3.873016e-02
R6938 n2_3708_849 n2_3708_882 2.095238e-02
R6939 n2_3708_882 n2_3708_1065 1.161905e-01
R6940 n2_3708_1065 n2_3708_1098 2.095238e-02
R6941 n2_3708_1098 n2_3708_1281 1.161905e-01
R6942 n2_3708_1281 n2_3708_1314 2.095238e-02
R6943 n2_3708_1314 n2_3708_1497 1.161905e-01
R6944 n2_3708_1497 n2_3708_1530 2.095238e-02
R6945 n2_3708_1530 n2_3708_1549 1.206349e-02
R6946 n2_3708_1549 n2_3708_1645 6.095238e-02
R6947 n2_3708_1645 n2_3708_1652 4.444444e-03
R6948 n2_3708_1652 n2_3708_1713 3.873016e-02
R6949 n2_3708_1713 n2_3708_1746 2.095238e-02
R6950 n2_3708_1746 n2_3708_1929 1.161905e-01
R6951 n2_3708_1929 n2_3708_1962 2.095238e-02
R6952 n2_3708_1962 n2_3708_1976 8.888889e-03
R6953 n2_3708_1976 n2_3708_2145 1.073016e-01
R6954 n2_3708_2145 n2_3708_2178 2.095238e-02
R6955 n2_3708_2178 n2_3708_2361 1.161905e-01
R6956 n2_3708_2361 n2_3708_2394 2.095238e-02
R6957 n2_3708_2394 n2_3708_2577 1.161905e-01
R6958 n2_3708_2577 n2_3708_2610 2.095238e-02
R6959 n2_3708_2610 n2_3708_2674 4.063492e-02
R6960 n2_3708_2674 n2_3708_2770 6.095238e-02
R6961 n2_3708_2770 n2_3708_2793 1.460317e-02
R6962 n2_3708_2793 n2_3708_2826 2.095238e-02
R6963 n2_3708_2826 n2_3708_3009 1.161905e-01
R6964 n2_3708_3009 n2_3708_3042 2.095238e-02
R6965 n2_3708_3042 n2_3708_3225 1.161905e-01
R6966 n2_3708_3225 n2_3708_3258 2.095238e-02
R6967 n2_3708_3258 n2_3708_3441 1.161905e-01
R6968 n2_3708_3441 n2_3708_3474 2.095238e-02
R6969 n2_3708_3474 n2_3708_3657 1.161905e-01
R6970 n2_3708_3657 n2_3708_3690 2.095238e-02
R6971 n2_3708_3690 n2_3708_3704 8.888889e-03
R6972 n2_3708_3704 n2_3708_3799 6.031746e-02
R6973 n2_3708_3799 n2_3708_3873 4.698413e-02
R6974 n2_3708_3873 n2_3708_3895 1.396825e-02
R6975 n2_3708_3895 n2_3708_3906 6.984127e-03
R6976 n2_3708_3906 n2_3708_3920 8.888889e-03
R6977 n2_3708_17265 n2_3708_17298 2.095238e-02
R6978 n2_3708_17298 n2_3708_17299 6.349206e-04
R6979 n2_3708_17299 n2_3708_17335 2.285714e-02
R6980 n2_3708_17335 n2_3708_17395 3.809524e-02
R6981 n2_3708_17395 n2_3708_17481 5.460317e-02
R6982 n2_3708_17481 n2_3708_17514 2.095238e-02
R6983 n2_3708_17514 n2_3708_17528 8.888889e-03
R6984 n2_3708_17528 n2_3708_17551 1.460317e-02
R6985 n2_3708_17551 n2_3708_17697 9.269841e-02
R6986 n2_3708_17697 n2_3708_17730 2.095238e-02
R6987 n2_3708_17730 n2_3708_17913 1.161905e-01
R6988 n2_3708_17913 n2_3708_17946 2.095238e-02
R6989 n2_3708_17946 n2_3708_18129 1.161905e-01
R6990 n2_3708_18129 n2_3708_18162 2.095238e-02
R6991 n2_3708_18162 n2_3708_18345 1.161905e-01
R6992 n2_3708_18345 n2_3708_18378 2.095238e-02
R6993 n2_3708_18378 n2_3708_18424 2.920635e-02
R6994 n2_3708_18424 n2_3708_18520 6.095238e-02
R6995 n2_3708_18520 n2_3708_18561 2.603175e-02
R6996 n2_3708_18561 n2_3708_18594 2.095238e-02
R6997 n2_3708_18594 n2_3708_18777 1.161905e-01
R6998 n2_3708_18777 n2_3708_18810 2.095238e-02
R6999 n2_3708_18810 n2_3708_18993 1.161905e-01
R7000 n2_3708_18993 n2_3708_19026 2.095238e-02
R7001 n2_3708_19026 n2_3708_19209 1.161905e-01
R7002 n2_3708_19209 n2_3708_19242 2.095238e-02
R7003 n2_3708_19242 n2_3708_19425 1.161905e-01
R7004 n2_3708_19425 n2_3708_19458 2.095238e-02
R7005 n2_3708_19458 n2_3708_19549 5.777778e-02
R7006 n2_3708_19549 n2_3708_19641 5.841270e-02
R7007 n2_3708_19641 n2_3708_19645 2.539683e-03
R7008 n2_3708_19645 n2_3708_19674 1.841270e-02
R7009 n2_3708_19674 n2_3708_19857 1.161905e-01
R7010 n2_3708_19857 n2_3708_19890 2.095238e-02
R7011 n2_3708_19890 n2_3708_20073 1.161905e-01
R7012 n2_3708_20073 n2_3708_20106 2.095238e-02
R7013 n2_3708_20106 n2_3708_20289 1.161905e-01
R7014 n2_3708_20289 n2_3708_20322 2.095238e-02
R7015 n2_3708_20322 n2_3708_20505 1.161905e-01
R7016 n2_3708_20505 n2_3708_20538 2.095238e-02
R7017 n2_3708_20538 n2_3708_20674 8.634921e-02
R7018 n2_3708_20674 n2_3708_20721 2.984127e-02
R7019 n2_3708_20721 n2_3708_20754 2.095238e-02
R7020 n2_3708_20754 n2_3708_20770 1.015873e-02
R7021 n2_3708_20770 n2_3708_20937 1.060317e-01
R7022 n2_3708_20937 n2_3708_20970 2.095238e-02
R7023 n2_3804_201 n2_3804_234 2.095238e-02
R7024 n2_3804_234 n2_3804_356 7.746032e-02
R7025 n2_3804_356 n2_3804_417 3.873016e-02
R7026 n2_3804_417 n2_3804_424 4.444444e-03
R7027 n2_3804_424 n2_3804_450 1.650794e-02
R7028 n2_3804_450 n2_3804_520 4.444444e-02
R7029 n2_3804_520 n2_3804_633 7.174603e-02
R7030 n2_3804_633 n2_3804_666 2.095238e-02
R7031 n2_3804_666 n2_3804_788 7.746032e-02
R7032 n2_3804_788 n2_3804_849 3.873016e-02
R7033 n2_3804_849 n2_3804_882 2.095238e-02
R7034 n2_3804_882 n2_3804_1065 1.161905e-01
R7035 n2_3804_1065 n2_3804_1098 2.095238e-02
R7036 n2_3804_1098 n2_3804_1281 1.161905e-01
R7037 n2_3804_1281 n2_3804_1314 2.095238e-02
R7038 n2_3804_1314 n2_3804_1497 1.161905e-01
R7039 n2_3804_1497 n2_3804_1530 2.095238e-02
R7040 n2_3804_1530 n2_3804_1549 1.206349e-02
R7041 n2_3804_1549 n2_3804_1645 6.095238e-02
R7042 n2_3804_1645 n2_3804_1652 4.444444e-03
R7043 n2_3804_1652 n2_3804_1713 3.873016e-02
R7044 n2_3804_1713 n2_3804_1746 2.095238e-02
R7045 n2_3804_1746 n2_3804_1929 1.161905e-01
R7046 n2_3804_1929 n2_3804_1962 2.095238e-02
R7047 n2_3804_1962 n2_3804_1976 8.888889e-03
R7048 n2_3804_1976 n2_3804_2145 1.073016e-01
R7049 n2_3804_2145 n2_3804_2178 2.095238e-02
R7050 n2_3804_2178 n2_3804_2361 1.161905e-01
R7051 n2_3804_2361 n2_3804_2394 2.095238e-02
R7052 n2_3804_2394 n2_3804_2577 1.161905e-01
R7053 n2_3804_2577 n2_3804_2610 2.095238e-02
R7054 n2_3804_2610 n2_3804_2674 4.063492e-02
R7055 n2_3804_2674 n2_3804_2770 6.095238e-02
R7056 n2_3804_2770 n2_3804_2793 1.460317e-02
R7057 n2_3804_2793 n2_3804_2826 2.095238e-02
R7058 n2_3804_2826 n2_3804_3009 1.161905e-01
R7059 n2_3804_3009 n2_3804_3042 2.095238e-02
R7060 n2_3804_3042 n2_3804_3225 1.161905e-01
R7061 n2_3804_3225 n2_3804_3258 2.095238e-02
R7062 n2_3804_3258 n2_3804_3441 1.161905e-01
R7063 n2_3804_3441 n2_3804_3474 2.095238e-02
R7064 n2_3804_3474 n2_3804_3657 1.161905e-01
R7065 n2_3804_3657 n2_3804_3690 2.095238e-02
R7066 n2_3804_3690 n2_3804_3704 8.888889e-03
R7067 n2_3804_3704 n2_3804_3799 6.031746e-02
R7068 n2_3804_3799 n2_3804_3873 4.698413e-02
R7069 n2_3804_3873 n2_3804_3895 1.396825e-02
R7070 n2_3804_3895 n2_3804_3906 6.984127e-03
R7071 n2_3804_3906 n2_3804_3920 8.888889e-03
R7072 n2_3804_3920 n2_3804_4089 1.073016e-01
R7073 n2_3804_4089 n2_3804_4122 2.095238e-02
R7074 n2_3804_4122 n2_3804_4136 8.888889e-03
R7075 n2_3804_4136 n2_3804_4159 1.460317e-02
R7076 n2_3804_4159 n2_3804_4305 9.269841e-02
R7077 n2_3804_4305 n2_3804_4338 2.095238e-02
R7078 n2_3804_4338 n2_3804_4352 8.888889e-03
R7079 n2_3804_4352 n2_3804_4375 1.460317e-02
R7080 n2_3804_4375 n2_3804_4521 9.269841e-02
R7081 n2_3804_4521 n2_3804_4554 2.095238e-02
R7082 n2_3804_4554 n2_3804_4737 1.161905e-01
R7083 n2_3804_4737 n2_3804_4770 2.095238e-02
R7084 n2_3804_5169 n2_3804_5202 2.095238e-02
R7085 n2_3804_5202 n2_3804_5385 1.161905e-01
R7086 n2_3804_5385 n2_3804_5418 2.095238e-02
R7087 n2_3804_5418 n2_3804_5432 8.888889e-03
R7088 n2_3804_5432 n2_3804_5601 1.073016e-01
R7089 n2_3804_5601 n2_3804_5634 2.095238e-02
R7090 n2_3804_5634 n2_3804_5817 1.161905e-01
R7091 n2_3804_5817 n2_3804_5850 2.095238e-02
R7092 n2_3804_5850 n2_3804_6033 1.161905e-01
R7093 n2_3804_6033 n2_3804_6049 1.015873e-02
R7094 n2_3804_6049 n2_3804_6066 1.079365e-02
R7095 n2_3804_6066 n2_3804_6145 5.015873e-02
R7096 n2_3804_6145 n2_3804_6249 6.603175e-02
R7097 n2_3804_6249 n2_3804_6282 2.095238e-02
R7098 n2_3804_6282 n2_3804_6465 1.161905e-01
R7099 n2_3804_6465 n2_3804_6498 2.095238e-02
R7100 n2_3804_6498 n2_3804_6535 2.349206e-02
R7101 n2_3804_6535 n2_3804_6681 9.269841e-02
R7102 n2_3804_6681 n2_3804_6714 2.095238e-02
R7103 n2_3804_6714 n2_3804_6897 1.161905e-01
R7104 n2_3804_6897 n2_3804_6930 2.095238e-02
R7105 n2_3804_6930 n2_3804_7113 1.161905e-01
R7106 n2_3804_7329 n2_3804_7362 2.095238e-02
R7107 n2_3804_7362 n2_3804_7545 1.161905e-01
R7108 n2_3804_7545 n2_3804_7578 2.095238e-02
R7109 n2_3804_7578 n2_3804_7761 1.161905e-01
R7110 n2_3804_7761 n2_3804_7794 2.095238e-02
R7111 n2_3804_7794 n2_3804_7808 8.888889e-03
R7112 n2_3804_7808 n2_3804_7977 1.073016e-01
R7113 n2_3804_7977 n2_3804_8010 2.095238e-02
R7114 n2_3804_8010 n2_3804_8193 1.161905e-01
R7115 n2_3804_8193 n2_3804_8226 2.095238e-02
R7116 n2_3804_8226 n2_3804_8299 4.634921e-02
R7117 n2_3804_8299 n2_3804_8395 6.095238e-02
R7118 n2_3804_8395 n2_3804_8409 8.888889e-03
R7119 n2_3804_8409 n2_3804_8442 2.095238e-02
R7120 n2_3804_8442 n2_3804_8625 1.161905e-01
R7121 n2_3804_8625 n2_3804_8658 2.095238e-02
R7122 n2_3804_8658 n2_3804_8841 1.161905e-01
R7123 n2_3804_8841 n2_3804_8874 2.095238e-02
R7124 n2_3804_8874 n2_3804_8888 8.888889e-03
R7125 n2_3804_8888 n2_3804_8911 1.460317e-02
R7126 n2_3804_8911 n2_3804_9057 9.269841e-02
R7127 n2_3804_9057 n2_3804_9090 2.095238e-02
R7128 n2_3804_9090 n2_3804_9273 1.161905e-01
R7129 n2_3804_9273 n2_3804_9306 2.095238e-02
R7130 n2_3804_9705 n2_3804_9738 2.095238e-02
R7131 n2_3804_9738 n2_3804_9921 1.161905e-01
R7132 n2_3804_9921 n2_3804_9954 2.095238e-02
R7133 n2_3804_9954 n2_3804_9968 8.888889e-03
R7134 n2_3804_9968 n2_3804_10137 1.073016e-01
R7135 n2_3804_10137 n2_3804_10170 2.095238e-02
R7136 n2_3804_10170 n2_3804_10353 1.161905e-01
R7137 n2_3804_10353 n2_3804_10386 2.095238e-02
R7138 n2_3804_10386 n2_3804_10549 1.034921e-01
R7139 n2_3804_10549 n2_3804_10569 1.269841e-02
R7140 n2_3804_10569 n2_3804_10602 2.095238e-02
R7141 n2_3804_10602 n2_3804_10645 2.730159e-02
R7142 n2_3804_10645 n2_3804_10785 8.888889e-02
R7143 n2_3804_10785 n2_3804_10818 2.095238e-02
R7144 n2_3804_10818 n2_3804_11001 1.161905e-01
R7145 n2_3804_11001 n2_3804_11034 2.095238e-02
R7146 n2_3804_11034 n2_3804_11048 8.888889e-03
R7147 n2_3804_11048 n2_3804_11217 1.073016e-01
R7148 n2_3804_11217 n2_3804_11250 2.095238e-02
R7149 n2_3804_11250 n2_3804_11433 1.161905e-01
R7150 n2_3804_11433 n2_3804_11466 2.095238e-02
R7151 n2_3804_11865 n2_3804_11898 2.095238e-02
R7152 n2_3804_11898 n2_3804_12081 1.161905e-01
R7153 n2_3804_12081 n2_3804_12114 2.095238e-02
R7154 n2_3804_12114 n2_3804_12128 8.888889e-03
R7155 n2_3804_12128 n2_3804_12151 1.460317e-02
R7156 n2_3804_12151 n2_3804_12297 9.269841e-02
R7157 n2_3804_12297 n2_3804_12330 2.095238e-02
R7158 n2_3804_12330 n2_3804_12513 1.161905e-01
R7159 n2_3804_12513 n2_3804_12546 2.095238e-02
R7160 n2_3804_12546 n2_3804_12729 1.161905e-01
R7161 n2_3804_12729 n2_3804_12762 2.095238e-02
R7162 n2_3804_12762 n2_3804_12799 2.349206e-02
R7163 n2_3804_12799 n2_3804_12895 6.095238e-02
R7164 n2_3804_12895 n2_3804_12945 3.174603e-02
R7165 n2_3804_12945 n2_3804_12978 2.095238e-02
R7166 n2_3804_12978 n2_3804_13161 1.161905e-01
R7167 n2_3804_13161 n2_3804_13194 2.095238e-02
R7168 n2_3804_13194 n2_3804_13377 1.161905e-01
R7169 n2_3804_13377 n2_3804_13410 2.095238e-02
R7170 n2_3804_13410 n2_3804_13424 8.888889e-03
R7171 n2_3804_13424 n2_3804_13593 1.073016e-01
R7172 n2_3804_13593 n2_3804_13626 2.095238e-02
R7173 n2_3804_13626 n2_3804_13640 8.888889e-03
R7174 n2_3804_13640 n2_3804_13809 1.073016e-01
R7175 n2_3804_13809 n2_3804_13842 2.095238e-02
R7176 n2_3804_14100 n2_3804_14241 8.952381e-02
R7177 n2_3804_14241 n2_3804_14274 2.095238e-02
R7178 n2_3804_14274 n2_3804_14457 1.161905e-01
R7179 n2_3804_14457 n2_3804_14490 2.095238e-02
R7180 n2_3804_14490 n2_3804_14536 2.920635e-02
R7181 n2_3804_14536 n2_3804_14673 8.698413e-02
R7182 n2_3804_14673 n2_3804_14706 2.095238e-02
R7183 n2_3804_14706 n2_3804_14889 1.161905e-01
R7184 n2_3804_14889 n2_3804_14922 2.095238e-02
R7185 n2_3804_14922 n2_3804_15049 8.063492e-02
R7186 n2_3804_15049 n2_3804_15105 3.555556e-02
R7187 n2_3804_15105 n2_3804_15138 2.095238e-02
R7188 n2_3804_15138 n2_3804_15145 4.444444e-03
R7189 n2_3804_15145 n2_3804_15321 1.117460e-01
R7190 n2_3804_15321 n2_3804_15354 2.095238e-02
R7191 n2_3804_15354 n2_3804_15368 8.888889e-03
R7192 n2_3804_15368 n2_3804_15537 1.073016e-01
R7193 n2_3804_15537 n2_3804_15570 2.095238e-02
R7194 n2_3804_15570 n2_3804_15584 8.888889e-03
R7195 n2_3804_15584 n2_3804_15753 1.073016e-01
R7196 n2_3804_15753 n2_3804_15786 2.095238e-02
R7197 n2_3804_15786 n2_3804_15969 1.161905e-01
R7198 n2_3804_15969 n2_3804_16002 2.095238e-02
R7199 n2_3804_16401 n2_3804_16434 2.095238e-02
R7200 n2_3804_16434 n2_3804_16471 2.349206e-02
R7201 n2_3804_16471 n2_3804_16617 9.269841e-02
R7202 n2_3804_16617 n2_3804_16650 2.095238e-02
R7203 n2_3804_16650 n2_3804_16664 8.888889e-03
R7204 n2_3804_16664 n2_3804_16833 1.073016e-01
R7205 n2_3804_16833 n2_3804_16866 2.095238e-02
R7206 n2_3804_16866 n2_3804_16880 8.888889e-03
R7207 n2_3804_16880 n2_3804_17049 1.073016e-01
R7208 n2_3804_17049 n2_3804_17082 2.095238e-02
R7209 n2_3804_17082 n2_3804_17265 1.161905e-01
R7210 n2_3804_17265 n2_3804_17298 2.095238e-02
R7211 n2_3804_17298 n2_3804_17299 6.349206e-04
R7212 n2_3804_17299 n2_3804_17335 2.285714e-02
R7213 n2_3804_17335 n2_3804_17395 3.809524e-02
R7214 n2_3804_17395 n2_3804_17481 5.460317e-02
R7215 n2_3804_17481 n2_3804_17514 2.095238e-02
R7216 n2_3804_17514 n2_3804_17528 8.888889e-03
R7217 n2_3804_17528 n2_3804_17551 1.460317e-02
R7218 n2_3804_17551 n2_3804_17697 9.269841e-02
R7219 n2_3804_17697 n2_3804_17730 2.095238e-02
R7220 n2_3804_17730 n2_3804_17913 1.161905e-01
R7221 n2_3804_17913 n2_3804_17946 2.095238e-02
R7222 n2_3804_17946 n2_3804_18129 1.161905e-01
R7223 n2_3804_18129 n2_3804_18162 2.095238e-02
R7224 n2_3804_18162 n2_3804_18345 1.161905e-01
R7225 n2_3804_18345 n2_3804_18378 2.095238e-02
R7226 n2_3804_18378 n2_3804_18424 2.920635e-02
R7227 n2_3804_18424 n2_3804_18520 6.095238e-02
R7228 n2_3804_18520 n2_3804_18561 2.603175e-02
R7229 n2_3804_18561 n2_3804_18594 2.095238e-02
R7230 n2_3804_18594 n2_3804_18777 1.161905e-01
R7231 n2_3804_18777 n2_3804_18810 2.095238e-02
R7232 n2_3804_18810 n2_3804_18993 1.161905e-01
R7233 n2_3804_18993 n2_3804_19026 2.095238e-02
R7234 n2_3804_19026 n2_3804_19209 1.161905e-01
R7235 n2_3804_19209 n2_3804_19242 2.095238e-02
R7236 n2_3804_19242 n2_3804_19425 1.161905e-01
R7237 n2_3804_19425 n2_3804_19458 2.095238e-02
R7238 n2_3804_19458 n2_3804_19549 5.777778e-02
R7239 n2_3804_19549 n2_3804_19641 5.841270e-02
R7240 n2_3804_19641 n2_3804_19645 2.539683e-03
R7241 n2_3804_19645 n2_3804_19674 1.841270e-02
R7242 n2_3804_19674 n2_3804_19857 1.161905e-01
R7243 n2_3804_19857 n2_3804_19890 2.095238e-02
R7244 n2_3804_19890 n2_3804_20073 1.161905e-01
R7245 n2_3804_20073 n2_3804_20106 2.095238e-02
R7246 n2_3804_20106 n2_3804_20289 1.161905e-01
R7247 n2_3804_20289 n2_3804_20322 2.095238e-02
R7248 n2_3804_20322 n2_3804_20505 1.161905e-01
R7249 n2_3804_20505 n2_3804_20538 2.095238e-02
R7250 n2_3804_20538 n2_3804_20674 8.634921e-02
R7251 n2_3804_20674 n2_3804_20721 2.984127e-02
R7252 n2_3804_20721 n2_3804_20754 2.095238e-02
R7253 n2_3804_20754 n2_3804_20770 1.015873e-02
R7254 n2_3804_20770 n2_3804_20937 1.060317e-01
R7255 n2_3804_20937 n2_3804_20970 2.095238e-02
R7256 n2_3896_201 n2_3896_234 2.095238e-02
R7257 n2_3896_234 n2_3896_356 7.746032e-02
R7258 n2_3896_356 n2_3896_417 3.873016e-02
R7259 n2_3896_417 n2_3896_424 4.444444e-03
R7260 n2_3896_424 n2_3896_450 1.650794e-02
R7261 n2_3896_520 n2_3896_633 7.174603e-02
R7262 n2_3896_633 n2_3896_666 2.095238e-02
R7263 n2_3896_666 n2_3896_788 7.746032e-02
R7264 n2_3896_788 n2_3896_849 3.873016e-02
R7265 n2_3896_849 n2_3896_882 2.095238e-02
R7266 n2_3896_882 n2_3896_1065 1.161905e-01
R7267 n2_3896_1065 n2_3896_1098 2.095238e-02
R7268 n2_3896_1098 n2_3896_1281 1.161905e-01
R7269 n2_3896_1281 n2_3896_1314 2.095238e-02
R7270 n2_3896_1314 n2_3896_1497 1.161905e-01
R7271 n2_3896_1497 n2_3896_1530 2.095238e-02
R7272 n2_3896_1530 n2_3896_1549 1.206349e-02
R7273 n2_3896_1645 n2_3896_1652 4.444444e-03
R7274 n2_3896_1652 n2_3896_1713 3.873016e-02
R7275 n2_3896_1713 n2_3896_1746 2.095238e-02
R7276 n2_3896_1746 n2_3896_1929 1.161905e-01
R7277 n2_3896_1929 n2_3896_1962 2.095238e-02
R7278 n2_3896_1962 n2_3896_1976 8.888889e-03
R7279 n2_3896_1976 n2_3896_2145 1.073016e-01
R7280 n2_3896_2145 n2_3896_2178 2.095238e-02
R7281 n2_3896_2178 n2_3896_2361 1.161905e-01
R7282 n2_3896_2361 n2_3896_2394 2.095238e-02
R7283 n2_3896_2394 n2_3896_2577 1.161905e-01
R7284 n2_3896_2577 n2_3896_2610 2.095238e-02
R7285 n2_3896_2610 n2_3896_2674 4.063492e-02
R7286 n2_3896_2770 n2_3896_2793 1.460317e-02
R7287 n2_3896_2793 n2_3896_2826 2.095238e-02
R7288 n2_3896_2826 n2_3896_3009 1.161905e-01
R7289 n2_3896_3009 n2_3896_3042 2.095238e-02
R7290 n2_3896_3042 n2_3896_3225 1.161905e-01
R7291 n2_3896_3225 n2_3896_3258 2.095238e-02
R7292 n2_3896_3258 n2_3896_3441 1.161905e-01
R7293 n2_3896_3441 n2_3896_3474 2.095238e-02
R7294 n2_3896_3474 n2_3896_3657 1.161905e-01
R7295 n2_3896_3657 n2_3896_3690 2.095238e-02
R7296 n2_3896_3690 n2_3896_3704 8.888889e-03
R7297 n2_3896_3704 n2_3896_3799 6.031746e-02
R7298 n2_3896_17395 n2_3896_17481 5.460317e-02
R7299 n2_3896_17481 n2_3896_17514 2.095238e-02
R7300 n2_3896_17514 n2_3896_17528 8.888889e-03
R7301 n2_3896_17528 n2_3896_17551 1.460317e-02
R7302 n2_3896_17551 n2_3896_17697 9.269841e-02
R7303 n2_3896_17697 n2_3896_17730 2.095238e-02
R7304 n2_3896_17730 n2_3896_17913 1.161905e-01
R7305 n2_3896_17913 n2_3896_17946 2.095238e-02
R7306 n2_3896_17946 n2_3896_18129 1.161905e-01
R7307 n2_3896_18129 n2_3896_18162 2.095238e-02
R7308 n2_3896_18162 n2_3896_18345 1.161905e-01
R7309 n2_3896_18345 n2_3896_18378 2.095238e-02
R7310 n2_3896_18378 n2_3896_18424 2.920635e-02
R7311 n2_3896_18520 n2_3896_18561 2.603175e-02
R7312 n2_3896_18561 n2_3896_18594 2.095238e-02
R7313 n2_3896_18594 n2_3896_18777 1.161905e-01
R7314 n2_3896_18777 n2_3896_18810 2.095238e-02
R7315 n2_3896_18810 n2_3896_18993 1.161905e-01
R7316 n2_3896_18993 n2_3896_19026 2.095238e-02
R7317 n2_3896_19026 n2_3896_19209 1.161905e-01
R7318 n2_3896_19209 n2_3896_19242 2.095238e-02
R7319 n2_3896_19242 n2_3896_19425 1.161905e-01
R7320 n2_3896_19425 n2_3896_19458 2.095238e-02
R7321 n2_3896_19458 n2_3896_19549 5.777778e-02
R7322 n2_3896_19641 n2_3896_19645 2.539683e-03
R7323 n2_3896_19645 n2_3896_19674 1.841270e-02
R7324 n2_3896_19674 n2_3896_19857 1.161905e-01
R7325 n2_3896_19857 n2_3896_19890 2.095238e-02
R7326 n2_3896_19890 n2_3896_20073 1.161905e-01
R7327 n2_3896_20073 n2_3896_20106 2.095238e-02
R7328 n2_3896_20106 n2_3896_20289 1.161905e-01
R7329 n2_3896_20289 n2_3896_20322 2.095238e-02
R7330 n2_3896_20322 n2_3896_20505 1.161905e-01
R7331 n2_3896_20505 n2_3896_20538 2.095238e-02
R7332 n2_3896_20538 n2_3896_20674 8.634921e-02
R7333 n2_3896_20754 n2_3896_20770 1.015873e-02
R7334 n2_3896_20770 n2_3896_20937 1.060317e-01
R7335 n2_3896_20937 n2_3896_20970 2.095238e-02
R7336 n2_4741_5169 n2_4741_5202 2.095238e-02
R7337 n2_4741_5202 n2_4741_5385 1.161905e-01
R7338 n2_4741_5385 n2_4741_5418 2.095238e-02
R7339 n2_4741_5418 n2_4741_5432 8.888889e-03
R7340 n2_4741_5432 n2_4741_5601 1.073016e-01
R7341 n2_4741_5601 n2_4741_5634 2.095238e-02
R7342 n2_4741_5634 n2_4741_5817 1.161905e-01
R7343 n2_4741_5817 n2_4741_5850 2.095238e-02
R7344 n2_4741_5850 n2_4741_6033 1.161905e-01
R7345 n2_4741_6033 n2_4741_6049 1.015873e-02
R7346 n2_4741_6049 n2_4741_6066 1.079365e-02
R7347 n2_4741_6145 n2_4741_6249 6.603175e-02
R7348 n2_4741_6249 n2_4741_6282 2.095238e-02
R7349 n2_4741_6282 n2_4741_6465 1.161905e-01
R7350 n2_4741_6465 n2_4741_6498 2.095238e-02
R7351 n2_4741_6498 n2_4741_6535 2.349206e-02
R7352 n2_4741_6535 n2_4741_6681 9.269841e-02
R7353 n2_4741_6681 n2_4741_6714 2.095238e-02
R7354 n2_4741_6714 n2_4741_6897 1.161905e-01
R7355 n2_4741_6897 n2_4741_6930 2.095238e-02
R7356 n2_4741_6930 n2_4741_7113 1.161905e-01
R7357 n2_4741_7113 n2_4741_7146 2.095238e-02
R7358 n2_4741_7146 n2_4741_7329 1.161905e-01
R7359 n2_4741_7329 n2_4741_7362 2.095238e-02
R7360 n2_4741_7362 n2_4741_7545 1.161905e-01
R7361 n2_4741_7545 n2_4741_7578 2.095238e-02
R7362 n2_4741_7578 n2_4741_7761 1.161905e-01
R7363 n2_4741_7761 n2_4741_7794 2.095238e-02
R7364 n2_4741_7794 n2_4741_7808 8.888889e-03
R7365 n2_4741_7808 n2_4741_7977 1.073016e-01
R7366 n2_4741_7977 n2_4741_8010 2.095238e-02
R7367 n2_4741_8010 n2_4741_8193 1.161905e-01
R7368 n2_4741_8193 n2_4741_8226 2.095238e-02
R7369 n2_4741_8226 n2_4741_8299 4.634921e-02
R7370 n2_4741_8395 n2_4741_8409 8.888889e-03
R7371 n2_4741_8409 n2_4741_8442 2.095238e-02
R7372 n2_4741_8442 n2_4741_8625 1.161905e-01
R7373 n2_4741_8625 n2_4741_8658 2.095238e-02
R7374 n2_4741_8658 n2_4741_8841 1.161905e-01
R7375 n2_4741_8841 n2_4741_8874 2.095238e-02
R7376 n2_4741_8874 n2_4741_8888 8.888889e-03
R7377 n2_4741_8888 n2_4741_8911 1.460317e-02
R7378 n2_4741_8911 n2_4741_9057 9.269841e-02
R7379 n2_4741_9057 n2_4741_9090 2.095238e-02
R7380 n2_4741_9090 n2_4741_9273 1.161905e-01
R7381 n2_4741_9273 n2_4741_9306 2.095238e-02
R7382 n2_4741_9306 n2_4741_9489 1.161905e-01
R7383 n2_4741_9489 n2_4741_9522 2.095238e-02
R7384 n2_4741_9522 n2_4741_9705 1.161905e-01
R7385 n2_4741_9705 n2_4741_9738 2.095238e-02
R7386 n2_4741_9738 n2_4741_9921 1.161905e-01
R7387 n2_4741_9921 n2_4741_9954 2.095238e-02
R7388 n2_4741_9954 n2_4741_9968 8.888889e-03
R7389 n2_4741_9968 n2_4741_10137 1.073016e-01
R7390 n2_4741_10137 n2_4741_10170 2.095238e-02
R7391 n2_4741_10170 n2_4741_10353 1.161905e-01
R7392 n2_4741_10353 n2_4741_10386 2.095238e-02
R7393 n2_4741_10386 n2_4741_10549 1.034921e-01
R7394 n2_4741_10549 n2_4741_10569 1.269841e-02
R7395 n2_4741_10645 n2_4741_10785 8.888889e-02
R7396 n2_4741_10785 n2_4741_10818 2.095238e-02
R7397 n2_4741_10818 n2_4741_11001 1.161905e-01
R7398 n2_4741_11001 n2_4741_11034 2.095238e-02
R7399 n2_4741_11034 n2_4741_11048 8.888889e-03
R7400 n2_4741_11048 n2_4741_11071 1.460317e-02
R7401 n2_4741_11071 n2_4741_11217 9.269841e-02
R7402 n2_4741_11217 n2_4741_11250 2.095238e-02
R7403 n2_4741_11250 n2_4741_11433 1.161905e-01
R7404 n2_4741_11433 n2_4741_11466 2.095238e-02
R7405 n2_4741_11466 n2_4741_11649 1.161905e-01
R7406 n2_4741_11649 n2_4741_11682 2.095238e-02
R7407 n2_4741_11682 n2_4741_11865 1.161905e-01
R7408 n2_4741_11865 n2_4741_11898 2.095238e-02
R7409 n2_4741_11898 n2_4741_12081 1.161905e-01
R7410 n2_4741_12081 n2_4741_12114 2.095238e-02
R7411 n2_4741_12114 n2_4741_12128 8.888889e-03
R7412 n2_4741_12128 n2_4741_12297 1.073016e-01
R7413 n2_4741_12297 n2_4741_12330 2.095238e-02
R7414 n2_4741_12330 n2_4741_12513 1.161905e-01
R7415 n2_4741_12513 n2_4741_12546 2.095238e-02
R7416 n2_4741_12546 n2_4741_12729 1.161905e-01
R7417 n2_4741_12729 n2_4741_12762 2.095238e-02
R7418 n2_4741_12762 n2_4741_12799 2.349206e-02
R7419 n2_4741_12895 n2_4741_12945 3.174603e-02
R7420 n2_4741_12945 n2_4741_12978 2.095238e-02
R7421 n2_4741_12978 n2_4741_13161 1.161905e-01
R7422 n2_4741_13161 n2_4741_13194 2.095238e-02
R7423 n2_4741_13194 n2_4741_13377 1.161905e-01
R7424 n2_4741_13377 n2_4741_13410 2.095238e-02
R7425 n2_4741_13410 n2_4741_13424 8.888889e-03
R7426 n2_4741_13424 n2_4741_13593 1.073016e-01
R7427 n2_4741_13593 n2_4741_13626 2.095238e-02
R7428 n2_4741_13626 n2_4741_13809 1.161905e-01
R7429 n2_4741_13809 n2_4741_13842 2.095238e-02
R7430 n2_4741_13842 n2_4741_13879 2.349206e-02
R7431 n2_4741_13879 n2_4741_14025 9.269841e-02
R7432 n2_4741_14025 n2_4741_14058 2.095238e-02
R7433 n2_4741_14058 n2_4741_14100 2.666667e-02
R7434 n2_4741_14100 n2_4741_14241 8.952381e-02
R7435 n2_4741_14241 n2_4741_14274 2.095238e-02
R7436 n2_4741_14274 n2_4741_14457 1.161905e-01
R7437 n2_4741_14457 n2_4741_14490 2.095238e-02
R7438 n2_4741_14490 n2_4741_14536 2.920635e-02
R7439 n2_4741_14536 n2_4741_14673 8.698413e-02
R7440 n2_4741_14673 n2_4741_14706 2.095238e-02
R7441 n2_4741_14706 n2_4741_14889 1.161905e-01
R7442 n2_4741_14889 n2_4741_14922 2.095238e-02
R7443 n2_4741_14922 n2_4741_15049 8.063492e-02
R7444 n2_4741_15138 n2_4741_15145 4.444444e-03
R7445 n2_4741_15145 n2_4741_15321 1.117460e-01
R7446 n2_4741_15321 n2_4741_15354 2.095238e-02
R7447 n2_4741_15354 n2_4741_15368 8.888889e-03
R7448 n2_4741_15368 n2_4741_15537 1.073016e-01
R7449 n2_4741_15537 n2_4741_15570 2.095238e-02
R7450 n2_4741_15570 n2_4741_15584 8.888889e-03
R7451 n2_4741_15584 n2_4741_15753 1.073016e-01
R7452 n2_4741_15753 n2_4741_15786 2.095238e-02
R7453 n2_4741_15786 n2_4741_15969 1.161905e-01
R7454 n2_4741_15969 n2_4741_16002 2.095238e-02
R7455 n2_4741_16002 n2_4741_16016 8.888889e-03
R7456 n2_4741_16016 n2_4741_16185 1.073016e-01
R7457 n2_4741_6049 n2_4880_6049 8.825397e-02
R7458 n2_4880_6049 n2_4929_6049 3.111111e-02
R7459 n2_4741_6145 n2_4880_6145 8.825397e-02
R7460 n2_4880_6145 n2_4929_6145 3.111111e-02
R7461 n2_4741_8299 n2_4880_8299 8.825397e-02
R7462 n2_4880_8299 n2_4929_8299 3.111111e-02
R7463 n2_4741_8395 n2_4880_8395 8.825397e-02
R7464 n2_4880_8395 n2_4929_8395 3.111111e-02
R7465 n2_4741_10549 n2_4880_10549 8.825397e-02
R7466 n2_4880_10549 n2_4929_10549 3.111111e-02
R7467 n2_4741_10645 n2_4880_10645 8.825397e-02
R7468 n2_4880_10645 n2_4929_10645 3.111111e-02
R7469 n2_4741_12799 n2_4880_12799 8.825397e-02
R7470 n2_4880_12799 n2_4929_12799 3.111111e-02
R7471 n2_4741_12895 n2_4880_12895 8.825397e-02
R7472 n2_4880_12895 n2_4929_12895 3.111111e-02
R7473 n2_4741_15049 n2_4880_15049 8.825397e-02
R7474 n2_4880_15049 n2_4929_15049 3.111111e-02
R7475 n2_4741_15145 n2_4880_15145 8.825397e-02
R7476 n2_4880_15145 n2_4929_15145 3.111111e-02
R7477 n2_4929_5169 n2_4929_5202 2.095238e-02
R7478 n2_4929_5202 n2_4929_5385 1.161905e-01
R7479 n2_4929_5385 n2_4929_5418 2.095238e-02
R7480 n2_4929_5418 n2_4929_5432 8.888889e-03
R7481 n2_4929_5432 n2_4929_5601 1.073016e-01
R7482 n2_4929_5601 n2_4929_5634 2.095238e-02
R7483 n2_4929_5634 n2_4929_5817 1.161905e-01
R7484 n2_4929_5817 n2_4929_5850 2.095238e-02
R7485 n2_4929_5850 n2_4929_6033 1.161905e-01
R7486 n2_4929_6033 n2_4929_6049 1.015873e-02
R7487 n2_4929_6049 n2_4929_6066 1.079365e-02
R7488 n2_4929_6066 n2_4929_6145 5.015873e-02
R7489 n2_4929_6145 n2_4929_6249 6.603175e-02
R7490 n2_4929_6249 n2_4929_6282 2.095238e-02
R7491 n2_4929_6282 n2_4929_6465 1.161905e-01
R7492 n2_4929_6465 n2_4929_6498 2.095238e-02
R7493 n2_4929_6498 n2_4929_6535 2.349206e-02
R7494 n2_4929_6535 n2_4929_6681 9.269841e-02
R7495 n2_4929_6681 n2_4929_6714 2.095238e-02
R7496 n2_4929_6714 n2_4929_6897 1.161905e-01
R7497 n2_4929_6897 n2_4929_6930 2.095238e-02
R7498 n2_4929_6930 n2_4929_7113 1.161905e-01
R7499 n2_4929_7329 n2_4929_7362 2.095238e-02
R7500 n2_4929_7362 n2_4929_7545 1.161905e-01
R7501 n2_4929_7545 n2_4929_7578 2.095238e-02
R7502 n2_4929_7578 n2_4929_7761 1.161905e-01
R7503 n2_4929_7761 n2_4929_7794 2.095238e-02
R7504 n2_4929_7794 n2_4929_7808 8.888889e-03
R7505 n2_4929_7808 n2_4929_7977 1.073016e-01
R7506 n2_4929_7977 n2_4929_8010 2.095238e-02
R7507 n2_4929_8010 n2_4929_8193 1.161905e-01
R7508 n2_4929_8193 n2_4929_8226 2.095238e-02
R7509 n2_4929_8226 n2_4929_8299 4.634921e-02
R7510 n2_4929_8299 n2_4929_8395 6.095238e-02
R7511 n2_4929_8395 n2_4929_8409 8.888889e-03
R7512 n2_4929_8409 n2_4929_8442 2.095238e-02
R7513 n2_4929_8442 n2_4929_8625 1.161905e-01
R7514 n2_4929_8625 n2_4929_8658 2.095238e-02
R7515 n2_4929_8658 n2_4929_8841 1.161905e-01
R7516 n2_4929_8841 n2_4929_8874 2.095238e-02
R7517 n2_4929_8874 n2_4929_8888 8.888889e-03
R7518 n2_4929_8888 n2_4929_8911 1.460317e-02
R7519 n2_4929_8911 n2_4929_9057 9.269841e-02
R7520 n2_4929_9057 n2_4929_9090 2.095238e-02
R7521 n2_4929_9090 n2_4929_9273 1.161905e-01
R7522 n2_4929_9273 n2_4929_9306 2.095238e-02
R7523 n2_4929_9705 n2_4929_9738 2.095238e-02
R7524 n2_4929_9738 n2_4929_9921 1.161905e-01
R7525 n2_4929_9921 n2_4929_9954 2.095238e-02
R7526 n2_4929_9954 n2_4929_9968 8.888889e-03
R7527 n2_4929_9968 n2_4929_10137 1.073016e-01
R7528 n2_4929_10137 n2_4929_10170 2.095238e-02
R7529 n2_4929_10170 n2_4929_10353 1.161905e-01
R7530 n2_4929_10353 n2_4929_10386 2.095238e-02
R7531 n2_4929_10386 n2_4929_10549 1.034921e-01
R7532 n2_4929_10549 n2_4929_10569 1.269841e-02
R7533 n2_4929_10569 n2_4929_10602 2.095238e-02
R7534 n2_4929_10602 n2_4929_10645 2.730159e-02
R7535 n2_4929_10645 n2_4929_10785 8.888889e-02
R7536 n2_4929_10785 n2_4929_10818 2.095238e-02
R7537 n2_4929_10818 n2_4929_11001 1.161905e-01
R7538 n2_4929_11001 n2_4929_11034 2.095238e-02
R7539 n2_4929_11034 n2_4929_11048 8.888889e-03
R7540 n2_4929_11048 n2_4929_11071 1.460317e-02
R7541 n2_4929_11071 n2_4929_11217 9.269841e-02
R7542 n2_4929_11217 n2_4929_11250 2.095238e-02
R7543 n2_4929_11250 n2_4929_11433 1.161905e-01
R7544 n2_4929_11433 n2_4929_11466 2.095238e-02
R7545 n2_4929_11865 n2_4929_11898 2.095238e-02
R7546 n2_4929_11898 n2_4929_12081 1.161905e-01
R7547 n2_4929_12081 n2_4929_12114 2.095238e-02
R7548 n2_4929_12114 n2_4929_12128 8.888889e-03
R7549 n2_4929_12128 n2_4929_12297 1.073016e-01
R7550 n2_4929_12297 n2_4929_12330 2.095238e-02
R7551 n2_4929_12330 n2_4929_12513 1.161905e-01
R7552 n2_4929_12513 n2_4929_12546 2.095238e-02
R7553 n2_4929_12546 n2_4929_12729 1.161905e-01
R7554 n2_4929_12729 n2_4929_12762 2.095238e-02
R7555 n2_4929_12762 n2_4929_12799 2.349206e-02
R7556 n2_4929_12799 n2_4929_12895 6.095238e-02
R7557 n2_4929_12895 n2_4929_12945 3.174603e-02
R7558 n2_4929_12945 n2_4929_12978 2.095238e-02
R7559 n2_4929_12978 n2_4929_13161 1.161905e-01
R7560 n2_4929_13161 n2_4929_13194 2.095238e-02
R7561 n2_4929_13194 n2_4929_13377 1.161905e-01
R7562 n2_4929_13377 n2_4929_13410 2.095238e-02
R7563 n2_4929_13410 n2_4929_13424 8.888889e-03
R7564 n2_4929_13424 n2_4929_13593 1.073016e-01
R7565 n2_4929_13593 n2_4929_13626 2.095238e-02
R7566 n2_4929_13626 n2_4929_13809 1.161905e-01
R7567 n2_4929_13809 n2_4929_13842 2.095238e-02
R7568 n2_4929_14100 n2_4929_14241 8.952381e-02
R7569 n2_4929_14241 n2_4929_14274 2.095238e-02
R7570 n2_4929_14274 n2_4929_14457 1.161905e-01
R7571 n2_4929_14457 n2_4929_14490 2.095238e-02
R7572 n2_4929_14490 n2_4929_14536 2.920635e-02
R7573 n2_4929_14536 n2_4929_14673 8.698413e-02
R7574 n2_4929_14673 n2_4929_14706 2.095238e-02
R7575 n2_4929_14706 n2_4929_14889 1.161905e-01
R7576 n2_4929_14889 n2_4929_14922 2.095238e-02
R7577 n2_4929_14922 n2_4929_15049 8.063492e-02
R7578 n2_4929_15049 n2_4929_15105 3.555556e-02
R7579 n2_4929_15105 n2_4929_15138 2.095238e-02
R7580 n2_4929_15138 n2_4929_15145 4.444444e-03
R7581 n2_4929_15145 n2_4929_15321 1.117460e-01
R7582 n2_4929_15321 n2_4929_15354 2.095238e-02
R7583 n2_4929_15354 n2_4929_15368 8.888889e-03
R7584 n2_4929_15368 n2_4929_15537 1.073016e-01
R7585 n2_4929_15537 n2_4929_15570 2.095238e-02
R7586 n2_4929_15570 n2_4929_15584 8.888889e-03
R7587 n2_4929_15584 n2_4929_15753 1.073016e-01
R7588 n2_4929_15753 n2_4929_15786 2.095238e-02
R7589 n2_4929_15786 n2_4929_15969 1.161905e-01
R7590 n2_4929_15969 n2_4929_16002 2.095238e-02
R7591 n2_4929_16002 n2_4929_16016 8.888889e-03
R7592 n2_5866_201 n2_5866_234 2.095238e-02
R7593 n2_5866_234 n2_5866_356 7.746032e-02
R7594 n2_5866_356 n2_5866_417 3.873016e-02
R7595 n2_5866_417 n2_5866_424 4.444444e-03
R7596 n2_5866_424 n2_5866_450 1.650794e-02
R7597 n2_5866_520 n2_5866_633 7.174603e-02
R7598 n2_5866_633 n2_5866_666 2.095238e-02
R7599 n2_5866_666 n2_5866_788 7.746032e-02
R7600 n2_5866_788 n2_5866_849 3.873016e-02
R7601 n2_5866_849 n2_5866_882 2.095238e-02
R7602 n2_5866_882 n2_5866_1065 1.161905e-01
R7603 n2_5866_1065 n2_5866_1098 2.095238e-02
R7604 n2_5866_1098 n2_5866_1281 1.161905e-01
R7605 n2_5866_1281 n2_5866_1314 2.095238e-02
R7606 n2_5866_1314 n2_5866_1497 1.161905e-01
R7607 n2_5866_1497 n2_5866_1530 2.095238e-02
R7608 n2_5866_1530 n2_5866_1549 1.206349e-02
R7609 n2_5866_1645 n2_5866_1713 4.317460e-02
R7610 n2_5866_1713 n2_5866_1746 2.095238e-02
R7611 n2_5866_1746 n2_5866_1760 8.888889e-03
R7612 n2_5866_1760 n2_5866_1929 1.073016e-01
R7613 n2_5866_1929 n2_5866_1962 2.095238e-02
R7614 n2_5866_1962 n2_5866_2145 1.161905e-01
R7615 n2_5866_2145 n2_5866_2178 2.095238e-02
R7616 n2_5866_2178 n2_5866_2361 1.161905e-01
R7617 n2_5866_2361 n2_5866_2394 2.095238e-02
R7618 n2_5866_2394 n2_5866_2408 8.888889e-03
R7619 n2_5866_2408 n2_5866_2577 1.073016e-01
R7620 n2_5866_2577 n2_5866_2610 2.095238e-02
R7621 n2_5866_2610 n2_5866_2674 4.063492e-02
R7622 n2_5866_2770 n2_5866_2793 1.460317e-02
R7623 n2_5866_2793 n2_5866_2826 2.095238e-02
R7624 n2_5866_2826 n2_5866_2840 8.888889e-03
R7625 n2_5866_2840 n2_5866_3009 1.073016e-01
R7626 n2_5866_3009 n2_5866_3042 2.095238e-02
R7627 n2_5866_3042 n2_5866_3056 8.888889e-03
R7628 n2_5866_3056 n2_5866_3225 1.073016e-01
R7629 n2_5866_3225 n2_5866_3258 2.095238e-02
R7630 n2_5866_3258 n2_5866_3441 1.161905e-01
R7631 n2_5866_3441 n2_5866_3474 2.095238e-02
R7632 n2_5866_3474 n2_5866_3488 8.888889e-03
R7633 n2_5866_3488 n2_5866_3657 1.073016e-01
R7634 n2_5866_3657 n2_5866_3690 2.095238e-02
R7635 n2_5866_3690 n2_5866_3799 6.920635e-02
R7636 n2_5866_3873 n2_5866_3895 1.396825e-02
R7637 n2_5866_3895 n2_5866_3906 6.984127e-03
R7638 n2_5866_3906 n2_5866_4089 1.161905e-01
R7639 n2_5866_4089 n2_5866_4122 2.095238e-02
R7640 n2_5866_4122 n2_5866_4136 8.888889e-03
R7641 n2_5866_4136 n2_5866_4305 1.073016e-01
R7642 n2_5866_4305 n2_5866_4338 2.095238e-02
R7643 n2_5866_4338 n2_5866_4352 8.888889e-03
R7644 n2_5866_4352 n2_5866_4375 1.460317e-02
R7645 n2_5866_4375 n2_5866_4521 9.269841e-02
R7646 n2_5866_4521 n2_5866_4554 2.095238e-02
R7647 n2_5866_4554 n2_5866_4568 8.888889e-03
R7648 n2_5866_4568 n2_5866_4737 1.073016e-01
R7649 n2_5866_4737 n2_5866_4770 2.095238e-02
R7650 n2_5866_4770 n2_5866_4924 9.777778e-02
R7651 n2_5866_4924 n2_5866_4953 1.841270e-02
R7652 n2_5866_5020 n2_5866_5169 9.460317e-02
R7653 n2_5866_5169 n2_5866_5202 2.095238e-02
R7654 n2_5866_5202 n2_5866_5216 8.888889e-03
R7655 n2_5866_5216 n2_5866_5385 1.073016e-01
R7656 n2_5866_5385 n2_5866_5418 2.095238e-02
R7657 n2_5866_5418 n2_5866_5432 8.888889e-03
R7658 n2_5866_5432 n2_5866_5455 1.460317e-02
R7659 n2_5866_5455 n2_5866_5601 9.269841e-02
R7660 n2_5866_5601 n2_5866_5634 2.095238e-02
R7661 n2_5866_5634 n2_5866_5817 1.161905e-01
R7662 n2_5866_5817 n2_5866_5850 2.095238e-02
R7663 n2_5866_5850 n2_5866_6033 1.161905e-01
R7664 n2_5866_6033 n2_5866_6049 1.015873e-02
R7665 n2_5866_6049 n2_5866_6066 1.079365e-02
R7666 n2_5866_6145 n2_5866_6249 6.603175e-02
R7667 n2_5866_6249 n2_5866_6282 2.095238e-02
R7668 n2_5866_6282 n2_5866_6465 1.161905e-01
R7669 n2_5866_6465 n2_5866_6498 2.095238e-02
R7670 n2_5866_6498 n2_5866_6535 2.349206e-02
R7671 n2_5866_6535 n2_5866_6681 9.269841e-02
R7672 n2_5866_6681 n2_5866_6714 2.095238e-02
R7673 n2_5866_6714 n2_5866_6897 1.161905e-01
R7674 n2_5866_6897 n2_5866_6930 2.095238e-02
R7675 n2_5866_6930 n2_5866_7113 1.161905e-01
R7676 n2_5866_7113 n2_5866_7146 2.095238e-02
R7677 n2_5866_7146 n2_5866_7329 1.161905e-01
R7678 n2_5866_7329 n2_5866_7362 2.095238e-02
R7679 n2_5866_7362 n2_5866_7545 1.161905e-01
R7680 n2_5866_7545 n2_5866_7578 2.095238e-02
R7681 n2_5866_7578 n2_5866_7761 1.161905e-01
R7682 n2_5866_7761 n2_5866_7794 2.095238e-02
R7683 n2_5866_7794 n2_5866_7808 8.888889e-03
R7684 n2_5866_7808 n2_5866_7977 1.073016e-01
R7685 n2_5866_7977 n2_5866_8010 2.095238e-02
R7686 n2_5866_8010 n2_5866_8193 1.161905e-01
R7687 n2_5866_8193 n2_5866_8226 2.095238e-02
R7688 n2_5866_8226 n2_5866_8299 4.634921e-02
R7689 n2_5866_8395 n2_5866_8409 8.888889e-03
R7690 n2_5866_8409 n2_5866_8442 2.095238e-02
R7691 n2_5866_8442 n2_5866_8625 1.161905e-01
R7692 n2_5866_8625 n2_5866_8658 2.095238e-02
R7693 n2_5866_8658 n2_5866_8841 1.161905e-01
R7694 n2_5866_8841 n2_5866_8874 2.095238e-02
R7695 n2_5866_8874 n2_5866_8888 8.888889e-03
R7696 n2_5866_8888 n2_5866_8911 1.460317e-02
R7697 n2_5866_8911 n2_5866_9057 9.269841e-02
R7698 n2_5866_9057 n2_5866_9090 2.095238e-02
R7699 n2_5866_9090 n2_5866_9273 1.161905e-01
R7700 n2_5866_9273 n2_5866_9306 2.095238e-02
R7701 n2_5866_9306 n2_5866_9489 1.161905e-01
R7702 n2_5866_9489 n2_5866_9522 2.095238e-02
R7703 n2_5866_9522 n2_5866_9705 1.161905e-01
R7704 n2_5866_9705 n2_5866_9738 2.095238e-02
R7705 n2_5866_9738 n2_5866_9921 1.161905e-01
R7706 n2_5866_9921 n2_5866_9954 2.095238e-02
R7707 n2_5866_9954 n2_5866_9968 8.888889e-03
R7708 n2_5866_9968 n2_5866_10137 1.073016e-01
R7709 n2_5866_10137 n2_5866_10170 2.095238e-02
R7710 n2_5866_10170 n2_5866_10353 1.161905e-01
R7711 n2_5866_10353 n2_5866_10386 2.095238e-02
R7712 n2_5866_10386 n2_5866_10549 1.034921e-01
R7713 n2_5866_10549 n2_5866_10569 1.269841e-02
R7714 n2_5866_10645 n2_5866_10785 8.888889e-02
R7715 n2_5866_10785 n2_5866_10818 2.095238e-02
R7716 n2_5866_10818 n2_5866_11001 1.161905e-01
R7717 n2_5866_11001 n2_5866_11034 2.095238e-02
R7718 n2_5866_11034 n2_5866_11048 8.888889e-03
R7719 n2_5866_11048 n2_5866_11071 1.460317e-02
R7720 n2_5866_11071 n2_5866_11217 9.269841e-02
R7721 n2_5866_11217 n2_5866_11250 2.095238e-02
R7722 n2_5866_11250 n2_5866_11433 1.161905e-01
R7723 n2_5866_11433 n2_5866_11466 2.095238e-02
R7724 n2_5866_11466 n2_5866_11649 1.161905e-01
R7725 n2_5866_11649 n2_5866_11682 2.095238e-02
R7726 n2_5866_11682 n2_5866_11865 1.161905e-01
R7727 n2_5866_11865 n2_5866_11898 2.095238e-02
R7728 n2_5866_11898 n2_5866_12081 1.161905e-01
R7729 n2_5866_12081 n2_5866_12114 2.095238e-02
R7730 n2_5866_12114 n2_5866_12128 8.888889e-03
R7731 n2_5866_12128 n2_5866_12297 1.073016e-01
R7732 n2_5866_12297 n2_5866_12330 2.095238e-02
R7733 n2_5866_12330 n2_5866_12513 1.161905e-01
R7734 n2_5866_12513 n2_5866_12546 2.095238e-02
R7735 n2_5866_12546 n2_5866_12729 1.161905e-01
R7736 n2_5866_12729 n2_5866_12762 2.095238e-02
R7737 n2_5866_12762 n2_5866_12799 2.349206e-02
R7738 n2_5866_12895 n2_5866_12945 3.174603e-02
R7739 n2_5866_12945 n2_5866_12978 2.095238e-02
R7740 n2_5866_12978 n2_5866_13161 1.161905e-01
R7741 n2_5866_13161 n2_5866_13194 2.095238e-02
R7742 n2_5866_13194 n2_5866_13377 1.161905e-01
R7743 n2_5866_13377 n2_5866_13410 2.095238e-02
R7744 n2_5866_13410 n2_5866_13424 8.888889e-03
R7745 n2_5866_13424 n2_5866_13593 1.073016e-01
R7746 n2_5866_13593 n2_5866_13626 2.095238e-02
R7747 n2_5866_13626 n2_5866_13809 1.161905e-01
R7748 n2_5866_13809 n2_5866_13842 2.095238e-02
R7749 n2_5866_13842 n2_5866_13879 2.349206e-02
R7750 n2_5866_13879 n2_5866_14025 9.269841e-02
R7751 n2_5866_14025 n2_5866_14058 2.095238e-02
R7752 n2_5866_14058 n2_5866_14241 1.161905e-01
R7753 n2_5866_14241 n2_5866_14274 2.095238e-02
R7754 n2_5866_14274 n2_5866_14457 1.161905e-01
R7755 n2_5866_14457 n2_5866_14490 2.095238e-02
R7756 n2_5866_14490 n2_5866_14536 2.920635e-02
R7757 n2_5866_14536 n2_5866_14673 8.698413e-02
R7758 n2_5866_14673 n2_5866_14706 2.095238e-02
R7759 n2_5866_14706 n2_5866_14889 1.161905e-01
R7760 n2_5866_14889 n2_5866_14922 2.095238e-02
R7761 n2_5866_14922 n2_5866_15049 8.063492e-02
R7762 n2_5866_15138 n2_5866_15145 4.444444e-03
R7763 n2_5866_15145 n2_5866_15321 1.117460e-01
R7764 n2_5866_15321 n2_5866_15354 2.095238e-02
R7765 n2_5866_15354 n2_5866_15537 1.161905e-01
R7766 n2_5866_15537 n2_5866_15570 2.095238e-02
R7767 n2_5866_15570 n2_5866_15584 8.888889e-03
R7768 n2_5866_15584 n2_5866_15753 1.073016e-01
R7769 n2_5866_15753 n2_5866_15786 2.095238e-02
R7770 n2_5866_15786 n2_5866_15800 8.888889e-03
R7771 n2_5866_15800 n2_5866_15969 1.073016e-01
R7772 n2_5866_15969 n2_5866_16002 2.095238e-02
R7773 n2_5866_16002 n2_5866_16016 8.888889e-03
R7774 n2_5866_16016 n2_5866_16174 1.003175e-01
R7775 n2_5866_16174 n2_5866_16185 6.984127e-03
R7776 n2_5866_16270 n2_5866_16401 8.317460e-02
R7777 n2_5866_16401 n2_5866_16434 2.095238e-02
R7778 n2_5866_16434 n2_5866_16617 1.161905e-01
R7779 n2_5866_16617 n2_5866_16650 2.095238e-02
R7780 n2_5866_16650 n2_5866_16833 1.161905e-01
R7781 n2_5866_16833 n2_5866_16866 2.095238e-02
R7782 n2_5866_16866 n2_5866_17049 1.161905e-01
R7783 n2_5866_17049 n2_5866_17082 2.095238e-02
R7784 n2_5866_17082 n2_5866_17096 8.888889e-03
R7785 n2_5866_17096 n2_5866_17119 1.460317e-02
R7786 n2_5866_17119 n2_5866_17265 9.269841e-02
R7787 n2_5866_17265 n2_5866_17298 2.095238e-02
R7788 n2_5866_17298 n2_5866_17299 6.349206e-04
R7789 n2_5866_17299 n2_5866_17312 8.253968e-03
R7790 n2_5866_17395 n2_5866_17481 5.460317e-02
R7791 n2_5866_17481 n2_5866_17514 2.095238e-02
R7792 n2_5866_17514 n2_5866_17528 8.888889e-03
R7793 n2_5866_17528 n2_5866_17697 1.073016e-01
R7794 n2_5866_17697 n2_5866_17730 2.095238e-02
R7795 n2_5866_17730 n2_5866_17913 1.161905e-01
R7796 n2_5866_17913 n2_5866_17946 2.095238e-02
R7797 n2_5866_17946 n2_5866_18129 1.161905e-01
R7798 n2_5866_18129 n2_5866_18162 2.095238e-02
R7799 n2_5866_18162 n2_5866_18345 1.161905e-01
R7800 n2_5866_18345 n2_5866_18378 2.095238e-02
R7801 n2_5866_18378 n2_5866_18392 8.888889e-03
R7802 n2_5866_18392 n2_5866_18424 2.031746e-02
R7803 n2_5866_18520 n2_5866_18561 2.603175e-02
R7804 n2_5866_18561 n2_5866_18594 2.095238e-02
R7805 n2_5866_18594 n2_5866_18608 8.888889e-03
R7806 n2_5866_18608 n2_5866_18777 1.073016e-01
R7807 n2_5866_18777 n2_5866_18810 2.095238e-02
R7808 n2_5866_18810 n2_5866_18824 8.888889e-03
R7809 n2_5866_18824 n2_5866_18993 1.073016e-01
R7810 n2_5866_18993 n2_5866_19026 2.095238e-02
R7811 n2_5866_19026 n2_5866_19040 8.888889e-03
R7812 n2_5866_19040 n2_5866_19209 1.073016e-01
R7813 n2_5866_19209 n2_5866_19242 2.095238e-02
R7814 n2_5866_19242 n2_5866_19425 1.161905e-01
R7815 n2_5866_19425 n2_5866_19458 2.095238e-02
R7816 n2_5866_19458 n2_5866_19472 8.888889e-03
R7817 n2_5866_19472 n2_5866_19549 4.888889e-02
R7818 n2_5866_19641 n2_5866_19645 2.539683e-03
R7819 n2_5866_19645 n2_5866_19674 1.841270e-02
R7820 n2_5866_19674 n2_5866_19857 1.161905e-01
R7821 n2_5866_19857 n2_5866_19890 2.095238e-02
R7822 n2_5866_19890 n2_5866_20073 1.161905e-01
R7823 n2_5866_20073 n2_5866_20106 2.095238e-02
R7824 n2_5866_20106 n2_5866_20289 1.161905e-01
R7825 n2_5866_20289 n2_5866_20322 2.095238e-02
R7826 n2_5866_20322 n2_5866_20505 1.161905e-01
R7827 n2_5866_20505 n2_5866_20538 2.095238e-02
R7828 n2_5866_20538 n2_5866_20674 8.634921e-02
R7829 n2_5866_20754 n2_5866_20770 1.015873e-02
R7830 n2_5866_20770 n2_5866_20937 1.060317e-01
R7831 n2_5866_20937 n2_5866_20970 2.095238e-02
R7832 n2_5866_6145 n2_5958_6145 5.841270e-02
R7833 n2_5958_6145 n2_6005_6145 2.984127e-02
R7834 n2_6005_6145 n2_6054_6145 3.111111e-02
R7835 n2_5866_8299 n2_6005_8299 8.825397e-02
R7836 n2_6005_8299 n2_6054_8299 3.111111e-02
R7837 n2_5866_8395 n2_6005_8395 8.825397e-02
R7838 n2_6005_8395 n2_6054_8395 3.111111e-02
R7839 n2_5866_10549 n2_6005_10549 8.825397e-02
R7840 n2_6005_10549 n2_6054_10549 3.111111e-02
R7841 n2_5866_10645 n2_6005_10645 8.825397e-02
R7842 n2_6005_10645 n2_6054_10645 3.111111e-02
R7843 n2_5866_12799 n2_6005_12799 8.825397e-02
R7844 n2_6005_12799 n2_6054_12799 3.111111e-02
R7845 n2_5866_12895 n2_6005_12895 8.825397e-02
R7846 n2_6005_12895 n2_6054_12895 3.111111e-02
R7847 n2_5866_15049 n2_5958_15049 5.841270e-02
R7848 n2_5958_15049 n2_6005_15049 2.984127e-02
R7849 n2_6005_15049 n2_6054_15049 3.111111e-02
R7850 n2_5866_424 n2_5958_424 5.841270e-02
R7851 n2_5958_424 n2_6005_424 2.984127e-02
R7852 n2_6005_424 n2_6054_424 3.111111e-02
R7853 n2_6054_424 n2_6146_424 5.841270e-02
R7854 n2_5866_520 n2_5958_520 5.841270e-02
R7855 n2_5958_520 n2_6005_520 2.984127e-02
R7856 n2_6005_520 n2_6054_520 3.111111e-02
R7857 n2_6054_520 n2_6146_520 5.841270e-02
R7858 n2_5866_1549 n2_5958_1549 5.841270e-02
R7859 n2_5958_1549 n2_6005_1549 2.984127e-02
R7860 n2_6005_1549 n2_6054_1549 3.111111e-02
R7861 n2_6054_1549 n2_6146_1549 5.841270e-02
R7862 n2_5866_1645 n2_5958_1645 5.841270e-02
R7863 n2_5958_1645 n2_6005_1645 2.984127e-02
R7864 n2_6005_1645 n2_6054_1645 3.111111e-02
R7865 n2_6054_1645 n2_6146_1645 5.841270e-02
R7866 n2_5866_2674 n2_5958_2674 5.841270e-02
R7867 n2_5958_2674 n2_6005_2674 2.984127e-02
R7868 n2_6005_2674 n2_6054_2674 3.111111e-02
R7869 n2_6054_2674 n2_6146_2674 5.841270e-02
R7870 n2_5866_2770 n2_5958_2770 5.841270e-02
R7871 n2_5958_2770 n2_6005_2770 2.984127e-02
R7872 n2_6005_2770 n2_6054_2770 3.111111e-02
R7873 n2_6054_2770 n2_6146_2770 5.841270e-02
R7874 n2_5866_3799 n2_5958_3799 5.841270e-02
R7875 n2_5958_3799 n2_6005_3799 2.984127e-02
R7876 n2_6005_3799 n2_6054_3799 3.111111e-02
R7877 n2_6054_3799 n2_6146_3799 5.841270e-02
R7878 n2_5866_3895 n2_5958_3895 5.841270e-02
R7879 n2_5958_3895 n2_6005_3895 2.984127e-02
R7880 n2_6005_3895 n2_6054_3895 3.111111e-02
R7881 n2_6054_3895 n2_6146_3895 5.841270e-02
R7882 n2_5866_4924 n2_5958_4924 5.841270e-02
R7883 n2_5958_4924 n2_6005_4924 2.984127e-02
R7884 n2_6005_4924 n2_6054_4924 3.111111e-02
R7885 n2_6054_4924 n2_6146_4924 5.841270e-02
R7886 n2_5866_5020 n2_5958_5020 5.841270e-02
R7887 n2_5958_5020 n2_6005_5020 2.984127e-02
R7888 n2_6005_5020 n2_6054_5020 3.111111e-02
R7889 n2_6054_5020 n2_6146_5020 5.841270e-02
R7890 n2_5866_6049 n2_5958_6049 5.841270e-02
R7891 n2_5958_6049 n2_6005_6049 2.984127e-02
R7892 n2_6005_6049 n2_6054_6049 3.111111e-02
R7893 n2_6054_6049 n2_6146_6049 5.841270e-02
R7894 n2_5866_15145 n2_5958_15145 5.841270e-02
R7895 n2_5958_15145 n2_6005_15145 2.984127e-02
R7896 n2_6005_15145 n2_6054_15145 3.111111e-02
R7897 n2_6054_15145 n2_6146_15145 5.841270e-02
R7898 n2_5866_16174 n2_5958_16174 5.841270e-02
R7899 n2_5958_16174 n2_6005_16174 2.984127e-02
R7900 n2_6005_16174 n2_6054_16174 3.111111e-02
R7901 n2_6054_16174 n2_6146_16174 5.841270e-02
R7902 n2_5866_16270 n2_5958_16270 5.841270e-02
R7903 n2_5958_16270 n2_6005_16270 2.984127e-02
R7904 n2_6005_16270 n2_6054_16270 3.111111e-02
R7905 n2_6054_16270 n2_6146_16270 5.841270e-02
R7906 n2_5866_17299 n2_5958_17299 5.841270e-02
R7907 n2_5958_17299 n2_6005_17299 2.984127e-02
R7908 n2_6005_17299 n2_6054_17299 3.111111e-02
R7909 n2_6054_17299 n2_6146_17299 5.841270e-02
R7910 n2_5866_17395 n2_5958_17395 5.841270e-02
R7911 n2_5958_17395 n2_6005_17395 2.984127e-02
R7912 n2_6005_17395 n2_6054_17395 3.111111e-02
R7913 n2_6054_17395 n2_6146_17395 5.841270e-02
R7914 n2_5866_18424 n2_5958_18424 5.841270e-02
R7915 n2_5958_18424 n2_6005_18424 2.984127e-02
R7916 n2_6005_18424 n2_6054_18424 3.111111e-02
R7917 n2_6054_18424 n2_6146_18424 5.841270e-02
R7918 n2_5866_18520 n2_5958_18520 5.841270e-02
R7919 n2_5958_18520 n2_6005_18520 2.984127e-02
R7920 n2_6005_18520 n2_6054_18520 3.111111e-02
R7921 n2_6054_18520 n2_6146_18520 5.841270e-02
R7922 n2_5866_19549 n2_5958_19549 5.841270e-02
R7923 n2_5958_19549 n2_6005_19549 2.984127e-02
R7924 n2_6005_19549 n2_6054_19549 3.111111e-02
R7925 n2_6054_19549 n2_6146_19549 5.841270e-02
R7926 n2_5866_19645 n2_5958_19645 5.841270e-02
R7927 n2_5958_19645 n2_6005_19645 2.984127e-02
R7928 n2_6005_19645 n2_6054_19645 3.111111e-02
R7929 n2_6054_19645 n2_6146_19645 5.841270e-02
R7930 n2_5866_20674 n2_5958_20674 5.841270e-02
R7931 n2_5958_20674 n2_6005_20674 2.984127e-02
R7932 n2_6005_20674 n2_6054_20674 3.111111e-02
R7933 n2_6054_20674 n2_6146_20674 5.841270e-02
R7934 n2_5866_20770 n2_5958_20770 5.841270e-02
R7935 n2_5958_20770 n2_6005_20770 2.984127e-02
R7936 n2_6005_20770 n2_6054_20770 3.111111e-02
R7937 n2_6054_20770 n2_6146_20770 5.841270e-02
R7938 n2_5958_201 n2_5958_234 2.095238e-02
R7939 n2_5958_234 n2_5958_356 7.746032e-02
R7940 n2_5958_356 n2_5958_417 3.873016e-02
R7941 n2_5958_417 n2_5958_424 4.444444e-03
R7942 n2_5958_424 n2_5958_450 1.650794e-02
R7943 n2_5958_450 n2_5958_520 4.444444e-02
R7944 n2_5958_520 n2_5958_633 7.174603e-02
R7945 n2_5958_633 n2_5958_666 2.095238e-02
R7946 n2_5958_666 n2_5958_788 7.746032e-02
R7947 n2_5958_788 n2_5958_849 3.873016e-02
R7948 n2_5958_849 n2_5958_882 2.095238e-02
R7949 n2_5958_882 n2_5958_1065 1.161905e-01
R7950 n2_5958_1065 n2_5958_1098 2.095238e-02
R7951 n2_5958_1098 n2_5958_1281 1.161905e-01
R7952 n2_5958_1281 n2_5958_1314 2.095238e-02
R7953 n2_5958_1314 n2_5958_1497 1.161905e-01
R7954 n2_5958_1497 n2_5958_1530 2.095238e-02
R7955 n2_5958_1530 n2_5958_1549 1.206349e-02
R7956 n2_5958_1549 n2_5958_1645 6.095238e-02
R7957 n2_5958_1645 n2_5958_1713 4.317460e-02
R7958 n2_5958_1713 n2_5958_1746 2.095238e-02
R7959 n2_5958_1746 n2_5958_1760 8.888889e-03
R7960 n2_5958_1760 n2_5958_1929 1.073016e-01
R7961 n2_5958_1929 n2_5958_1962 2.095238e-02
R7962 n2_5958_1962 n2_5958_2145 1.161905e-01
R7963 n2_5958_2145 n2_5958_2178 2.095238e-02
R7964 n2_5958_2178 n2_5958_2361 1.161905e-01
R7965 n2_5958_2361 n2_5958_2394 2.095238e-02
R7966 n2_5958_2394 n2_5958_2408 8.888889e-03
R7967 n2_5958_2408 n2_5958_2577 1.073016e-01
R7968 n2_5958_2577 n2_5958_2610 2.095238e-02
R7969 n2_5958_2610 n2_5958_2674 4.063492e-02
R7970 n2_5958_2674 n2_5958_2770 6.095238e-02
R7971 n2_5958_2770 n2_5958_2793 1.460317e-02
R7972 n2_5958_2793 n2_5958_2826 2.095238e-02
R7973 n2_5958_2826 n2_5958_2840 8.888889e-03
R7974 n2_5958_2840 n2_5958_3009 1.073016e-01
R7975 n2_5958_3009 n2_5958_3042 2.095238e-02
R7976 n2_5958_3042 n2_5958_3056 8.888889e-03
R7977 n2_5958_3056 n2_5958_3225 1.073016e-01
R7978 n2_5958_3225 n2_5958_3258 2.095238e-02
R7979 n2_5958_3258 n2_5958_3441 1.161905e-01
R7980 n2_5958_3441 n2_5958_3474 2.095238e-02
R7981 n2_5958_3474 n2_5958_3488 8.888889e-03
R7982 n2_5958_3488 n2_5958_3657 1.073016e-01
R7983 n2_5958_3657 n2_5958_3690 2.095238e-02
R7984 n2_5958_3690 n2_5958_3799 6.920635e-02
R7985 n2_5958_3799 n2_5958_3873 4.698413e-02
R7986 n2_5958_3873 n2_5958_3895 1.396825e-02
R7987 n2_5958_3895 n2_5958_3906 6.984127e-03
R7988 n2_5958_3906 n2_5958_4089 1.161905e-01
R7989 n2_5958_4089 n2_5958_4122 2.095238e-02
R7990 n2_5958_4122 n2_5958_4136 8.888889e-03
R7991 n2_5958_4136 n2_5958_4305 1.073016e-01
R7992 n2_5958_4305 n2_5958_4338 2.095238e-02
R7993 n2_5958_4338 n2_5958_4352 8.888889e-03
R7994 n2_5958_4352 n2_5958_4375 1.460317e-02
R7995 n2_5958_4375 n2_5958_4521 9.269841e-02
R7996 n2_5958_4521 n2_5958_4554 2.095238e-02
R7997 n2_5958_4554 n2_5958_4568 8.888889e-03
R7998 n2_5958_4568 n2_5958_4737 1.073016e-01
R7999 n2_5958_4737 n2_5958_4770 2.095238e-02
R8000 n2_5958_4770 n2_5958_4924 9.777778e-02
R8001 n2_5958_4924 n2_5958_4953 1.841270e-02
R8002 n2_5958_4953 n2_5958_4986 2.095238e-02
R8003 n2_5958_4986 n2_5958_5020 2.158730e-02
R8004 n2_5958_5020 n2_5958_5169 9.460317e-02
R8005 n2_5958_5169 n2_5958_5202 2.095238e-02
R8006 n2_5958_5202 n2_5958_5216 8.888889e-03
R8007 n2_5958_5216 n2_5958_5385 1.073016e-01
R8008 n2_5958_5385 n2_5958_5418 2.095238e-02
R8009 n2_5958_5418 n2_5958_5432 8.888889e-03
R8010 n2_5958_5432 n2_5958_5455 1.460317e-02
R8011 n2_5958_5455 n2_5958_5601 9.269841e-02
R8012 n2_5958_5601 n2_5958_5634 2.095238e-02
R8013 n2_5958_5634 n2_5958_5817 1.161905e-01
R8014 n2_5958_5817 n2_5958_5850 2.095238e-02
R8015 n2_5958_5850 n2_5958_6033 1.161905e-01
R8016 n2_5958_6033 n2_5958_6049 1.015873e-02
R8017 n2_5958_6049 n2_5958_6066 1.079365e-02
R8018 n2_5958_6066 n2_5958_6145 5.015873e-02
R8019 n2_5958_15049 n2_5958_15105 3.555556e-02
R8020 n2_5958_15105 n2_5958_15138 2.095238e-02
R8021 n2_5958_15138 n2_5958_15145 4.444444e-03
R8022 n2_5958_15145 n2_5958_15321 1.117460e-01
R8023 n2_5958_15321 n2_5958_15354 2.095238e-02
R8024 n2_5958_15354 n2_5958_15537 1.161905e-01
R8025 n2_5958_15537 n2_5958_15570 2.095238e-02
R8026 n2_5958_15570 n2_5958_15584 8.888889e-03
R8027 n2_5958_15584 n2_5958_15753 1.073016e-01
R8028 n2_5958_15753 n2_5958_15786 2.095238e-02
R8029 n2_5958_15786 n2_5958_15800 8.888889e-03
R8030 n2_5958_15800 n2_5958_15969 1.073016e-01
R8031 n2_5958_15969 n2_5958_16002 2.095238e-02
R8032 n2_5958_16002 n2_5958_16016 8.888889e-03
R8033 n2_5958_16016 n2_5958_16174 1.003175e-01
R8034 n2_5958_16174 n2_5958_16185 6.984127e-03
R8035 n2_5958_16185 n2_5958_16218 2.095238e-02
R8036 n2_5958_16218 n2_5958_16270 3.301587e-02
R8037 n2_5958_16270 n2_5958_16401 8.317460e-02
R8038 n2_5958_16401 n2_5958_16434 2.095238e-02
R8039 n2_5958_16434 n2_5958_16617 1.161905e-01
R8040 n2_5958_16617 n2_5958_16650 2.095238e-02
R8041 n2_5958_16650 n2_5958_16833 1.161905e-01
R8042 n2_5958_16833 n2_5958_16866 2.095238e-02
R8043 n2_5958_16866 n2_5958_17049 1.161905e-01
R8044 n2_5958_17049 n2_5958_17082 2.095238e-02
R8045 n2_5958_17082 n2_5958_17096 8.888889e-03
R8046 n2_5958_17096 n2_5958_17119 1.460317e-02
R8047 n2_5958_17119 n2_5958_17265 9.269841e-02
R8048 n2_5958_17265 n2_5958_17298 2.095238e-02
R8049 n2_5958_17298 n2_5958_17299 6.349206e-04
R8050 n2_5958_17299 n2_5958_17312 8.253968e-03
R8051 n2_5958_17312 n2_5958_17335 1.460317e-02
R8052 n2_5958_17335 n2_5958_17395 3.809524e-02
R8053 n2_5958_17395 n2_5958_17481 5.460317e-02
R8054 n2_5958_17481 n2_5958_17514 2.095238e-02
R8055 n2_5958_17514 n2_5958_17528 8.888889e-03
R8056 n2_5958_17528 n2_5958_17697 1.073016e-01
R8057 n2_5958_17697 n2_5958_17730 2.095238e-02
R8058 n2_5958_17730 n2_5958_17913 1.161905e-01
R8059 n2_5958_17913 n2_5958_17946 2.095238e-02
R8060 n2_5958_17946 n2_5958_18129 1.161905e-01
R8061 n2_5958_18129 n2_5958_18162 2.095238e-02
R8062 n2_5958_18162 n2_5958_18345 1.161905e-01
R8063 n2_5958_18345 n2_5958_18378 2.095238e-02
R8064 n2_5958_18378 n2_5958_18392 8.888889e-03
R8065 n2_5958_18392 n2_5958_18424 2.031746e-02
R8066 n2_5958_18424 n2_5958_18520 6.095238e-02
R8067 n2_5958_18520 n2_5958_18561 2.603175e-02
R8068 n2_5958_18561 n2_5958_18594 2.095238e-02
R8069 n2_5958_18594 n2_5958_18608 8.888889e-03
R8070 n2_5958_18608 n2_5958_18777 1.073016e-01
R8071 n2_5958_18777 n2_5958_18810 2.095238e-02
R8072 n2_5958_18810 n2_5958_18824 8.888889e-03
R8073 n2_5958_18824 n2_5958_18993 1.073016e-01
R8074 n2_5958_18993 n2_5958_19026 2.095238e-02
R8075 n2_5958_19026 n2_5958_19040 8.888889e-03
R8076 n2_5958_19040 n2_5958_19209 1.073016e-01
R8077 n2_5958_19209 n2_5958_19242 2.095238e-02
R8078 n2_5958_19242 n2_5958_19425 1.161905e-01
R8079 n2_5958_19425 n2_5958_19458 2.095238e-02
R8080 n2_5958_19458 n2_5958_19472 8.888889e-03
R8081 n2_5958_19472 n2_5958_19549 4.888889e-02
R8082 n2_5958_19549 n2_5958_19641 5.841270e-02
R8083 n2_5958_19641 n2_5958_19645 2.539683e-03
R8084 n2_5958_19645 n2_5958_19674 1.841270e-02
R8085 n2_5958_19674 n2_5958_19857 1.161905e-01
R8086 n2_5958_19857 n2_5958_19890 2.095238e-02
R8087 n2_5958_19890 n2_5958_20073 1.161905e-01
R8088 n2_5958_20073 n2_5958_20106 2.095238e-02
R8089 n2_5958_20106 n2_5958_20289 1.161905e-01
R8090 n2_5958_20289 n2_5958_20322 2.095238e-02
R8091 n2_5958_20322 n2_5958_20505 1.161905e-01
R8092 n2_5958_20505 n2_5958_20538 2.095238e-02
R8093 n2_5958_20538 n2_5958_20674 8.634921e-02
R8094 n2_5958_20674 n2_5958_20721 2.984127e-02
R8095 n2_5958_20721 n2_5958_20754 2.095238e-02
R8096 n2_5958_20754 n2_5958_20770 1.015873e-02
R8097 n2_5958_20770 n2_5958_20937 1.060317e-01
R8098 n2_5958_20937 n2_5958_20970 2.095238e-02
R8099 n2_6054_201 n2_6054_234 2.095238e-02
R8100 n2_6054_234 n2_6054_356 7.746032e-02
R8101 n2_6054_356 n2_6054_417 3.873016e-02
R8102 n2_6054_417 n2_6054_424 4.444444e-03
R8103 n2_6054_424 n2_6054_450 1.650794e-02
R8104 n2_6054_450 n2_6054_520 4.444444e-02
R8105 n2_6054_520 n2_6054_633 7.174603e-02
R8106 n2_6054_633 n2_6054_666 2.095238e-02
R8107 n2_6054_666 n2_6054_788 7.746032e-02
R8108 n2_6054_788 n2_6054_849 3.873016e-02
R8109 n2_6054_849 n2_6054_882 2.095238e-02
R8110 n2_6054_882 n2_6054_1065 1.161905e-01
R8111 n2_6054_1065 n2_6054_1098 2.095238e-02
R8112 n2_6054_1098 n2_6054_1281 1.161905e-01
R8113 n2_6054_1281 n2_6054_1314 2.095238e-02
R8114 n2_6054_1314 n2_6054_1497 1.161905e-01
R8115 n2_6054_1497 n2_6054_1530 2.095238e-02
R8116 n2_6054_1530 n2_6054_1549 1.206349e-02
R8117 n2_6054_1549 n2_6054_1645 6.095238e-02
R8118 n2_6054_1645 n2_6054_1713 4.317460e-02
R8119 n2_6054_1713 n2_6054_1746 2.095238e-02
R8120 n2_6054_1746 n2_6054_1760 8.888889e-03
R8121 n2_6054_1760 n2_6054_1929 1.073016e-01
R8122 n2_6054_1929 n2_6054_1962 2.095238e-02
R8123 n2_6054_1962 n2_6054_2145 1.161905e-01
R8124 n2_6054_2145 n2_6054_2178 2.095238e-02
R8125 n2_6054_2178 n2_6054_2361 1.161905e-01
R8126 n2_6054_2361 n2_6054_2394 2.095238e-02
R8127 n2_6054_2394 n2_6054_2408 8.888889e-03
R8128 n2_6054_2408 n2_6054_2577 1.073016e-01
R8129 n2_6054_2577 n2_6054_2610 2.095238e-02
R8130 n2_6054_2610 n2_6054_2674 4.063492e-02
R8131 n2_6054_2674 n2_6054_2770 6.095238e-02
R8132 n2_6054_2770 n2_6054_2793 1.460317e-02
R8133 n2_6054_2793 n2_6054_2826 2.095238e-02
R8134 n2_6054_2826 n2_6054_2840 8.888889e-03
R8135 n2_6054_2840 n2_6054_3009 1.073016e-01
R8136 n2_6054_3009 n2_6054_3042 2.095238e-02
R8137 n2_6054_3042 n2_6054_3056 8.888889e-03
R8138 n2_6054_3056 n2_6054_3225 1.073016e-01
R8139 n2_6054_3225 n2_6054_3258 2.095238e-02
R8140 n2_6054_3258 n2_6054_3441 1.161905e-01
R8141 n2_6054_3441 n2_6054_3474 2.095238e-02
R8142 n2_6054_3474 n2_6054_3488 8.888889e-03
R8143 n2_6054_3488 n2_6054_3657 1.073016e-01
R8144 n2_6054_3657 n2_6054_3690 2.095238e-02
R8145 n2_6054_3690 n2_6054_3799 6.920635e-02
R8146 n2_6054_3799 n2_6054_3873 4.698413e-02
R8147 n2_6054_3873 n2_6054_3895 1.396825e-02
R8148 n2_6054_3895 n2_6054_3906 6.984127e-03
R8149 n2_6054_3906 n2_6054_4089 1.161905e-01
R8150 n2_6054_4089 n2_6054_4122 2.095238e-02
R8151 n2_6054_4122 n2_6054_4136 8.888889e-03
R8152 n2_6054_4136 n2_6054_4305 1.073016e-01
R8153 n2_6054_4305 n2_6054_4338 2.095238e-02
R8154 n2_6054_4338 n2_6054_4352 8.888889e-03
R8155 n2_6054_4352 n2_6054_4375 1.460317e-02
R8156 n2_6054_4375 n2_6054_4521 9.269841e-02
R8157 n2_6054_4521 n2_6054_4554 2.095238e-02
R8158 n2_6054_4554 n2_6054_4568 8.888889e-03
R8159 n2_6054_4568 n2_6054_4737 1.073016e-01
R8160 n2_6054_4737 n2_6054_4770 2.095238e-02
R8161 n2_6054_4770 n2_6054_4924 9.777778e-02
R8162 n2_6054_4924 n2_6054_4953 1.841270e-02
R8163 n2_6054_4953 n2_6054_4986 2.095238e-02
R8164 n2_6054_4986 n2_6054_5020 2.158730e-02
R8165 n2_6054_5020 n2_6054_5169 9.460317e-02
R8166 n2_6054_5169 n2_6054_5202 2.095238e-02
R8167 n2_6054_5202 n2_6054_5216 8.888889e-03
R8168 n2_6054_5216 n2_6054_5385 1.073016e-01
R8169 n2_6054_5385 n2_6054_5418 2.095238e-02
R8170 n2_6054_5418 n2_6054_5432 8.888889e-03
R8171 n2_6054_5432 n2_6054_5455 1.460317e-02
R8172 n2_6054_5455 n2_6054_5601 9.269841e-02
R8173 n2_6054_5601 n2_6054_5634 2.095238e-02
R8174 n2_6054_5634 n2_6054_5817 1.161905e-01
R8175 n2_6054_5817 n2_6054_5850 2.095238e-02
R8176 n2_6054_5850 n2_6054_6033 1.161905e-01
R8177 n2_6054_6033 n2_6054_6049 1.015873e-02
R8178 n2_6054_6049 n2_6054_6066 1.079365e-02
R8179 n2_6054_6066 n2_6054_6145 5.015873e-02
R8180 n2_6054_6145 n2_6054_6249 6.603175e-02
R8181 n2_6054_6249 n2_6054_6282 2.095238e-02
R8182 n2_6054_6282 n2_6054_6465 1.161905e-01
R8183 n2_6054_6465 n2_6054_6498 2.095238e-02
R8184 n2_6054_6498 n2_6054_6535 2.349206e-02
R8185 n2_6054_6535 n2_6054_6681 9.269841e-02
R8186 n2_6054_6681 n2_6054_6714 2.095238e-02
R8187 n2_6054_6714 n2_6054_6897 1.161905e-01
R8188 n2_6054_6897 n2_6054_6930 2.095238e-02
R8189 n2_6054_6930 n2_6054_7113 1.161905e-01
R8190 n2_6054_7329 n2_6054_7362 2.095238e-02
R8191 n2_6054_7362 n2_6054_7545 1.161905e-01
R8192 n2_6054_7545 n2_6054_7578 2.095238e-02
R8193 n2_6054_7578 n2_6054_7761 1.161905e-01
R8194 n2_6054_7761 n2_6054_7794 2.095238e-02
R8195 n2_6054_7794 n2_6054_7808 8.888889e-03
R8196 n2_6054_7808 n2_6054_7977 1.073016e-01
R8197 n2_6054_7977 n2_6054_8010 2.095238e-02
R8198 n2_6054_8010 n2_6054_8193 1.161905e-01
R8199 n2_6054_8193 n2_6054_8226 2.095238e-02
R8200 n2_6054_8226 n2_6054_8299 4.634921e-02
R8201 n2_6054_8299 n2_6054_8395 6.095238e-02
R8202 n2_6054_8395 n2_6054_8409 8.888889e-03
R8203 n2_6054_8409 n2_6054_8442 2.095238e-02
R8204 n2_6054_8442 n2_6054_8625 1.161905e-01
R8205 n2_6054_8625 n2_6054_8658 2.095238e-02
R8206 n2_6054_8658 n2_6054_8841 1.161905e-01
R8207 n2_6054_8841 n2_6054_8874 2.095238e-02
R8208 n2_6054_8874 n2_6054_8888 8.888889e-03
R8209 n2_6054_8888 n2_6054_8911 1.460317e-02
R8210 n2_6054_8911 n2_6054_9057 9.269841e-02
R8211 n2_6054_9057 n2_6054_9090 2.095238e-02
R8212 n2_6054_9090 n2_6054_9273 1.161905e-01
R8213 n2_6054_9273 n2_6054_9306 2.095238e-02
R8214 n2_6054_9705 n2_6054_9738 2.095238e-02
R8215 n2_6054_9738 n2_6054_9921 1.161905e-01
R8216 n2_6054_9921 n2_6054_9954 2.095238e-02
R8217 n2_6054_9954 n2_6054_9968 8.888889e-03
R8218 n2_6054_9968 n2_6054_10137 1.073016e-01
R8219 n2_6054_10137 n2_6054_10170 2.095238e-02
R8220 n2_6054_10170 n2_6054_10353 1.161905e-01
R8221 n2_6054_10353 n2_6054_10386 2.095238e-02
R8222 n2_6054_10386 n2_6054_10549 1.034921e-01
R8223 n2_6054_10549 n2_6054_10569 1.269841e-02
R8224 n2_6054_10569 n2_6054_10602 2.095238e-02
R8225 n2_6054_10602 n2_6054_10645 2.730159e-02
R8226 n2_6054_10645 n2_6054_10785 8.888889e-02
R8227 n2_6054_10785 n2_6054_10818 2.095238e-02
R8228 n2_6054_10818 n2_6054_11001 1.161905e-01
R8229 n2_6054_11001 n2_6054_11034 2.095238e-02
R8230 n2_6054_11034 n2_6054_11048 8.888889e-03
R8231 n2_6054_11048 n2_6054_11071 1.460317e-02
R8232 n2_6054_11071 n2_6054_11217 9.269841e-02
R8233 n2_6054_11217 n2_6054_11250 2.095238e-02
R8234 n2_6054_11250 n2_6054_11433 1.161905e-01
R8235 n2_6054_11433 n2_6054_11466 2.095238e-02
R8236 n2_6054_11865 n2_6054_11898 2.095238e-02
R8237 n2_6054_11898 n2_6054_12081 1.161905e-01
R8238 n2_6054_12081 n2_6054_12114 2.095238e-02
R8239 n2_6054_12114 n2_6054_12128 8.888889e-03
R8240 n2_6054_12128 n2_6054_12297 1.073016e-01
R8241 n2_6054_12297 n2_6054_12330 2.095238e-02
R8242 n2_6054_12330 n2_6054_12513 1.161905e-01
R8243 n2_6054_12513 n2_6054_12546 2.095238e-02
R8244 n2_6054_12546 n2_6054_12729 1.161905e-01
R8245 n2_6054_12729 n2_6054_12762 2.095238e-02
R8246 n2_6054_12762 n2_6054_12799 2.349206e-02
R8247 n2_6054_12799 n2_6054_12895 6.095238e-02
R8248 n2_6054_12895 n2_6054_12945 3.174603e-02
R8249 n2_6054_12945 n2_6054_12978 2.095238e-02
R8250 n2_6054_12978 n2_6054_13161 1.161905e-01
R8251 n2_6054_13161 n2_6054_13194 2.095238e-02
R8252 n2_6054_13194 n2_6054_13377 1.161905e-01
R8253 n2_6054_13377 n2_6054_13410 2.095238e-02
R8254 n2_6054_13410 n2_6054_13424 8.888889e-03
R8255 n2_6054_13424 n2_6054_13593 1.073016e-01
R8256 n2_6054_13593 n2_6054_13626 2.095238e-02
R8257 n2_6054_13626 n2_6054_13809 1.161905e-01
R8258 n2_6054_13809 n2_6054_13842 2.095238e-02
R8259 n2_6054_14241 n2_6054_14274 2.095238e-02
R8260 n2_6054_14274 n2_6054_14457 1.161905e-01
R8261 n2_6054_14457 n2_6054_14490 2.095238e-02
R8262 n2_6054_14490 n2_6054_14536 2.920635e-02
R8263 n2_6054_14536 n2_6054_14673 8.698413e-02
R8264 n2_6054_14673 n2_6054_14706 2.095238e-02
R8265 n2_6054_14706 n2_6054_14889 1.161905e-01
R8266 n2_6054_14889 n2_6054_14922 2.095238e-02
R8267 n2_6054_14922 n2_6054_15049 8.063492e-02
R8268 n2_6054_15049 n2_6054_15105 3.555556e-02
R8269 n2_6054_15105 n2_6054_15138 2.095238e-02
R8270 n2_6054_15138 n2_6054_15145 4.444444e-03
R8271 n2_6054_15145 n2_6054_15321 1.117460e-01
R8272 n2_6054_15321 n2_6054_15354 2.095238e-02
R8273 n2_6054_15354 n2_6054_15537 1.161905e-01
R8274 n2_6054_15537 n2_6054_15570 2.095238e-02
R8275 n2_6054_15570 n2_6054_15584 8.888889e-03
R8276 n2_6054_15584 n2_6054_15753 1.073016e-01
R8277 n2_6054_15753 n2_6054_15786 2.095238e-02
R8278 n2_6054_15786 n2_6054_15800 8.888889e-03
R8279 n2_6054_15800 n2_6054_15969 1.073016e-01
R8280 n2_6054_15969 n2_6054_16002 2.095238e-02
R8281 n2_6054_16002 n2_6054_16016 8.888889e-03
R8282 n2_6054_16016 n2_6054_16174 1.003175e-01
R8283 n2_6054_16174 n2_6054_16185 6.984127e-03
R8284 n2_6054_16185 n2_6054_16218 2.095238e-02
R8285 n2_6054_16218 n2_6054_16270 3.301587e-02
R8286 n2_6054_16270 n2_6054_16401 8.317460e-02
R8287 n2_6054_16401 n2_6054_16434 2.095238e-02
R8288 n2_6054_16434 n2_6054_16617 1.161905e-01
R8289 n2_6054_16617 n2_6054_16650 2.095238e-02
R8290 n2_6054_16650 n2_6054_16833 1.161905e-01
R8291 n2_6054_16833 n2_6054_16866 2.095238e-02
R8292 n2_6054_16866 n2_6054_17049 1.161905e-01
R8293 n2_6054_17049 n2_6054_17082 2.095238e-02
R8294 n2_6054_17082 n2_6054_17096 8.888889e-03
R8295 n2_6054_17096 n2_6054_17119 1.460317e-02
R8296 n2_6054_17119 n2_6054_17265 9.269841e-02
R8297 n2_6054_17265 n2_6054_17298 2.095238e-02
R8298 n2_6054_17298 n2_6054_17299 6.349206e-04
R8299 n2_6054_17299 n2_6054_17312 8.253968e-03
R8300 n2_6054_17312 n2_6054_17335 1.460317e-02
R8301 n2_6054_17335 n2_6054_17395 3.809524e-02
R8302 n2_6054_17395 n2_6054_17481 5.460317e-02
R8303 n2_6054_17481 n2_6054_17514 2.095238e-02
R8304 n2_6054_17514 n2_6054_17528 8.888889e-03
R8305 n2_6054_17528 n2_6054_17697 1.073016e-01
R8306 n2_6054_17697 n2_6054_17730 2.095238e-02
R8307 n2_6054_17730 n2_6054_17913 1.161905e-01
R8308 n2_6054_17913 n2_6054_17946 2.095238e-02
R8309 n2_6054_17946 n2_6054_18129 1.161905e-01
R8310 n2_6054_18129 n2_6054_18162 2.095238e-02
R8311 n2_6054_18162 n2_6054_18345 1.161905e-01
R8312 n2_6054_18345 n2_6054_18378 2.095238e-02
R8313 n2_6054_18378 n2_6054_18392 8.888889e-03
R8314 n2_6054_18392 n2_6054_18424 2.031746e-02
R8315 n2_6054_18424 n2_6054_18520 6.095238e-02
R8316 n2_6054_18520 n2_6054_18561 2.603175e-02
R8317 n2_6054_18561 n2_6054_18594 2.095238e-02
R8318 n2_6054_18594 n2_6054_18608 8.888889e-03
R8319 n2_6054_18608 n2_6054_18777 1.073016e-01
R8320 n2_6054_18777 n2_6054_18810 2.095238e-02
R8321 n2_6054_18810 n2_6054_18824 8.888889e-03
R8322 n2_6054_18824 n2_6054_18993 1.073016e-01
R8323 n2_6054_18993 n2_6054_19026 2.095238e-02
R8324 n2_6054_19026 n2_6054_19040 8.888889e-03
R8325 n2_6054_19040 n2_6054_19209 1.073016e-01
R8326 n2_6054_19209 n2_6054_19242 2.095238e-02
R8327 n2_6054_19242 n2_6054_19425 1.161905e-01
R8328 n2_6054_19425 n2_6054_19458 2.095238e-02
R8329 n2_6054_19458 n2_6054_19472 8.888889e-03
R8330 n2_6054_19472 n2_6054_19549 4.888889e-02
R8331 n2_6054_19549 n2_6054_19641 5.841270e-02
R8332 n2_6054_19641 n2_6054_19645 2.539683e-03
R8333 n2_6054_19645 n2_6054_19674 1.841270e-02
R8334 n2_6054_19674 n2_6054_19857 1.161905e-01
R8335 n2_6054_19857 n2_6054_19890 2.095238e-02
R8336 n2_6054_19890 n2_6054_20073 1.161905e-01
R8337 n2_6054_20073 n2_6054_20106 2.095238e-02
R8338 n2_6054_20106 n2_6054_20289 1.161905e-01
R8339 n2_6054_20289 n2_6054_20322 2.095238e-02
R8340 n2_6054_20322 n2_6054_20505 1.161905e-01
R8341 n2_6054_20505 n2_6054_20538 2.095238e-02
R8342 n2_6054_20538 n2_6054_20674 8.634921e-02
R8343 n2_6054_20674 n2_6054_20721 2.984127e-02
R8344 n2_6054_20721 n2_6054_20754 2.095238e-02
R8345 n2_6054_20754 n2_6054_20770 1.015873e-02
R8346 n2_6054_20770 n2_6054_20937 1.060317e-01
R8347 n2_6054_20937 n2_6054_20970 2.095238e-02
R8348 n2_6146_201 n2_6146_234 2.095238e-02
R8349 n2_6146_234 n2_6146_356 7.746032e-02
R8350 n2_6146_356 n2_6146_417 3.873016e-02
R8351 n2_6146_417 n2_6146_424 4.444444e-03
R8352 n2_6146_424 n2_6146_450 1.650794e-02
R8353 n2_6146_520 n2_6146_633 7.174603e-02
R8354 n2_6146_633 n2_6146_666 2.095238e-02
R8355 n2_6146_666 n2_6146_788 7.746032e-02
R8356 n2_6146_788 n2_6146_849 3.873016e-02
R8357 n2_6146_849 n2_6146_882 2.095238e-02
R8358 n2_6146_882 n2_6146_1065 1.161905e-01
R8359 n2_6146_1065 n2_6146_1098 2.095238e-02
R8360 n2_6146_1098 n2_6146_1281 1.161905e-01
R8361 n2_6146_1281 n2_6146_1314 2.095238e-02
R8362 n2_6146_1314 n2_6146_1497 1.161905e-01
R8363 n2_6146_1497 n2_6146_1530 2.095238e-02
R8364 n2_6146_1530 n2_6146_1549 1.206349e-02
R8365 n2_6146_1645 n2_6146_1713 4.317460e-02
R8366 n2_6146_1713 n2_6146_1746 2.095238e-02
R8367 n2_6146_1746 n2_6146_1760 8.888889e-03
R8368 n2_6146_1760 n2_6146_1929 1.073016e-01
R8369 n2_6146_1929 n2_6146_1962 2.095238e-02
R8370 n2_6146_1962 n2_6146_2145 1.161905e-01
R8371 n2_6146_2145 n2_6146_2178 2.095238e-02
R8372 n2_6146_2178 n2_6146_2361 1.161905e-01
R8373 n2_6146_2361 n2_6146_2394 2.095238e-02
R8374 n2_6146_2394 n2_6146_2408 8.888889e-03
R8375 n2_6146_2408 n2_6146_2577 1.073016e-01
R8376 n2_6146_2577 n2_6146_2610 2.095238e-02
R8377 n2_6146_2610 n2_6146_2674 4.063492e-02
R8378 n2_6146_2770 n2_6146_2793 1.460317e-02
R8379 n2_6146_2793 n2_6146_2826 2.095238e-02
R8380 n2_6146_2826 n2_6146_2840 8.888889e-03
R8381 n2_6146_2840 n2_6146_3009 1.073016e-01
R8382 n2_6146_3009 n2_6146_3042 2.095238e-02
R8383 n2_6146_3042 n2_6146_3056 8.888889e-03
R8384 n2_6146_3056 n2_6146_3225 1.073016e-01
R8385 n2_6146_3225 n2_6146_3258 2.095238e-02
R8386 n2_6146_3258 n2_6146_3441 1.161905e-01
R8387 n2_6146_3441 n2_6146_3474 2.095238e-02
R8388 n2_6146_3474 n2_6146_3488 8.888889e-03
R8389 n2_6146_3488 n2_6146_3657 1.073016e-01
R8390 n2_6146_3657 n2_6146_3690 2.095238e-02
R8391 n2_6146_3690 n2_6146_3799 6.920635e-02
R8392 n2_6146_3873 n2_6146_3895 1.396825e-02
R8393 n2_6146_3895 n2_6146_3906 6.984127e-03
R8394 n2_6146_3906 n2_6146_4089 1.161905e-01
R8395 n2_6146_4089 n2_6146_4122 2.095238e-02
R8396 n2_6146_4122 n2_6146_4136 8.888889e-03
R8397 n2_6146_4136 n2_6146_4305 1.073016e-01
R8398 n2_6146_4305 n2_6146_4338 2.095238e-02
R8399 n2_6146_4338 n2_6146_4352 8.888889e-03
R8400 n2_6146_4352 n2_6146_4375 1.460317e-02
R8401 n2_6146_4375 n2_6146_4521 9.269841e-02
R8402 n2_6146_4521 n2_6146_4554 2.095238e-02
R8403 n2_6146_4554 n2_6146_4568 8.888889e-03
R8404 n2_6146_4568 n2_6146_4737 1.073016e-01
R8405 n2_6146_4737 n2_6146_4770 2.095238e-02
R8406 n2_6146_4770 n2_6146_4924 9.777778e-02
R8407 n2_6146_4924 n2_6146_4953 1.841270e-02
R8408 n2_6146_5020 n2_6146_5169 9.460317e-02
R8409 n2_6146_5169 n2_6146_5202 2.095238e-02
R8410 n2_6146_5202 n2_6146_5216 8.888889e-03
R8411 n2_6146_5216 n2_6146_5385 1.073016e-01
R8412 n2_6146_5385 n2_6146_5418 2.095238e-02
R8413 n2_6146_5418 n2_6146_5432 8.888889e-03
R8414 n2_6146_5432 n2_6146_5455 1.460317e-02
R8415 n2_6146_5455 n2_6146_5601 9.269841e-02
R8416 n2_6146_5601 n2_6146_5634 2.095238e-02
R8417 n2_6146_5634 n2_6146_5817 1.161905e-01
R8418 n2_6146_5817 n2_6146_5850 2.095238e-02
R8419 n2_6146_5850 n2_6146_6033 1.161905e-01
R8420 n2_6146_6033 n2_6146_6049 1.015873e-02
R8421 n2_6146_6049 n2_6146_6066 1.079365e-02
R8422 n2_6146_15138 n2_6146_15145 4.444444e-03
R8423 n2_6146_15145 n2_6146_15321 1.117460e-01
R8424 n2_6146_15321 n2_6146_15354 2.095238e-02
R8425 n2_6146_15354 n2_6146_15537 1.161905e-01
R8426 n2_6146_15537 n2_6146_15570 2.095238e-02
R8427 n2_6146_15570 n2_6146_15584 8.888889e-03
R8428 n2_6146_15584 n2_6146_15753 1.073016e-01
R8429 n2_6146_15753 n2_6146_15786 2.095238e-02
R8430 n2_6146_15786 n2_6146_15800 8.888889e-03
R8431 n2_6146_15800 n2_6146_15969 1.073016e-01
R8432 n2_6146_15969 n2_6146_16002 2.095238e-02
R8433 n2_6146_16002 n2_6146_16016 8.888889e-03
R8434 n2_6146_16016 n2_6146_16174 1.003175e-01
R8435 n2_6146_16174 n2_6146_16185 6.984127e-03
R8436 n2_6146_16270 n2_6146_16401 8.317460e-02
R8437 n2_6146_16401 n2_6146_16434 2.095238e-02
R8438 n2_6146_16434 n2_6146_16617 1.161905e-01
R8439 n2_6146_16617 n2_6146_16650 2.095238e-02
R8440 n2_6146_16650 n2_6146_16833 1.161905e-01
R8441 n2_6146_16833 n2_6146_16866 2.095238e-02
R8442 n2_6146_16866 n2_6146_17049 1.161905e-01
R8443 n2_6146_17049 n2_6146_17082 2.095238e-02
R8444 n2_6146_17082 n2_6146_17096 8.888889e-03
R8445 n2_6146_17096 n2_6146_17119 1.460317e-02
R8446 n2_6146_17119 n2_6146_17265 9.269841e-02
R8447 n2_6146_17265 n2_6146_17298 2.095238e-02
R8448 n2_6146_17298 n2_6146_17299 6.349206e-04
R8449 n2_6146_17299 n2_6146_17312 8.253968e-03
R8450 n2_6146_17395 n2_6146_17481 5.460317e-02
R8451 n2_6146_17481 n2_6146_17514 2.095238e-02
R8452 n2_6146_17514 n2_6146_17528 8.888889e-03
R8453 n2_6146_17528 n2_6146_17697 1.073016e-01
R8454 n2_6146_17697 n2_6146_17730 2.095238e-02
R8455 n2_6146_17730 n2_6146_17913 1.161905e-01
R8456 n2_6146_17913 n2_6146_17946 2.095238e-02
R8457 n2_6146_17946 n2_6146_18129 1.161905e-01
R8458 n2_6146_18129 n2_6146_18162 2.095238e-02
R8459 n2_6146_18162 n2_6146_18345 1.161905e-01
R8460 n2_6146_18345 n2_6146_18378 2.095238e-02
R8461 n2_6146_18378 n2_6146_18392 8.888889e-03
R8462 n2_6146_18392 n2_6146_18424 2.031746e-02
R8463 n2_6146_18520 n2_6146_18561 2.603175e-02
R8464 n2_6146_18561 n2_6146_18594 2.095238e-02
R8465 n2_6146_18594 n2_6146_18608 8.888889e-03
R8466 n2_6146_18608 n2_6146_18777 1.073016e-01
R8467 n2_6146_18777 n2_6146_18810 2.095238e-02
R8468 n2_6146_18810 n2_6146_18824 8.888889e-03
R8469 n2_6146_18824 n2_6146_18993 1.073016e-01
R8470 n2_6146_18993 n2_6146_19026 2.095238e-02
R8471 n2_6146_19026 n2_6146_19040 8.888889e-03
R8472 n2_6146_19040 n2_6146_19209 1.073016e-01
R8473 n2_6146_19209 n2_6146_19242 2.095238e-02
R8474 n2_6146_19242 n2_6146_19425 1.161905e-01
R8475 n2_6146_19425 n2_6146_19458 2.095238e-02
R8476 n2_6146_19458 n2_6146_19472 8.888889e-03
R8477 n2_6146_19472 n2_6146_19549 4.888889e-02
R8478 n2_6146_19641 n2_6146_19645 2.539683e-03
R8479 n2_6146_19645 n2_6146_19674 1.841270e-02
R8480 n2_6146_19674 n2_6146_19857 1.161905e-01
R8481 n2_6146_19857 n2_6146_19890 2.095238e-02
R8482 n2_6146_19890 n2_6146_20073 1.161905e-01
R8483 n2_6146_20073 n2_6146_20106 2.095238e-02
R8484 n2_6146_20106 n2_6146_20289 1.161905e-01
R8485 n2_6146_20289 n2_6146_20322 2.095238e-02
R8486 n2_6146_20322 n2_6146_20505 1.161905e-01
R8487 n2_6146_20505 n2_6146_20538 2.095238e-02
R8488 n2_6146_20538 n2_6146_20674 8.634921e-02
R8489 n2_6146_20754 n2_6146_20770 1.015873e-02
R8490 n2_6146_20770 n2_6146_20937 1.060317e-01
R8491 n2_6146_20937 n2_6146_20970 2.095238e-02
R8492 n2_6991_7329 n2_6991_7362 2.095238e-02
R8493 n2_6991_7362 n2_6991_7545 1.161905e-01
R8494 n2_6991_7545 n2_6991_7578 2.095238e-02
R8495 n2_6991_7578 n2_6991_7761 1.161905e-01
R8496 n2_6991_7761 n2_6991_7794 2.095238e-02
R8497 n2_6991_7794 n2_6991_7808 8.888889e-03
R8498 n2_6991_7808 n2_6991_7977 1.073016e-01
R8499 n2_6991_7977 n2_6991_8010 2.095238e-02
R8500 n2_6991_8010 n2_6991_8193 1.161905e-01
R8501 n2_6991_8193 n2_6991_8226 2.095238e-02
R8502 n2_6991_8226 n2_6991_8299 4.634921e-02
R8503 n2_6991_8395 n2_6991_8409 8.888889e-03
R8504 n2_6991_8409 n2_6991_8442 2.095238e-02
R8505 n2_6991_8442 n2_6991_8625 1.161905e-01
R8506 n2_6991_8625 n2_6991_8658 2.095238e-02
R8507 n2_6991_8658 n2_6991_8841 1.161905e-01
R8508 n2_6991_8841 n2_6991_8874 2.095238e-02
R8509 n2_6991_8874 n2_6991_8888 8.888889e-03
R8510 n2_6991_8888 n2_6991_9057 1.073016e-01
R8511 n2_6991_9057 n2_6991_9090 2.095238e-02
R8512 n2_6991_9090 n2_6991_9273 1.161905e-01
R8513 n2_6991_9273 n2_6991_9306 2.095238e-02
R8514 n2_6991_9306 n2_6991_9489 1.161905e-01
R8515 n2_6991_9489 n2_6991_9522 2.095238e-02
R8516 n2_6991_9522 n2_6991_9705 1.161905e-01
R8517 n2_6991_9705 n2_6991_9738 2.095238e-02
R8518 n2_6991_9738 n2_6991_9921 1.161905e-01
R8519 n2_6991_9921 n2_6991_9954 2.095238e-02
R8520 n2_6991_9954 n2_6991_9968 8.888889e-03
R8521 n2_6991_9968 n2_6991_10137 1.073016e-01
R8522 n2_6991_10137 n2_6991_10170 2.095238e-02
R8523 n2_6991_10170 n2_6991_10353 1.161905e-01
R8524 n2_6991_10353 n2_6991_10386 2.095238e-02
R8525 n2_6991_10386 n2_6991_10549 1.034921e-01
R8526 n2_6991_10549 n2_6991_10569 1.269841e-02
R8527 n2_6991_10645 n2_6991_10785 8.888889e-02
R8528 n2_6991_10785 n2_6991_10818 2.095238e-02
R8529 n2_6991_10818 n2_6991_11001 1.161905e-01
R8530 n2_6991_11001 n2_6991_11034 2.095238e-02
R8531 n2_6991_11034 n2_6991_11048 8.888889e-03
R8532 n2_6991_11048 n2_6991_11217 1.073016e-01
R8533 n2_6991_11217 n2_6991_11250 2.095238e-02
R8534 n2_6991_11250 n2_6991_11433 1.161905e-01
R8535 n2_6991_11433 n2_6991_11466 2.095238e-02
R8536 n2_6991_11466 n2_6991_11649 1.161905e-01
R8537 n2_6991_11649 n2_6991_11682 2.095238e-02
R8538 n2_6991_11682 n2_6991_11865 1.161905e-01
R8539 n2_6991_11865 n2_6991_11898 2.095238e-02
R8540 n2_6991_11898 n2_6991_12081 1.161905e-01
R8541 n2_6991_12081 n2_6991_12114 2.095238e-02
R8542 n2_6991_12114 n2_6991_12128 8.888889e-03
R8543 n2_6991_12128 n2_6991_12297 1.073016e-01
R8544 n2_6991_12297 n2_6991_12330 2.095238e-02
R8545 n2_6991_12330 n2_6991_12513 1.161905e-01
R8546 n2_6991_12513 n2_6991_12546 2.095238e-02
R8547 n2_6991_12546 n2_6991_12729 1.161905e-01
R8548 n2_6991_12729 n2_6991_12762 2.095238e-02
R8549 n2_6991_12762 n2_6991_12799 2.349206e-02
R8550 n2_6991_12895 n2_6991_12945 3.174603e-02
R8551 n2_6991_12945 n2_6991_12978 2.095238e-02
R8552 n2_6991_12978 n2_6991_13161 1.161905e-01
R8553 n2_6991_13161 n2_6991_13194 2.095238e-02
R8554 n2_6991_13194 n2_6991_13377 1.161905e-01
R8555 n2_6991_13377 n2_6991_13410 2.095238e-02
R8556 n2_6991_13410 n2_6991_13424 8.888889e-03
R8557 n2_6991_13424 n2_6991_13593 1.073016e-01
R8558 n2_6991_13593 n2_6991_13626 2.095238e-02
R8559 n2_6991_13626 n2_6991_13809 1.161905e-01
R8560 n2_6991_13809 n2_6991_13842 2.095238e-02
R8561 n2_6991_8299 n2_7130_8299 8.825397e-02
R8562 n2_7130_8299 n2_7179_8299 3.111111e-02
R8563 n2_6991_8395 n2_7130_8395 8.825397e-02
R8564 n2_7130_8395 n2_7179_8395 3.111111e-02
R8565 n2_6991_10549 n2_7130_10549 8.825397e-02
R8566 n2_7130_10549 n2_7179_10549 3.111111e-02
R8567 n2_6991_10645 n2_7130_10645 8.825397e-02
R8568 n2_7130_10645 n2_7179_10645 3.111111e-02
R8569 n2_6991_12799 n2_7130_12799 8.825397e-02
R8570 n2_7130_12799 n2_7179_12799 3.111111e-02
R8571 n2_6991_12895 n2_7130_12895 8.825397e-02
R8572 n2_7130_12895 n2_7179_12895 3.111111e-02
R8573 n2_7179_7329 n2_7179_7362 2.095238e-02
R8574 n2_7179_7362 n2_7179_7545 1.161905e-01
R8575 n2_7179_7545 n2_7179_7578 2.095238e-02
R8576 n2_7179_7578 n2_7179_7761 1.161905e-01
R8577 n2_7179_7761 n2_7179_7794 2.095238e-02
R8578 n2_7179_7794 n2_7179_7808 8.888889e-03
R8579 n2_7179_7808 n2_7179_7977 1.073016e-01
R8580 n2_7179_7977 n2_7179_8010 2.095238e-02
R8581 n2_7179_8010 n2_7179_8193 1.161905e-01
R8582 n2_7179_8193 n2_7179_8226 2.095238e-02
R8583 n2_7179_8226 n2_7179_8299 4.634921e-02
R8584 n2_7179_8299 n2_7179_8395 6.095238e-02
R8585 n2_7179_8395 n2_7179_8409 8.888889e-03
R8586 n2_7179_8409 n2_7179_8442 2.095238e-02
R8587 n2_7179_8442 n2_7179_8625 1.161905e-01
R8588 n2_7179_8625 n2_7179_8658 2.095238e-02
R8589 n2_7179_8658 n2_7179_8841 1.161905e-01
R8590 n2_7179_8841 n2_7179_8874 2.095238e-02
R8591 n2_7179_8874 n2_7179_8888 8.888889e-03
R8592 n2_7179_8888 n2_7179_9057 1.073016e-01
R8593 n2_7179_9057 n2_7179_9090 2.095238e-02
R8594 n2_7179_9090 n2_7179_9273 1.161905e-01
R8595 n2_7179_9273 n2_7179_9306 2.095238e-02
R8596 n2_7179_9705 n2_7179_9738 2.095238e-02
R8597 n2_7179_9738 n2_7179_9921 1.161905e-01
R8598 n2_7179_9921 n2_7179_9954 2.095238e-02
R8599 n2_7179_9954 n2_7179_9968 8.888889e-03
R8600 n2_7179_9968 n2_7179_10137 1.073016e-01
R8601 n2_7179_10137 n2_7179_10170 2.095238e-02
R8602 n2_7179_10170 n2_7179_10353 1.161905e-01
R8603 n2_7179_10353 n2_7179_10386 2.095238e-02
R8604 n2_7179_10386 n2_7179_10549 1.034921e-01
R8605 n2_7179_10549 n2_7179_10569 1.269841e-02
R8606 n2_7179_10569 n2_7179_10602 2.095238e-02
R8607 n2_7179_10602 n2_7179_10645 2.730159e-02
R8608 n2_7179_10645 n2_7179_10785 8.888889e-02
R8609 n2_7179_10785 n2_7179_10818 2.095238e-02
R8610 n2_7179_10818 n2_7179_11001 1.161905e-01
R8611 n2_7179_11001 n2_7179_11034 2.095238e-02
R8612 n2_7179_11034 n2_7179_11048 8.888889e-03
R8613 n2_7179_11048 n2_7179_11217 1.073016e-01
R8614 n2_7179_11217 n2_7179_11250 2.095238e-02
R8615 n2_7179_11250 n2_7179_11433 1.161905e-01
R8616 n2_7179_11433 n2_7179_11466 2.095238e-02
R8617 n2_7179_11865 n2_7179_11898 2.095238e-02
R8618 n2_7179_11898 n2_7179_12081 1.161905e-01
R8619 n2_7179_12081 n2_7179_12114 2.095238e-02
R8620 n2_7179_12114 n2_7179_12128 8.888889e-03
R8621 n2_7179_12128 n2_7179_12297 1.073016e-01
R8622 n2_7179_12297 n2_7179_12330 2.095238e-02
R8623 n2_7179_12330 n2_7179_12513 1.161905e-01
R8624 n2_7179_12513 n2_7179_12546 2.095238e-02
R8625 n2_7179_12546 n2_7179_12729 1.161905e-01
R8626 n2_7179_12729 n2_7179_12762 2.095238e-02
R8627 n2_7179_12762 n2_7179_12799 2.349206e-02
R8628 n2_7179_12799 n2_7179_12895 6.095238e-02
R8629 n2_7179_12895 n2_7179_12945 3.174603e-02
R8630 n2_7179_12945 n2_7179_12978 2.095238e-02
R8631 n2_7179_12978 n2_7179_13161 1.161905e-01
R8632 n2_7179_13161 n2_7179_13194 2.095238e-02
R8633 n2_7179_13194 n2_7179_13377 1.161905e-01
R8634 n2_7179_13377 n2_7179_13410 2.095238e-02
R8635 n2_7179_13410 n2_7179_13424 8.888889e-03
R8636 n2_7179_13424 n2_7179_13593 1.073016e-01
R8637 n2_7179_13593 n2_7179_13626 2.095238e-02
R8638 n2_7179_13626 n2_7179_13809 1.161905e-01
R8639 n2_7179_13809 n2_7179_13842 2.095238e-02
R8640 n2_8116_201 n2_8116_234 2.095238e-02
R8641 n2_8116_234 n2_8116_417 1.161905e-01
R8642 n2_8116_417 n2_8116_424 4.444444e-03
R8643 n2_8116_424 n2_8116_450 1.650794e-02
R8644 n2_8116_520 n2_8116_633 7.174603e-02
R8645 n2_8116_633 n2_8116_666 2.095238e-02
R8646 n2_8116_666 n2_8116_849 1.161905e-01
R8647 n2_8116_849 n2_8116_882 2.095238e-02
R8648 n2_8116_882 n2_8116_1065 1.161905e-01
R8649 n2_8116_1065 n2_8116_1098 2.095238e-02
R8650 n2_8116_1098 n2_8116_1281 1.161905e-01
R8651 n2_8116_1281 n2_8116_1314 2.095238e-02
R8652 n2_8116_1314 n2_8116_1497 1.161905e-01
R8653 n2_8116_1497 n2_8116_1530 2.095238e-02
R8654 n2_8116_1530 n2_8116_1549 1.206349e-02
R8655 n2_8116_1645 n2_8116_1713 4.317460e-02
R8656 n2_8116_1713 n2_8116_1746 2.095238e-02
R8657 n2_8116_1746 n2_8116_1760 8.888889e-03
R8658 n2_8116_1760 n2_8116_1783 1.460317e-02
R8659 n2_8116_1783 n2_8116_1929 9.269841e-02
R8660 n2_8116_1929 n2_8116_1962 2.095238e-02
R8661 n2_8116_1962 n2_8116_2145 1.161905e-01
R8662 n2_8116_2145 n2_8116_2178 2.095238e-02
R8663 n2_8116_2178 n2_8116_2361 1.161905e-01
R8664 n2_8116_2361 n2_8116_2394 2.095238e-02
R8665 n2_8116_2394 n2_8116_2408 8.888889e-03
R8666 n2_8116_2408 n2_8116_2577 1.073016e-01
R8667 n2_8116_2577 n2_8116_2610 2.095238e-02
R8668 n2_8116_2610 n2_8116_2674 4.063492e-02
R8669 n2_8116_2770 n2_8116_2793 1.460317e-02
R8670 n2_8116_2793 n2_8116_2826 2.095238e-02
R8671 n2_8116_2826 n2_8116_2840 8.888889e-03
R8672 n2_8116_2840 n2_8116_2863 1.460317e-02
R8673 n2_8116_2863 n2_8116_3009 9.269841e-02
R8674 n2_8116_3009 n2_8116_3042 2.095238e-02
R8675 n2_8116_3042 n2_8116_3225 1.161905e-01
R8676 n2_8116_3225 n2_8116_3258 2.095238e-02
R8677 n2_8116_3258 n2_8116_3441 1.161905e-01
R8678 n2_8116_3441 n2_8116_3474 2.095238e-02
R8679 n2_8116_3474 n2_8116_3488 8.888889e-03
R8680 n2_8116_3488 n2_8116_3657 1.073016e-01
R8681 n2_8116_3657 n2_8116_3690 2.095238e-02
R8682 n2_8116_3690 n2_8116_3799 6.920635e-02
R8683 n2_8116_3873 n2_8116_3895 1.396825e-02
R8684 n2_8116_3895 n2_8116_3906 6.984127e-03
R8685 n2_8116_3906 n2_8116_4089 1.161905e-01
R8686 n2_8116_4089 n2_8116_4122 2.095238e-02
R8687 n2_8116_4122 n2_8116_4136 8.888889e-03
R8688 n2_8116_4136 n2_8116_4305 1.073016e-01
R8689 n2_8116_4305 n2_8116_4338 2.095238e-02
R8690 n2_8116_4338 n2_8116_4521 1.161905e-01
R8691 n2_8116_4521 n2_8116_4554 2.095238e-02
R8692 n2_8116_4554 n2_8116_4568 8.888889e-03
R8693 n2_8116_4568 n2_8116_4737 1.073016e-01
R8694 n2_8116_4737 n2_8116_4770 2.095238e-02
R8695 n2_8116_4770 n2_8116_4924 9.777778e-02
R8696 n2_8116_4924 n2_8116_4953 1.841270e-02
R8697 n2_8116_5020 n2_8116_5169 9.460317e-02
R8698 n2_8116_5169 n2_8116_5202 2.095238e-02
R8699 n2_8116_5202 n2_8116_5216 8.888889e-03
R8700 n2_8116_5216 n2_8116_5239 1.460317e-02
R8701 n2_8116_5239 n2_8116_5385 9.269841e-02
R8702 n2_8116_5385 n2_8116_5418 2.095238e-02
R8703 n2_8116_5418 n2_8116_5432 8.888889e-03
R8704 n2_8116_5432 n2_8116_5455 1.460317e-02
R8705 n2_8116_5455 n2_8116_5601 9.269841e-02
R8706 n2_8116_5601 n2_8116_5634 2.095238e-02
R8707 n2_8116_5634 n2_8116_5817 1.161905e-01
R8708 n2_8116_5817 n2_8116_5850 2.095238e-02
R8709 n2_8116_5850 n2_8116_6033 1.161905e-01
R8710 n2_8116_6033 n2_8116_6049 1.015873e-02
R8711 n2_8116_6049 n2_8116_6066 1.079365e-02
R8712 n2_8116_6145 n2_8116_6249 6.603175e-02
R8713 n2_8116_6249 n2_8116_6282 2.095238e-02
R8714 n2_8116_6282 n2_8116_6465 1.161905e-01
R8715 n2_8116_6465 n2_8116_6498 2.095238e-02
R8716 n2_8116_6498 n2_8116_6512 8.888889e-03
R8717 n2_8116_6512 n2_8116_6535 1.460317e-02
R8718 n2_8116_6535 n2_8116_6681 9.269841e-02
R8719 n2_8116_6681 n2_8116_6714 2.095238e-02
R8720 n2_8116_6714 n2_8116_6897 1.161905e-01
R8721 n2_8116_6897 n2_8116_6930 2.095238e-02
R8722 n2_8116_6930 n2_8116_6944 8.888889e-03
R8723 n2_8116_6944 n2_8116_7113 1.073016e-01
R8724 n2_8116_7113 n2_8116_7146 2.095238e-02
R8725 n2_8116_7146 n2_8116_7160 8.888889e-03
R8726 n2_8116_7160 n2_8116_7174 8.888889e-03
R8727 n2_8116_7270 n2_8116_7329 3.746032e-02
R8728 n2_8116_7329 n2_8116_7362 2.095238e-02
R8729 n2_8116_7362 n2_8116_7376 8.888889e-03
R8730 n2_8116_7376 n2_8116_7545 1.073016e-01
R8731 n2_8116_7545 n2_8116_7578 2.095238e-02
R8732 n2_8116_7578 n2_8116_7761 1.161905e-01
R8733 n2_8116_7761 n2_8116_7794 2.095238e-02
R8734 n2_8116_7794 n2_8116_7808 8.888889e-03
R8735 n2_8116_7808 n2_8116_7977 1.073016e-01
R8736 n2_8116_7977 n2_8116_8010 2.095238e-02
R8737 n2_8116_8010 n2_8116_8193 1.161905e-01
R8738 n2_8116_8193 n2_8116_8226 2.095238e-02
R8739 n2_8116_8226 n2_8116_8299 4.634921e-02
R8740 n2_8116_8395 n2_8116_8409 8.888889e-03
R8741 n2_8116_8409 n2_8116_8442 2.095238e-02
R8742 n2_8116_8442 n2_8116_8625 1.161905e-01
R8743 n2_8116_8625 n2_8116_8658 2.095238e-02
R8744 n2_8116_8658 n2_8116_8841 1.161905e-01
R8745 n2_8116_8841 n2_8116_8874 2.095238e-02
R8746 n2_8116_8874 n2_8116_8888 8.888889e-03
R8747 n2_8116_8888 n2_8116_9057 1.073016e-01
R8748 n2_8116_9057 n2_8116_9090 2.095238e-02
R8749 n2_8116_9090 n2_8116_9273 1.161905e-01
R8750 n2_8116_9273 n2_8116_9306 2.095238e-02
R8751 n2_8116_9306 n2_8116_9489 1.161905e-01
R8752 n2_8116_9489 n2_8116_9522 2.095238e-02
R8753 n2_8116_9522 n2_8116_9705 1.161905e-01
R8754 n2_8116_9705 n2_8116_9738 2.095238e-02
R8755 n2_8116_9738 n2_8116_9921 1.161905e-01
R8756 n2_8116_9921 n2_8116_9954 2.095238e-02
R8757 n2_8116_9954 n2_8116_9968 8.888889e-03
R8758 n2_8116_9968 n2_8116_10137 1.073016e-01
R8759 n2_8116_10137 n2_8116_10170 2.095238e-02
R8760 n2_8116_10170 n2_8116_10353 1.161905e-01
R8761 n2_8116_10353 n2_8116_10386 2.095238e-02
R8762 n2_8116_10386 n2_8116_10549 1.034921e-01
R8763 n2_8116_10549 n2_8116_10569 1.269841e-02
R8764 n2_8116_10645 n2_8116_10785 8.888889e-02
R8765 n2_8116_10785 n2_8116_10818 2.095238e-02
R8766 n2_8116_10818 n2_8116_11001 1.161905e-01
R8767 n2_8116_11001 n2_8116_11034 2.095238e-02
R8768 n2_8116_11034 n2_8116_11048 8.888889e-03
R8769 n2_8116_11048 n2_8116_11217 1.073016e-01
R8770 n2_8116_11217 n2_8116_11250 2.095238e-02
R8771 n2_8116_11250 n2_8116_11433 1.161905e-01
R8772 n2_8116_11433 n2_8116_11466 2.095238e-02
R8773 n2_8116_11466 n2_8116_11649 1.161905e-01
R8774 n2_8116_11649 n2_8116_11682 2.095238e-02
R8775 n2_8116_11682 n2_8116_11865 1.161905e-01
R8776 n2_8116_11865 n2_8116_11898 2.095238e-02
R8777 n2_8116_11898 n2_8116_12081 1.161905e-01
R8778 n2_8116_12081 n2_8116_12114 2.095238e-02
R8779 n2_8116_12114 n2_8116_12128 8.888889e-03
R8780 n2_8116_12128 n2_8116_12297 1.073016e-01
R8781 n2_8116_12297 n2_8116_12330 2.095238e-02
R8782 n2_8116_12330 n2_8116_12513 1.161905e-01
R8783 n2_8116_12513 n2_8116_12546 2.095238e-02
R8784 n2_8116_12546 n2_8116_12729 1.161905e-01
R8785 n2_8116_12729 n2_8116_12762 2.095238e-02
R8786 n2_8116_12762 n2_8116_12799 2.349206e-02
R8787 n2_8116_12895 n2_8116_12945 3.174603e-02
R8788 n2_8116_12945 n2_8116_12978 2.095238e-02
R8789 n2_8116_12978 n2_8116_13161 1.161905e-01
R8790 n2_8116_13161 n2_8116_13194 2.095238e-02
R8791 n2_8116_13194 n2_8116_13377 1.161905e-01
R8792 n2_8116_13377 n2_8116_13410 2.095238e-02
R8793 n2_8116_13410 n2_8116_13424 8.888889e-03
R8794 n2_8116_13424 n2_8116_13593 1.073016e-01
R8795 n2_8116_13593 n2_8116_13626 2.095238e-02
R8796 n2_8116_13626 n2_8116_13640 8.888889e-03
R8797 n2_8116_13640 n2_8116_13809 1.073016e-01
R8798 n2_8116_13809 n2_8116_13842 2.095238e-02
R8799 n2_8116_13842 n2_8116_13856 8.888889e-03
R8800 n2_8116_13856 n2_8116_13924 4.317460e-02
R8801 n2_8116_14020 n2_8116_14025 3.174603e-03
R8802 n2_8116_14025 n2_8116_14058 2.095238e-02
R8803 n2_8116_14058 n2_8116_14072 8.888889e-03
R8804 n2_8116_14072 n2_8116_14241 1.073016e-01
R8805 n2_8116_14241 n2_8116_14274 2.095238e-02
R8806 n2_8116_14274 n2_8116_14396 7.746032e-02
R8807 n2_8116_14396 n2_8116_14457 3.873016e-02
R8808 n2_8116_14457 n2_8116_14490 2.095238e-02
R8809 n2_8116_14490 n2_8116_14504 8.888889e-03
R8810 n2_8116_14504 n2_8116_14673 1.073016e-01
R8811 n2_8116_14673 n2_8116_14706 2.095238e-02
R8812 n2_8116_14706 n2_8116_14889 1.161905e-01
R8813 n2_8116_14889 n2_8116_14922 2.095238e-02
R8814 n2_8116_14922 n2_8116_15049 8.063492e-02
R8815 n2_8116_15138 n2_8116_15145 4.444444e-03
R8816 n2_8116_15145 n2_8116_15321 1.117460e-01
R8817 n2_8116_15321 n2_8116_15354 2.095238e-02
R8818 n2_8116_15354 n2_8116_15537 1.161905e-01
R8819 n2_8116_15537 n2_8116_15570 2.095238e-02
R8820 n2_8116_15570 n2_8116_15584 8.888889e-03
R8821 n2_8116_15584 n2_8116_15753 1.073016e-01
R8822 n2_8116_15753 n2_8116_15786 2.095238e-02
R8823 n2_8116_15786 n2_8116_15800 8.888889e-03
R8824 n2_8116_15800 n2_8116_15969 1.073016e-01
R8825 n2_8116_15969 n2_8116_16002 2.095238e-02
R8826 n2_8116_16002 n2_8116_16016 8.888889e-03
R8827 n2_8116_16016 n2_8116_16174 1.003175e-01
R8828 n2_8116_16174 n2_8116_16185 6.984127e-03
R8829 n2_8116_16270 n2_8116_16401 8.317460e-02
R8830 n2_8116_16401 n2_8116_16434 2.095238e-02
R8831 n2_8116_16434 n2_8116_16617 1.161905e-01
R8832 n2_8116_16617 n2_8116_16650 2.095238e-02
R8833 n2_8116_16650 n2_8116_16833 1.161905e-01
R8834 n2_8116_16833 n2_8116_16866 2.095238e-02
R8835 n2_8116_16866 n2_8116_17049 1.161905e-01
R8836 n2_8116_17049 n2_8116_17082 2.095238e-02
R8837 n2_8116_17082 n2_8116_17096 8.888889e-03
R8838 n2_8116_17096 n2_8116_17119 1.460317e-02
R8839 n2_8116_17119 n2_8116_17265 9.269841e-02
R8840 n2_8116_17265 n2_8116_17298 2.095238e-02
R8841 n2_8116_17298 n2_8116_17299 6.349206e-04
R8842 n2_8116_17299 n2_8116_17312 8.253968e-03
R8843 n2_8116_17395 n2_8116_17481 5.460317e-02
R8844 n2_8116_17481 n2_8116_17514 2.095238e-02
R8845 n2_8116_17514 n2_8116_17697 1.161905e-01
R8846 n2_8116_17697 n2_8116_17730 2.095238e-02
R8847 n2_8116_17730 n2_8116_17913 1.161905e-01
R8848 n2_8116_17913 n2_8116_17946 2.095238e-02
R8849 n2_8116_17946 n2_8116_18129 1.161905e-01
R8850 n2_8116_18129 n2_8116_18162 2.095238e-02
R8851 n2_8116_18162 n2_8116_18345 1.161905e-01
R8852 n2_8116_18345 n2_8116_18378 2.095238e-02
R8853 n2_8116_18378 n2_8116_18392 8.888889e-03
R8854 n2_8116_18392 n2_8116_18421 1.841270e-02
R8855 n2_8116_18421 n2_8116_18424 1.904762e-03
R8856 n2_8116_18520 n2_8116_18561 2.603175e-02
R8857 n2_8116_18561 n2_8116_18594 2.095238e-02
R8858 n2_8116_18594 n2_8116_18608 8.888889e-03
R8859 n2_8116_18608 n2_8116_18777 1.073016e-01
R8860 n2_8116_18777 n2_8116_18810 2.095238e-02
R8861 n2_8116_18810 n2_8116_18993 1.161905e-01
R8862 n2_8116_18993 n2_8116_19026 2.095238e-02
R8863 n2_8116_19026 n2_8116_19209 1.161905e-01
R8864 n2_8116_19209 n2_8116_19242 2.095238e-02
R8865 n2_8116_19242 n2_8116_19256 8.888889e-03
R8866 n2_8116_19256 n2_8116_19279 1.460317e-02
R8867 n2_8116_19279 n2_8116_19425 9.269841e-02
R8868 n2_8116_19425 n2_8116_19458 2.095238e-02
R8869 n2_8116_19458 n2_8116_19549 5.777778e-02
R8870 n2_8116_19641 n2_8116_19645 2.539683e-03
R8871 n2_8116_19645 n2_8116_19674 1.841270e-02
R8872 n2_8116_19674 n2_8116_19857 1.161905e-01
R8873 n2_8116_19857 n2_8116_19890 2.095238e-02
R8874 n2_8116_19890 n2_8116_20073 1.161905e-01
R8875 n2_8116_20073 n2_8116_20106 2.095238e-02
R8876 n2_8116_20106 n2_8116_20289 1.161905e-01
R8877 n2_8116_20289 n2_8116_20322 2.095238e-02
R8878 n2_8116_20322 n2_8116_20505 1.161905e-01
R8879 n2_8116_20505 n2_8116_20538 2.095238e-02
R8880 n2_8116_20538 n2_8116_20674 8.634921e-02
R8881 n2_8116_20754 n2_8116_20770 1.015873e-02
R8882 n2_8116_20770 n2_8116_20937 1.060317e-01
R8883 n2_8116_20937 n2_8116_20970 2.095238e-02
R8884 n2_8116_8395 n2_8208_8395 5.841270e-02
R8885 n2_8208_8395 n2_8255_8395 2.984127e-02
R8886 n2_8255_8395 n2_8304_8395 3.111111e-02
R8887 n2_8116_10549 n2_8255_10549 8.825397e-02
R8888 n2_8255_10549 n2_8304_10549 3.111111e-02
R8889 n2_8116_10645 n2_8255_10645 8.825397e-02
R8890 n2_8255_10645 n2_8304_10645 3.111111e-02
R8891 n2_8116_12799 n2_8208_12799 5.841270e-02
R8892 n2_8208_12799 n2_8255_12799 2.984127e-02
R8893 n2_8255_12799 n2_8304_12799 3.111111e-02
R8894 n2_8116_424 n2_8208_424 5.841270e-02
R8895 n2_8208_424 n2_8255_424 2.984127e-02
R8896 n2_8255_424 n2_8304_424 3.111111e-02
R8897 n2_8304_424 n2_8396_424 5.841270e-02
R8898 n2_8116_520 n2_8208_520 5.841270e-02
R8899 n2_8208_520 n2_8255_520 2.984127e-02
R8900 n2_8255_520 n2_8304_520 3.111111e-02
R8901 n2_8304_520 n2_8396_520 5.841270e-02
R8902 n2_8116_1549 n2_8208_1549 5.841270e-02
R8903 n2_8208_1549 n2_8255_1549 2.984127e-02
R8904 n2_8255_1549 n2_8304_1549 3.111111e-02
R8905 n2_8304_1549 n2_8396_1549 5.841270e-02
R8906 n2_8116_1645 n2_8208_1645 5.841270e-02
R8907 n2_8208_1645 n2_8255_1645 2.984127e-02
R8908 n2_8255_1645 n2_8304_1645 3.111111e-02
R8909 n2_8304_1645 n2_8396_1645 5.841270e-02
R8910 n2_8116_2674 n2_8208_2674 5.841270e-02
R8911 n2_8208_2674 n2_8255_2674 2.984127e-02
R8912 n2_8255_2674 n2_8304_2674 3.111111e-02
R8913 n2_8304_2674 n2_8396_2674 5.841270e-02
R8914 n2_8116_2770 n2_8208_2770 5.841270e-02
R8915 n2_8208_2770 n2_8255_2770 2.984127e-02
R8916 n2_8255_2770 n2_8304_2770 3.111111e-02
R8917 n2_8304_2770 n2_8396_2770 5.841270e-02
R8918 n2_8116_3799 n2_8208_3799 5.841270e-02
R8919 n2_8208_3799 n2_8255_3799 2.984127e-02
R8920 n2_8255_3799 n2_8304_3799 3.111111e-02
R8921 n2_8304_3799 n2_8396_3799 5.841270e-02
R8922 n2_8116_3895 n2_8208_3895 5.841270e-02
R8923 n2_8208_3895 n2_8255_3895 2.984127e-02
R8924 n2_8255_3895 n2_8304_3895 3.111111e-02
R8925 n2_8304_3895 n2_8396_3895 5.841270e-02
R8926 n2_8116_4924 n2_8208_4924 5.841270e-02
R8927 n2_8208_4924 n2_8255_4924 2.984127e-02
R8928 n2_8255_4924 n2_8304_4924 3.111111e-02
R8929 n2_8304_4924 n2_8396_4924 5.841270e-02
R8930 n2_8116_5020 n2_8208_5020 5.841270e-02
R8931 n2_8208_5020 n2_8255_5020 2.984127e-02
R8932 n2_8255_5020 n2_8304_5020 3.111111e-02
R8933 n2_8304_5020 n2_8396_5020 5.841270e-02
R8934 n2_8116_6049 n2_8208_6049 5.841270e-02
R8935 n2_8208_6049 n2_8255_6049 2.984127e-02
R8936 n2_8255_6049 n2_8304_6049 3.111111e-02
R8937 n2_8304_6049 n2_8396_6049 5.841270e-02
R8938 n2_8116_6145 n2_8208_6145 5.841270e-02
R8939 n2_8208_6145 n2_8255_6145 2.984127e-02
R8940 n2_8255_6145 n2_8304_6145 3.111111e-02
R8941 n2_8304_6145 n2_8396_6145 5.841270e-02
R8942 n2_8116_7174 n2_8208_7174 5.841270e-02
R8943 n2_8208_7174 n2_8255_7174 2.984127e-02
R8944 n2_8255_7174 n2_8304_7174 3.111111e-02
R8945 n2_8304_7174 n2_8396_7174 5.841270e-02
R8946 n2_8116_7270 n2_8208_7270 5.841270e-02
R8947 n2_8208_7270 n2_8255_7270 2.984127e-02
R8948 n2_8255_7270 n2_8304_7270 3.111111e-02
R8949 n2_8304_7270 n2_8396_7270 5.841270e-02
R8950 n2_8116_8299 n2_8208_8299 5.841270e-02
R8951 n2_8208_8299 n2_8255_8299 2.984127e-02
R8952 n2_8255_8299 n2_8304_8299 3.111111e-02
R8953 n2_8304_8299 n2_8396_8299 5.841270e-02
R8954 n2_8116_12895 n2_8208_12895 5.841270e-02
R8955 n2_8208_12895 n2_8255_12895 2.984127e-02
R8956 n2_8255_12895 n2_8304_12895 3.111111e-02
R8957 n2_8304_12895 n2_8396_12895 5.841270e-02
R8958 n2_8116_13924 n2_8208_13924 5.841270e-02
R8959 n2_8208_13924 n2_8255_13924 2.984127e-02
R8960 n2_8255_13924 n2_8304_13924 3.111111e-02
R8961 n2_8304_13924 n2_8396_13924 5.841270e-02
R8962 n2_8116_14020 n2_8208_14020 5.841270e-02
R8963 n2_8208_14020 n2_8255_14020 2.984127e-02
R8964 n2_8255_14020 n2_8304_14020 3.111111e-02
R8965 n2_8304_14020 n2_8396_14020 5.841270e-02
R8966 n2_8116_15049 n2_8208_15049 5.841270e-02
R8967 n2_8208_15049 n2_8255_15049 2.984127e-02
R8968 n2_8255_15049 n2_8304_15049 3.111111e-02
R8969 n2_8304_15049 n2_8396_15049 5.841270e-02
R8970 n2_8116_15145 n2_8208_15145 5.841270e-02
R8971 n2_8208_15145 n2_8255_15145 2.984127e-02
R8972 n2_8255_15145 n2_8304_15145 3.111111e-02
R8973 n2_8304_15145 n2_8396_15145 5.841270e-02
R8974 n2_8116_16174 n2_8208_16174 5.841270e-02
R8975 n2_8208_16174 n2_8255_16174 2.984127e-02
R8976 n2_8255_16174 n2_8304_16174 3.111111e-02
R8977 n2_8304_16174 n2_8396_16174 5.841270e-02
R8978 n2_8116_16270 n2_8208_16270 5.841270e-02
R8979 n2_8208_16270 n2_8255_16270 2.984127e-02
R8980 n2_8255_16270 n2_8304_16270 3.111111e-02
R8981 n2_8304_16270 n2_8396_16270 5.841270e-02
R8982 n2_8116_17299 n2_8208_17299 5.841270e-02
R8983 n2_8208_17299 n2_8255_17299 2.984127e-02
R8984 n2_8255_17299 n2_8304_17299 3.111111e-02
R8985 n2_8304_17299 n2_8396_17299 5.841270e-02
R8986 n2_8116_17395 n2_8208_17395 5.841270e-02
R8987 n2_8208_17395 n2_8255_17395 2.984127e-02
R8988 n2_8255_17395 n2_8304_17395 3.111111e-02
R8989 n2_8304_17395 n2_8396_17395 5.841270e-02
R8990 n2_8116_18424 n2_8208_18424 5.841270e-02
R8991 n2_8208_18424 n2_8255_18424 2.984127e-02
R8992 n2_8255_18424 n2_8304_18424 3.111111e-02
R8993 n2_8304_18424 n2_8396_18424 5.841270e-02
R8994 n2_8116_18520 n2_8208_18520 5.841270e-02
R8995 n2_8208_18520 n2_8255_18520 2.984127e-02
R8996 n2_8255_18520 n2_8304_18520 3.111111e-02
R8997 n2_8304_18520 n2_8396_18520 5.841270e-02
R8998 n2_8116_19549 n2_8208_19549 5.841270e-02
R8999 n2_8208_19549 n2_8255_19549 2.984127e-02
R9000 n2_8255_19549 n2_8304_19549 3.111111e-02
R9001 n2_8304_19549 n2_8396_19549 5.841270e-02
R9002 n2_8116_19645 n2_8208_19645 5.841270e-02
R9003 n2_8208_19645 n2_8255_19645 2.984127e-02
R9004 n2_8255_19645 n2_8304_19645 3.111111e-02
R9005 n2_8304_19645 n2_8396_19645 5.841270e-02
R9006 n2_8116_20674 n2_8208_20674 5.841270e-02
R9007 n2_8208_20674 n2_8255_20674 2.984127e-02
R9008 n2_8255_20674 n2_8304_20674 3.111111e-02
R9009 n2_8304_20674 n2_8396_20674 5.841270e-02
R9010 n2_8116_20770 n2_8208_20770 5.841270e-02
R9011 n2_8208_20770 n2_8255_20770 2.984127e-02
R9012 n2_8255_20770 n2_8304_20770 3.111111e-02
R9013 n2_8304_20770 n2_8396_20770 5.841270e-02
R9014 n2_8208_201 n2_8208_234 2.095238e-02
R9015 n2_8208_234 n2_8208_417 1.161905e-01
R9016 n2_8208_417 n2_8208_424 4.444444e-03
R9017 n2_8208_424 n2_8208_450 1.650794e-02
R9018 n2_8208_450 n2_8208_520 4.444444e-02
R9019 n2_8208_520 n2_8208_633 7.174603e-02
R9020 n2_8208_633 n2_8208_666 2.095238e-02
R9021 n2_8208_666 n2_8208_849 1.161905e-01
R9022 n2_8208_849 n2_8208_882 2.095238e-02
R9023 n2_8208_882 n2_8208_1065 1.161905e-01
R9024 n2_8208_1065 n2_8208_1098 2.095238e-02
R9025 n2_8208_1098 n2_8208_1281 1.161905e-01
R9026 n2_8208_1281 n2_8208_1314 2.095238e-02
R9027 n2_8208_1314 n2_8208_1497 1.161905e-01
R9028 n2_8208_1497 n2_8208_1530 2.095238e-02
R9029 n2_8208_1530 n2_8208_1549 1.206349e-02
R9030 n2_8208_1549 n2_8208_1645 6.095238e-02
R9031 n2_8208_1645 n2_8208_1713 4.317460e-02
R9032 n2_8208_1713 n2_8208_1746 2.095238e-02
R9033 n2_8208_1746 n2_8208_1760 8.888889e-03
R9034 n2_8208_1760 n2_8208_1783 1.460317e-02
R9035 n2_8208_1783 n2_8208_1929 9.269841e-02
R9036 n2_8208_1929 n2_8208_1962 2.095238e-02
R9037 n2_8208_1962 n2_8208_2145 1.161905e-01
R9038 n2_8208_2145 n2_8208_2178 2.095238e-02
R9039 n2_8208_2178 n2_8208_2361 1.161905e-01
R9040 n2_8208_2361 n2_8208_2394 2.095238e-02
R9041 n2_8208_2394 n2_8208_2408 8.888889e-03
R9042 n2_8208_2408 n2_8208_2577 1.073016e-01
R9043 n2_8208_2577 n2_8208_2610 2.095238e-02
R9044 n2_8208_2610 n2_8208_2674 4.063492e-02
R9045 n2_8208_2674 n2_8208_2770 6.095238e-02
R9046 n2_8208_2770 n2_8208_2793 1.460317e-02
R9047 n2_8208_2793 n2_8208_2826 2.095238e-02
R9048 n2_8208_2826 n2_8208_2840 8.888889e-03
R9049 n2_8208_2840 n2_8208_2863 1.460317e-02
R9050 n2_8208_2863 n2_8208_3009 9.269841e-02
R9051 n2_8208_3009 n2_8208_3042 2.095238e-02
R9052 n2_8208_3042 n2_8208_3225 1.161905e-01
R9053 n2_8208_3225 n2_8208_3258 2.095238e-02
R9054 n2_8208_3258 n2_8208_3441 1.161905e-01
R9055 n2_8208_3441 n2_8208_3474 2.095238e-02
R9056 n2_8208_3474 n2_8208_3488 8.888889e-03
R9057 n2_8208_3488 n2_8208_3657 1.073016e-01
R9058 n2_8208_3657 n2_8208_3690 2.095238e-02
R9059 n2_8208_3690 n2_8208_3799 6.920635e-02
R9060 n2_8208_3799 n2_8208_3873 4.698413e-02
R9061 n2_8208_3873 n2_8208_3895 1.396825e-02
R9062 n2_8208_3895 n2_8208_3906 6.984127e-03
R9063 n2_8208_3906 n2_8208_4089 1.161905e-01
R9064 n2_8208_4089 n2_8208_4122 2.095238e-02
R9065 n2_8208_4122 n2_8208_4136 8.888889e-03
R9066 n2_8208_4136 n2_8208_4305 1.073016e-01
R9067 n2_8208_4305 n2_8208_4338 2.095238e-02
R9068 n2_8208_4338 n2_8208_4521 1.161905e-01
R9069 n2_8208_4521 n2_8208_4554 2.095238e-02
R9070 n2_8208_4554 n2_8208_4568 8.888889e-03
R9071 n2_8208_4568 n2_8208_4737 1.073016e-01
R9072 n2_8208_4737 n2_8208_4770 2.095238e-02
R9073 n2_8208_4770 n2_8208_4924 9.777778e-02
R9074 n2_8208_4924 n2_8208_4953 1.841270e-02
R9075 n2_8208_4953 n2_8208_4986 2.095238e-02
R9076 n2_8208_4986 n2_8208_5020 2.158730e-02
R9077 n2_8208_5020 n2_8208_5169 9.460317e-02
R9078 n2_8208_5169 n2_8208_5202 2.095238e-02
R9079 n2_8208_5202 n2_8208_5216 8.888889e-03
R9080 n2_8208_5216 n2_8208_5239 1.460317e-02
R9081 n2_8208_5239 n2_8208_5385 9.269841e-02
R9082 n2_8208_5385 n2_8208_5418 2.095238e-02
R9083 n2_8208_5418 n2_8208_5432 8.888889e-03
R9084 n2_8208_5432 n2_8208_5455 1.460317e-02
R9085 n2_8208_5455 n2_8208_5601 9.269841e-02
R9086 n2_8208_5601 n2_8208_5634 2.095238e-02
R9087 n2_8208_5634 n2_8208_5817 1.161905e-01
R9088 n2_8208_5817 n2_8208_5850 2.095238e-02
R9089 n2_8208_5850 n2_8208_6033 1.161905e-01
R9090 n2_8208_6033 n2_8208_6049 1.015873e-02
R9091 n2_8208_6049 n2_8208_6066 1.079365e-02
R9092 n2_8208_6066 n2_8208_6145 5.015873e-02
R9093 n2_8208_6145 n2_8208_6249 6.603175e-02
R9094 n2_8208_6249 n2_8208_6282 2.095238e-02
R9095 n2_8208_6282 n2_8208_6465 1.161905e-01
R9096 n2_8208_6465 n2_8208_6498 2.095238e-02
R9097 n2_8208_6498 n2_8208_6512 8.888889e-03
R9098 n2_8208_6512 n2_8208_6535 1.460317e-02
R9099 n2_8208_6535 n2_8208_6681 9.269841e-02
R9100 n2_8208_6681 n2_8208_6714 2.095238e-02
R9101 n2_8208_6714 n2_8208_6897 1.161905e-01
R9102 n2_8208_6897 n2_8208_6930 2.095238e-02
R9103 n2_8208_6930 n2_8208_6944 8.888889e-03
R9104 n2_8208_6944 n2_8208_7113 1.073016e-01
R9105 n2_8208_7113 n2_8208_7146 2.095238e-02
R9106 n2_8208_7146 n2_8208_7160 8.888889e-03
R9107 n2_8208_7160 n2_8208_7174 8.888889e-03
R9108 n2_8208_7174 n2_8208_7270 6.095238e-02
R9109 n2_8208_7270 n2_8208_7329 3.746032e-02
R9110 n2_8208_7329 n2_8208_7362 2.095238e-02
R9111 n2_8208_7362 n2_8208_7376 8.888889e-03
R9112 n2_8208_7376 n2_8208_7545 1.073016e-01
R9113 n2_8208_7545 n2_8208_7578 2.095238e-02
R9114 n2_8208_7578 n2_8208_7761 1.161905e-01
R9115 n2_8208_7761 n2_8208_7794 2.095238e-02
R9116 n2_8208_7794 n2_8208_7808 8.888889e-03
R9117 n2_8208_7808 n2_8208_7977 1.073016e-01
R9118 n2_8208_7977 n2_8208_8010 2.095238e-02
R9119 n2_8208_8010 n2_8208_8193 1.161905e-01
R9120 n2_8208_8193 n2_8208_8226 2.095238e-02
R9121 n2_8208_8226 n2_8208_8299 4.634921e-02
R9122 n2_8208_8299 n2_8208_8395 6.095238e-02
R9123 n2_8208_8395 n2_8208_8409 8.888889e-03
R9124 n2_8208_8409 n2_8208_8442 2.095238e-02
R9125 n2_8208_12762 n2_8208_12799 2.349206e-02
R9126 n2_8208_12799 n2_8208_12895 6.095238e-02
R9127 n2_8208_12895 n2_8208_12945 3.174603e-02
R9128 n2_8208_12945 n2_8208_12978 2.095238e-02
R9129 n2_8208_12978 n2_8208_13161 1.161905e-01
R9130 n2_8208_13161 n2_8208_13194 2.095238e-02
R9131 n2_8208_13194 n2_8208_13377 1.161905e-01
R9132 n2_8208_13377 n2_8208_13410 2.095238e-02
R9133 n2_8208_13410 n2_8208_13424 8.888889e-03
R9134 n2_8208_13424 n2_8208_13593 1.073016e-01
R9135 n2_8208_13593 n2_8208_13626 2.095238e-02
R9136 n2_8208_13626 n2_8208_13640 8.888889e-03
R9137 n2_8208_13640 n2_8208_13809 1.073016e-01
R9138 n2_8208_13809 n2_8208_13842 2.095238e-02
R9139 n2_8208_13842 n2_8208_13856 8.888889e-03
R9140 n2_8208_13856 n2_8208_13924 4.317460e-02
R9141 n2_8208_13924 n2_8208_14020 6.095238e-02
R9142 n2_8208_14020 n2_8208_14025 3.174603e-03
R9143 n2_8208_14025 n2_8208_14058 2.095238e-02
R9144 n2_8208_14058 n2_8208_14072 8.888889e-03
R9145 n2_8208_14072 n2_8208_14241 1.073016e-01
R9146 n2_8208_14241 n2_8208_14274 2.095238e-02
R9147 n2_8208_14274 n2_8208_14396 7.746032e-02
R9148 n2_8208_14396 n2_8208_14457 3.873016e-02
R9149 n2_8208_14457 n2_8208_14490 2.095238e-02
R9150 n2_8208_14490 n2_8208_14504 8.888889e-03
R9151 n2_8208_14504 n2_8208_14673 1.073016e-01
R9152 n2_8208_14673 n2_8208_14706 2.095238e-02
R9153 n2_8208_14706 n2_8208_14889 1.161905e-01
R9154 n2_8208_14889 n2_8208_14922 2.095238e-02
R9155 n2_8208_14922 n2_8208_15049 8.063492e-02
R9156 n2_8208_15049 n2_8208_15105 3.555556e-02
R9157 n2_8208_15105 n2_8208_15138 2.095238e-02
R9158 n2_8208_15138 n2_8208_15145 4.444444e-03
R9159 n2_8208_15145 n2_8208_15321 1.117460e-01
R9160 n2_8208_15321 n2_8208_15354 2.095238e-02
R9161 n2_8208_15354 n2_8208_15537 1.161905e-01
R9162 n2_8208_15537 n2_8208_15570 2.095238e-02
R9163 n2_8208_15570 n2_8208_15584 8.888889e-03
R9164 n2_8208_15584 n2_8208_15753 1.073016e-01
R9165 n2_8208_15753 n2_8208_15786 2.095238e-02
R9166 n2_8208_15786 n2_8208_15800 8.888889e-03
R9167 n2_8208_15800 n2_8208_15969 1.073016e-01
R9168 n2_8208_15969 n2_8208_16002 2.095238e-02
R9169 n2_8208_16002 n2_8208_16016 8.888889e-03
R9170 n2_8208_16016 n2_8208_16174 1.003175e-01
R9171 n2_8208_16174 n2_8208_16185 6.984127e-03
R9172 n2_8208_16185 n2_8208_16218 2.095238e-02
R9173 n2_8208_16218 n2_8208_16270 3.301587e-02
R9174 n2_8208_16270 n2_8208_16401 8.317460e-02
R9175 n2_8208_16401 n2_8208_16434 2.095238e-02
R9176 n2_8208_16434 n2_8208_16617 1.161905e-01
R9177 n2_8208_16617 n2_8208_16650 2.095238e-02
R9178 n2_8208_16650 n2_8208_16833 1.161905e-01
R9179 n2_8208_16833 n2_8208_16866 2.095238e-02
R9180 n2_8208_16866 n2_8208_17049 1.161905e-01
R9181 n2_8208_17049 n2_8208_17082 2.095238e-02
R9182 n2_8208_17082 n2_8208_17096 8.888889e-03
R9183 n2_8208_17096 n2_8208_17119 1.460317e-02
R9184 n2_8208_17119 n2_8208_17265 9.269841e-02
R9185 n2_8208_17265 n2_8208_17298 2.095238e-02
R9186 n2_8208_17298 n2_8208_17299 6.349206e-04
R9187 n2_8208_17299 n2_8208_17312 8.253968e-03
R9188 n2_8208_17312 n2_8208_17395 5.269841e-02
R9189 n2_8208_17395 n2_8208_17481 5.460317e-02
R9190 n2_8208_17481 n2_8208_17514 2.095238e-02
R9191 n2_8208_17514 n2_8208_17697 1.161905e-01
R9192 n2_8208_17697 n2_8208_17730 2.095238e-02
R9193 n2_8208_17730 n2_8208_17913 1.161905e-01
R9194 n2_8208_17913 n2_8208_17946 2.095238e-02
R9195 n2_8208_17946 n2_8208_18129 1.161905e-01
R9196 n2_8208_18129 n2_8208_18162 2.095238e-02
R9197 n2_8208_18162 n2_8208_18345 1.161905e-01
R9198 n2_8208_18345 n2_8208_18378 2.095238e-02
R9199 n2_8208_18378 n2_8208_18392 8.888889e-03
R9200 n2_8208_18392 n2_8208_18421 1.841270e-02
R9201 n2_8208_18421 n2_8208_18424 1.904762e-03
R9202 n2_8208_18424 n2_8208_18520 6.095238e-02
R9203 n2_8208_18520 n2_8208_18561 2.603175e-02
R9204 n2_8208_18561 n2_8208_18594 2.095238e-02
R9205 n2_8208_18594 n2_8208_18608 8.888889e-03
R9206 n2_8208_18608 n2_8208_18777 1.073016e-01
R9207 n2_8208_18777 n2_8208_18810 2.095238e-02
R9208 n2_8208_18810 n2_8208_18993 1.161905e-01
R9209 n2_8208_18993 n2_8208_19026 2.095238e-02
R9210 n2_8208_19026 n2_8208_19209 1.161905e-01
R9211 n2_8208_19209 n2_8208_19242 2.095238e-02
R9212 n2_8208_19242 n2_8208_19256 8.888889e-03
R9213 n2_8208_19256 n2_8208_19279 1.460317e-02
R9214 n2_8208_19279 n2_8208_19425 9.269841e-02
R9215 n2_8208_19425 n2_8208_19458 2.095238e-02
R9216 n2_8208_19458 n2_8208_19549 5.777778e-02
R9217 n2_8208_19549 n2_8208_19641 5.841270e-02
R9218 n2_8208_19641 n2_8208_19645 2.539683e-03
R9219 n2_8208_19645 n2_8208_19674 1.841270e-02
R9220 n2_8208_19674 n2_8208_19857 1.161905e-01
R9221 n2_8208_19857 n2_8208_19890 2.095238e-02
R9222 n2_8208_19890 n2_8208_20073 1.161905e-01
R9223 n2_8208_20073 n2_8208_20106 2.095238e-02
R9224 n2_8208_20106 n2_8208_20289 1.161905e-01
R9225 n2_8208_20289 n2_8208_20322 2.095238e-02
R9226 n2_8208_20322 n2_8208_20505 1.161905e-01
R9227 n2_8208_20505 n2_8208_20538 2.095238e-02
R9228 n2_8208_20538 n2_8208_20674 8.634921e-02
R9229 n2_8208_20674 n2_8208_20721 2.984127e-02
R9230 n2_8208_20721 n2_8208_20754 2.095238e-02
R9231 n2_8208_20754 n2_8208_20770 1.015873e-02
R9232 n2_8208_20770 n2_8208_20937 1.060317e-01
R9233 n2_8208_20937 n2_8208_20970 2.095238e-02
R9234 n2_8304_201 n2_8304_234 2.095238e-02
R9235 n2_8304_234 n2_8304_417 1.161905e-01
R9236 n2_8304_417 n2_8304_424 4.444444e-03
R9237 n2_8304_424 n2_8304_450 1.650794e-02
R9238 n2_8304_450 n2_8304_520 4.444444e-02
R9239 n2_8304_520 n2_8304_633 7.174603e-02
R9240 n2_8304_633 n2_8304_666 2.095238e-02
R9241 n2_8304_666 n2_8304_849 1.161905e-01
R9242 n2_8304_849 n2_8304_882 2.095238e-02
R9243 n2_8304_882 n2_8304_1065 1.161905e-01
R9244 n2_8304_1065 n2_8304_1098 2.095238e-02
R9245 n2_8304_1098 n2_8304_1281 1.161905e-01
R9246 n2_8304_1281 n2_8304_1314 2.095238e-02
R9247 n2_8304_1314 n2_8304_1497 1.161905e-01
R9248 n2_8304_1497 n2_8304_1530 2.095238e-02
R9249 n2_8304_1530 n2_8304_1549 1.206349e-02
R9250 n2_8304_1549 n2_8304_1645 6.095238e-02
R9251 n2_8304_1645 n2_8304_1713 4.317460e-02
R9252 n2_8304_1713 n2_8304_1746 2.095238e-02
R9253 n2_8304_1746 n2_8304_1760 8.888889e-03
R9254 n2_8304_1760 n2_8304_1783 1.460317e-02
R9255 n2_8304_1783 n2_8304_1929 9.269841e-02
R9256 n2_8304_1929 n2_8304_1962 2.095238e-02
R9257 n2_8304_1962 n2_8304_2145 1.161905e-01
R9258 n2_8304_2145 n2_8304_2178 2.095238e-02
R9259 n2_8304_2178 n2_8304_2361 1.161905e-01
R9260 n2_8304_2361 n2_8304_2394 2.095238e-02
R9261 n2_8304_2394 n2_8304_2408 8.888889e-03
R9262 n2_8304_2408 n2_8304_2577 1.073016e-01
R9263 n2_8304_2577 n2_8304_2610 2.095238e-02
R9264 n2_8304_2610 n2_8304_2674 4.063492e-02
R9265 n2_8304_2674 n2_8304_2770 6.095238e-02
R9266 n2_8304_2770 n2_8304_2793 1.460317e-02
R9267 n2_8304_2793 n2_8304_2826 2.095238e-02
R9268 n2_8304_2826 n2_8304_2840 8.888889e-03
R9269 n2_8304_2840 n2_8304_2863 1.460317e-02
R9270 n2_8304_2863 n2_8304_3009 9.269841e-02
R9271 n2_8304_3009 n2_8304_3042 2.095238e-02
R9272 n2_8304_3042 n2_8304_3225 1.161905e-01
R9273 n2_8304_3225 n2_8304_3258 2.095238e-02
R9274 n2_8304_3258 n2_8304_3441 1.161905e-01
R9275 n2_8304_3441 n2_8304_3474 2.095238e-02
R9276 n2_8304_3474 n2_8304_3488 8.888889e-03
R9277 n2_8304_3488 n2_8304_3657 1.073016e-01
R9278 n2_8304_3657 n2_8304_3690 2.095238e-02
R9279 n2_8304_3690 n2_8304_3799 6.920635e-02
R9280 n2_8304_3799 n2_8304_3873 4.698413e-02
R9281 n2_8304_3873 n2_8304_3895 1.396825e-02
R9282 n2_8304_3895 n2_8304_3906 6.984127e-03
R9283 n2_8304_3906 n2_8304_4089 1.161905e-01
R9284 n2_8304_4089 n2_8304_4122 2.095238e-02
R9285 n2_8304_4122 n2_8304_4136 8.888889e-03
R9286 n2_8304_4136 n2_8304_4305 1.073016e-01
R9287 n2_8304_4305 n2_8304_4338 2.095238e-02
R9288 n2_8304_4338 n2_8304_4521 1.161905e-01
R9289 n2_8304_4521 n2_8304_4554 2.095238e-02
R9290 n2_8304_4554 n2_8304_4568 8.888889e-03
R9291 n2_8304_4568 n2_8304_4737 1.073016e-01
R9292 n2_8304_4737 n2_8304_4770 2.095238e-02
R9293 n2_8304_4770 n2_8304_4924 9.777778e-02
R9294 n2_8304_4924 n2_8304_4953 1.841270e-02
R9295 n2_8304_4953 n2_8304_4986 2.095238e-02
R9296 n2_8304_4986 n2_8304_5020 2.158730e-02
R9297 n2_8304_5020 n2_8304_5169 9.460317e-02
R9298 n2_8304_5169 n2_8304_5202 2.095238e-02
R9299 n2_8304_5202 n2_8304_5216 8.888889e-03
R9300 n2_8304_5216 n2_8304_5239 1.460317e-02
R9301 n2_8304_5239 n2_8304_5385 9.269841e-02
R9302 n2_8304_5385 n2_8304_5418 2.095238e-02
R9303 n2_8304_5418 n2_8304_5432 8.888889e-03
R9304 n2_8304_5432 n2_8304_5455 1.460317e-02
R9305 n2_8304_5455 n2_8304_5601 9.269841e-02
R9306 n2_8304_5601 n2_8304_5634 2.095238e-02
R9307 n2_8304_5634 n2_8304_5817 1.161905e-01
R9308 n2_8304_5817 n2_8304_5850 2.095238e-02
R9309 n2_8304_5850 n2_8304_6033 1.161905e-01
R9310 n2_8304_6033 n2_8304_6049 1.015873e-02
R9311 n2_8304_6049 n2_8304_6066 1.079365e-02
R9312 n2_8304_6066 n2_8304_6145 5.015873e-02
R9313 n2_8304_6145 n2_8304_6249 6.603175e-02
R9314 n2_8304_6249 n2_8304_6282 2.095238e-02
R9315 n2_8304_6282 n2_8304_6465 1.161905e-01
R9316 n2_8304_6465 n2_8304_6498 2.095238e-02
R9317 n2_8304_6498 n2_8304_6512 8.888889e-03
R9318 n2_8304_6512 n2_8304_6535 1.460317e-02
R9319 n2_8304_6535 n2_8304_6681 9.269841e-02
R9320 n2_8304_6681 n2_8304_6714 2.095238e-02
R9321 n2_8304_6714 n2_8304_6897 1.161905e-01
R9322 n2_8304_6897 n2_8304_6930 2.095238e-02
R9323 n2_8304_6930 n2_8304_6944 8.888889e-03
R9324 n2_8304_6944 n2_8304_7113 1.073016e-01
R9325 n2_8304_7113 n2_8304_7146 2.095238e-02
R9326 n2_8304_7146 n2_8304_7160 8.888889e-03
R9327 n2_8304_7160 n2_8304_7174 8.888889e-03
R9328 n2_8304_7174 n2_8304_7270 6.095238e-02
R9329 n2_8304_7270 n2_8304_7329 3.746032e-02
R9330 n2_8304_7329 n2_8304_7362 2.095238e-02
R9331 n2_8304_7362 n2_8304_7376 8.888889e-03
R9332 n2_8304_7376 n2_8304_7545 1.073016e-01
R9333 n2_8304_7545 n2_8304_7578 2.095238e-02
R9334 n2_8304_7578 n2_8304_7761 1.161905e-01
R9335 n2_8304_7761 n2_8304_7794 2.095238e-02
R9336 n2_8304_7794 n2_8304_7808 8.888889e-03
R9337 n2_8304_7808 n2_8304_7977 1.073016e-01
R9338 n2_8304_7977 n2_8304_8010 2.095238e-02
R9339 n2_8304_8010 n2_8304_8193 1.161905e-01
R9340 n2_8304_8193 n2_8304_8226 2.095238e-02
R9341 n2_8304_8226 n2_8304_8299 4.634921e-02
R9342 n2_8304_8299 n2_8304_8395 6.095238e-02
R9343 n2_8304_8395 n2_8304_8409 8.888889e-03
R9344 n2_8304_8409 n2_8304_8442 2.095238e-02
R9345 n2_8304_8442 n2_8304_8625 1.161905e-01
R9346 n2_8304_8625 n2_8304_8658 2.095238e-02
R9347 n2_8304_8658 n2_8304_8841 1.161905e-01
R9348 n2_8304_8841 n2_8304_8874 2.095238e-02
R9349 n2_8304_8874 n2_8304_8888 8.888889e-03
R9350 n2_8304_8888 n2_8304_8909 1.333333e-02
R9351 n2_8304_8909 n2_8304_9057 9.396825e-02
R9352 n2_8304_9057 n2_8304_9090 2.095238e-02
R9353 n2_8304_9090 n2_8304_9273 1.161905e-01
R9354 n2_8304_9273 n2_8304_9306 2.095238e-02
R9355 n2_8304_9705 n2_8304_9738 2.095238e-02
R9356 n2_8304_9738 n2_8304_9921 1.161905e-01
R9357 n2_8304_9921 n2_8304_9954 2.095238e-02
R9358 n2_8304_9954 n2_8304_9968 8.888889e-03
R9359 n2_8304_9968 n2_8304_10034 4.190476e-02
R9360 n2_8304_10034 n2_8304_10137 6.539683e-02
R9361 n2_8304_10137 n2_8304_10170 2.095238e-02
R9362 n2_8304_10170 n2_8304_10353 1.161905e-01
R9363 n2_8304_10353 n2_8304_10386 2.095238e-02
R9364 n2_8304_10386 n2_8304_10549 1.034921e-01
R9365 n2_8304_10549 n2_8304_10569 1.269841e-02
R9366 n2_8304_10569 n2_8304_10602 2.095238e-02
R9367 n2_8304_10602 n2_8304_10645 2.730159e-02
R9368 n2_8304_10645 n2_8304_10785 8.888889e-02
R9369 n2_8304_10785 n2_8304_10818 2.095238e-02
R9370 n2_8304_10818 n2_8304_11001 1.161905e-01
R9371 n2_8304_11001 n2_8304_11034 2.095238e-02
R9372 n2_8304_11034 n2_8304_11048 8.888889e-03
R9373 n2_8304_11048 n2_8304_11160 7.111111e-02
R9374 n2_8304_11160 n2_8304_11217 3.619048e-02
R9375 n2_8304_11217 n2_8304_11250 2.095238e-02
R9376 n2_8304_11250 n2_8304_11433 1.161905e-01
R9377 n2_8304_11433 n2_8304_11466 2.095238e-02
R9378 n2_8304_11865 n2_8304_11898 2.095238e-02
R9379 n2_8304_11898 n2_8304_12081 1.161905e-01
R9380 n2_8304_12081 n2_8304_12114 2.095238e-02
R9381 n2_8304_12114 n2_8304_12128 8.888889e-03
R9382 n2_8304_12128 n2_8304_12285 9.968254e-02
R9383 n2_8304_12285 n2_8304_12297 7.619048e-03
R9384 n2_8304_12297 n2_8304_12330 2.095238e-02
R9385 n2_8304_12330 n2_8304_12513 1.161905e-01
R9386 n2_8304_12513 n2_8304_12546 2.095238e-02
R9387 n2_8304_12546 n2_8304_12729 1.161905e-01
R9388 n2_8304_12729 n2_8304_12762 2.095238e-02
R9389 n2_8304_12762 n2_8304_12799 2.349206e-02
R9390 n2_8304_12799 n2_8304_12895 6.095238e-02
R9391 n2_8304_12895 n2_8304_12945 3.174603e-02
R9392 n2_8304_12945 n2_8304_12978 2.095238e-02
R9393 n2_8304_12978 n2_8304_13161 1.161905e-01
R9394 n2_8304_13161 n2_8304_13194 2.095238e-02
R9395 n2_8304_13194 n2_8304_13377 1.161905e-01
R9396 n2_8304_13377 n2_8304_13410 2.095238e-02
R9397 n2_8304_13410 n2_8304_13424 8.888889e-03
R9398 n2_8304_13424 n2_8304_13593 1.073016e-01
R9399 n2_8304_13593 n2_8304_13626 2.095238e-02
R9400 n2_8304_13626 n2_8304_13640 8.888889e-03
R9401 n2_8304_13640 n2_8304_13809 1.073016e-01
R9402 n2_8304_13809 n2_8304_13842 2.095238e-02
R9403 n2_8304_13842 n2_8304_13856 8.888889e-03
R9404 n2_8304_13856 n2_8304_13924 4.317460e-02
R9405 n2_8304_13924 n2_8304_14020 6.095238e-02
R9406 n2_8304_14020 n2_8304_14025 3.174603e-03
R9407 n2_8304_14025 n2_8304_14058 2.095238e-02
R9408 n2_8304_14058 n2_8304_14072 8.888889e-03
R9409 n2_8304_14072 n2_8304_14241 1.073016e-01
R9410 n2_8304_14241 n2_8304_14274 2.095238e-02
R9411 n2_8304_14274 n2_8304_14396 7.746032e-02
R9412 n2_8304_14396 n2_8304_14457 3.873016e-02
R9413 n2_8304_14457 n2_8304_14490 2.095238e-02
R9414 n2_8304_14490 n2_8304_14504 8.888889e-03
R9415 n2_8304_14504 n2_8304_14673 1.073016e-01
R9416 n2_8304_14673 n2_8304_14706 2.095238e-02
R9417 n2_8304_14706 n2_8304_14889 1.161905e-01
R9418 n2_8304_14889 n2_8304_14922 2.095238e-02
R9419 n2_8304_14922 n2_8304_15049 8.063492e-02
R9420 n2_8304_15049 n2_8304_15105 3.555556e-02
R9421 n2_8304_15105 n2_8304_15138 2.095238e-02
R9422 n2_8304_15138 n2_8304_15145 4.444444e-03
R9423 n2_8304_15145 n2_8304_15321 1.117460e-01
R9424 n2_8304_15321 n2_8304_15354 2.095238e-02
R9425 n2_8304_15354 n2_8304_15537 1.161905e-01
R9426 n2_8304_15537 n2_8304_15570 2.095238e-02
R9427 n2_8304_15570 n2_8304_15584 8.888889e-03
R9428 n2_8304_15584 n2_8304_15753 1.073016e-01
R9429 n2_8304_15753 n2_8304_15786 2.095238e-02
R9430 n2_8304_15786 n2_8304_15800 8.888889e-03
R9431 n2_8304_15800 n2_8304_15969 1.073016e-01
R9432 n2_8304_15969 n2_8304_16002 2.095238e-02
R9433 n2_8304_16002 n2_8304_16016 8.888889e-03
R9434 n2_8304_16016 n2_8304_16174 1.003175e-01
R9435 n2_8304_16174 n2_8304_16185 6.984127e-03
R9436 n2_8304_16185 n2_8304_16218 2.095238e-02
R9437 n2_8304_16218 n2_8304_16270 3.301587e-02
R9438 n2_8304_16270 n2_8304_16401 8.317460e-02
R9439 n2_8304_16401 n2_8304_16434 2.095238e-02
R9440 n2_8304_16434 n2_8304_16617 1.161905e-01
R9441 n2_8304_16617 n2_8304_16650 2.095238e-02
R9442 n2_8304_16650 n2_8304_16833 1.161905e-01
R9443 n2_8304_16833 n2_8304_16866 2.095238e-02
R9444 n2_8304_16866 n2_8304_17049 1.161905e-01
R9445 n2_8304_17049 n2_8304_17082 2.095238e-02
R9446 n2_8304_17082 n2_8304_17096 8.888889e-03
R9447 n2_8304_17096 n2_8304_17119 1.460317e-02
R9448 n2_8304_17119 n2_8304_17265 9.269841e-02
R9449 n2_8304_17265 n2_8304_17298 2.095238e-02
R9450 n2_8304_17298 n2_8304_17299 6.349206e-04
R9451 n2_8304_17299 n2_8304_17312 8.253968e-03
R9452 n2_8304_17312 n2_8304_17395 5.269841e-02
R9453 n2_8304_17395 n2_8304_17481 5.460317e-02
R9454 n2_8304_17481 n2_8304_17514 2.095238e-02
R9455 n2_8304_17514 n2_8304_17697 1.161905e-01
R9456 n2_8304_17697 n2_8304_17730 2.095238e-02
R9457 n2_8304_17730 n2_8304_17913 1.161905e-01
R9458 n2_8304_17913 n2_8304_17946 2.095238e-02
R9459 n2_8304_17946 n2_8304_18129 1.161905e-01
R9460 n2_8304_18129 n2_8304_18162 2.095238e-02
R9461 n2_8304_18162 n2_8304_18345 1.161905e-01
R9462 n2_8304_18345 n2_8304_18378 2.095238e-02
R9463 n2_8304_18378 n2_8304_18392 8.888889e-03
R9464 n2_8304_18392 n2_8304_18421 1.841270e-02
R9465 n2_8304_18421 n2_8304_18424 1.904762e-03
R9466 n2_8304_18424 n2_8304_18520 6.095238e-02
R9467 n2_8304_18520 n2_8304_18561 2.603175e-02
R9468 n2_8304_18561 n2_8304_18594 2.095238e-02
R9469 n2_8304_18594 n2_8304_18608 8.888889e-03
R9470 n2_8304_18608 n2_8304_18777 1.073016e-01
R9471 n2_8304_18777 n2_8304_18810 2.095238e-02
R9472 n2_8304_18810 n2_8304_18993 1.161905e-01
R9473 n2_8304_18993 n2_8304_19026 2.095238e-02
R9474 n2_8304_19026 n2_8304_19209 1.161905e-01
R9475 n2_8304_19209 n2_8304_19242 2.095238e-02
R9476 n2_8304_19242 n2_8304_19256 8.888889e-03
R9477 n2_8304_19256 n2_8304_19279 1.460317e-02
R9478 n2_8304_19279 n2_8304_19425 9.269841e-02
R9479 n2_8304_19425 n2_8304_19458 2.095238e-02
R9480 n2_8304_19458 n2_8304_19549 5.777778e-02
R9481 n2_8304_19549 n2_8304_19641 5.841270e-02
R9482 n2_8304_19641 n2_8304_19645 2.539683e-03
R9483 n2_8304_19645 n2_8304_19674 1.841270e-02
R9484 n2_8304_19674 n2_8304_19857 1.161905e-01
R9485 n2_8304_19857 n2_8304_19890 2.095238e-02
R9486 n2_8304_19890 n2_8304_20073 1.161905e-01
R9487 n2_8304_20073 n2_8304_20106 2.095238e-02
R9488 n2_8304_20106 n2_8304_20289 1.161905e-01
R9489 n2_8304_20289 n2_8304_20322 2.095238e-02
R9490 n2_8304_20322 n2_8304_20505 1.161905e-01
R9491 n2_8304_20505 n2_8304_20538 2.095238e-02
R9492 n2_8304_20538 n2_8304_20674 8.634921e-02
R9493 n2_8304_20674 n2_8304_20721 2.984127e-02
R9494 n2_8304_20721 n2_8304_20754 2.095238e-02
R9495 n2_8304_20754 n2_8304_20770 1.015873e-02
R9496 n2_8304_20770 n2_8304_20937 1.060317e-01
R9497 n2_8304_20937 n2_8304_20970 2.095238e-02
R9498 n2_8396_201 n2_8396_234 2.095238e-02
R9499 n2_8396_234 n2_8396_417 1.161905e-01
R9500 n2_8396_417 n2_8396_424 4.444444e-03
R9501 n2_8396_424 n2_8396_450 1.650794e-02
R9502 n2_8396_520 n2_8396_633 7.174603e-02
R9503 n2_8396_633 n2_8396_666 2.095238e-02
R9504 n2_8396_666 n2_8396_849 1.161905e-01
R9505 n2_8396_849 n2_8396_882 2.095238e-02
R9506 n2_8396_882 n2_8396_1065 1.161905e-01
R9507 n2_8396_1065 n2_8396_1098 2.095238e-02
R9508 n2_8396_1098 n2_8396_1281 1.161905e-01
R9509 n2_8396_1281 n2_8396_1314 2.095238e-02
R9510 n2_8396_1314 n2_8396_1497 1.161905e-01
R9511 n2_8396_1497 n2_8396_1530 2.095238e-02
R9512 n2_8396_1530 n2_8396_1549 1.206349e-02
R9513 n2_8396_1645 n2_8396_1713 4.317460e-02
R9514 n2_8396_1713 n2_8396_1746 2.095238e-02
R9515 n2_8396_1746 n2_8396_1760 8.888889e-03
R9516 n2_8396_1760 n2_8396_1783 1.460317e-02
R9517 n2_8396_1783 n2_8396_1929 9.269841e-02
R9518 n2_8396_1929 n2_8396_1962 2.095238e-02
R9519 n2_8396_1962 n2_8396_2145 1.161905e-01
R9520 n2_8396_2145 n2_8396_2178 2.095238e-02
R9521 n2_8396_2178 n2_8396_2361 1.161905e-01
R9522 n2_8396_2361 n2_8396_2394 2.095238e-02
R9523 n2_8396_2394 n2_8396_2408 8.888889e-03
R9524 n2_8396_2408 n2_8396_2577 1.073016e-01
R9525 n2_8396_2577 n2_8396_2610 2.095238e-02
R9526 n2_8396_2610 n2_8396_2674 4.063492e-02
R9527 n2_8396_2770 n2_8396_2793 1.460317e-02
R9528 n2_8396_2793 n2_8396_2826 2.095238e-02
R9529 n2_8396_2826 n2_8396_2840 8.888889e-03
R9530 n2_8396_2840 n2_8396_2863 1.460317e-02
R9531 n2_8396_2863 n2_8396_3009 9.269841e-02
R9532 n2_8396_3009 n2_8396_3042 2.095238e-02
R9533 n2_8396_3042 n2_8396_3225 1.161905e-01
R9534 n2_8396_3225 n2_8396_3258 2.095238e-02
R9535 n2_8396_3258 n2_8396_3441 1.161905e-01
R9536 n2_8396_3441 n2_8396_3474 2.095238e-02
R9537 n2_8396_3474 n2_8396_3488 8.888889e-03
R9538 n2_8396_3488 n2_8396_3657 1.073016e-01
R9539 n2_8396_3657 n2_8396_3690 2.095238e-02
R9540 n2_8396_3690 n2_8396_3799 6.920635e-02
R9541 n2_8396_3873 n2_8396_3895 1.396825e-02
R9542 n2_8396_3895 n2_8396_3906 6.984127e-03
R9543 n2_8396_3906 n2_8396_4089 1.161905e-01
R9544 n2_8396_4089 n2_8396_4122 2.095238e-02
R9545 n2_8396_4122 n2_8396_4136 8.888889e-03
R9546 n2_8396_4136 n2_8396_4305 1.073016e-01
R9547 n2_8396_4305 n2_8396_4338 2.095238e-02
R9548 n2_8396_4338 n2_8396_4521 1.161905e-01
R9549 n2_8396_4521 n2_8396_4554 2.095238e-02
R9550 n2_8396_4554 n2_8396_4568 8.888889e-03
R9551 n2_8396_4568 n2_8396_4737 1.073016e-01
R9552 n2_8396_4737 n2_8396_4770 2.095238e-02
R9553 n2_8396_4770 n2_8396_4924 9.777778e-02
R9554 n2_8396_4924 n2_8396_4953 1.841270e-02
R9555 n2_8396_5020 n2_8396_5169 9.460317e-02
R9556 n2_8396_5169 n2_8396_5202 2.095238e-02
R9557 n2_8396_5202 n2_8396_5216 8.888889e-03
R9558 n2_8396_5216 n2_8396_5239 1.460317e-02
R9559 n2_8396_5239 n2_8396_5385 9.269841e-02
R9560 n2_8396_5385 n2_8396_5418 2.095238e-02
R9561 n2_8396_5418 n2_8396_5432 8.888889e-03
R9562 n2_8396_5432 n2_8396_5455 1.460317e-02
R9563 n2_8396_5455 n2_8396_5601 9.269841e-02
R9564 n2_8396_5601 n2_8396_5634 2.095238e-02
R9565 n2_8396_5634 n2_8396_5817 1.161905e-01
R9566 n2_8396_5817 n2_8396_5850 2.095238e-02
R9567 n2_8396_5850 n2_8396_6033 1.161905e-01
R9568 n2_8396_6033 n2_8396_6049 1.015873e-02
R9569 n2_8396_6049 n2_8396_6066 1.079365e-02
R9570 n2_8396_6145 n2_8396_6249 6.603175e-02
R9571 n2_8396_6249 n2_8396_6282 2.095238e-02
R9572 n2_8396_6282 n2_8396_6465 1.161905e-01
R9573 n2_8396_6465 n2_8396_6498 2.095238e-02
R9574 n2_8396_6498 n2_8396_6512 8.888889e-03
R9575 n2_8396_6512 n2_8396_6535 1.460317e-02
R9576 n2_8396_6535 n2_8396_6681 9.269841e-02
R9577 n2_8396_6681 n2_8396_6714 2.095238e-02
R9578 n2_8396_6714 n2_8396_6897 1.161905e-01
R9579 n2_8396_6897 n2_8396_6930 2.095238e-02
R9580 n2_8396_6930 n2_8396_6944 8.888889e-03
R9581 n2_8396_6944 n2_8396_7113 1.073016e-01
R9582 n2_8396_7113 n2_8396_7146 2.095238e-02
R9583 n2_8396_7146 n2_8396_7160 8.888889e-03
R9584 n2_8396_7160 n2_8396_7174 8.888889e-03
R9585 n2_8396_7270 n2_8396_7329 3.746032e-02
R9586 n2_8396_7329 n2_8396_7362 2.095238e-02
R9587 n2_8396_7362 n2_8396_7376 8.888889e-03
R9588 n2_8396_7376 n2_8396_7545 1.073016e-01
R9589 n2_8396_7545 n2_8396_7578 2.095238e-02
R9590 n2_8396_7578 n2_8396_7761 1.161905e-01
R9591 n2_8396_7761 n2_8396_7794 2.095238e-02
R9592 n2_8396_7794 n2_8396_7808 8.888889e-03
R9593 n2_8396_7808 n2_8396_7977 1.073016e-01
R9594 n2_8396_7977 n2_8396_8010 2.095238e-02
R9595 n2_8396_8010 n2_8396_8193 1.161905e-01
R9596 n2_8396_8193 n2_8396_8226 2.095238e-02
R9597 n2_8396_8226 n2_8396_8299 4.634921e-02
R9598 n2_8396_12895 n2_8396_12945 3.174603e-02
R9599 n2_8396_12945 n2_8396_12978 2.095238e-02
R9600 n2_8396_12978 n2_8396_13161 1.161905e-01
R9601 n2_8396_13161 n2_8396_13194 2.095238e-02
R9602 n2_8396_13194 n2_8396_13377 1.161905e-01
R9603 n2_8396_13377 n2_8396_13410 2.095238e-02
R9604 n2_8396_13410 n2_8396_13424 8.888889e-03
R9605 n2_8396_13424 n2_8396_13593 1.073016e-01
R9606 n2_8396_13593 n2_8396_13626 2.095238e-02
R9607 n2_8396_13626 n2_8396_13640 8.888889e-03
R9608 n2_8396_13640 n2_8396_13809 1.073016e-01
R9609 n2_8396_13809 n2_8396_13842 2.095238e-02
R9610 n2_8396_13842 n2_8396_13856 8.888889e-03
R9611 n2_8396_13856 n2_8396_13924 4.317460e-02
R9612 n2_8396_14020 n2_8396_14025 3.174603e-03
R9613 n2_8396_14025 n2_8396_14058 2.095238e-02
R9614 n2_8396_14058 n2_8396_14072 8.888889e-03
R9615 n2_8396_14072 n2_8396_14241 1.073016e-01
R9616 n2_8396_14241 n2_8396_14274 2.095238e-02
R9617 n2_8396_14274 n2_8396_14396 7.746032e-02
R9618 n2_8396_14396 n2_8396_14457 3.873016e-02
R9619 n2_8396_14457 n2_8396_14490 2.095238e-02
R9620 n2_8396_14490 n2_8396_14504 8.888889e-03
R9621 n2_8396_14504 n2_8396_14673 1.073016e-01
R9622 n2_8396_14673 n2_8396_14706 2.095238e-02
R9623 n2_8396_14706 n2_8396_14889 1.161905e-01
R9624 n2_8396_14889 n2_8396_14922 2.095238e-02
R9625 n2_8396_14922 n2_8396_15049 8.063492e-02
R9626 n2_8396_15138 n2_8396_15145 4.444444e-03
R9627 n2_8396_15145 n2_8396_15321 1.117460e-01
R9628 n2_8396_15321 n2_8396_15354 2.095238e-02
R9629 n2_8396_15354 n2_8396_15537 1.161905e-01
R9630 n2_8396_15537 n2_8396_15570 2.095238e-02
R9631 n2_8396_15570 n2_8396_15584 8.888889e-03
R9632 n2_8396_15584 n2_8396_15753 1.073016e-01
R9633 n2_8396_15753 n2_8396_15786 2.095238e-02
R9634 n2_8396_15786 n2_8396_15800 8.888889e-03
R9635 n2_8396_15800 n2_8396_15969 1.073016e-01
R9636 n2_8396_15969 n2_8396_16002 2.095238e-02
R9637 n2_8396_16002 n2_8396_16016 8.888889e-03
R9638 n2_8396_16016 n2_8396_16174 1.003175e-01
R9639 n2_8396_16174 n2_8396_16185 6.984127e-03
R9640 n2_8396_16270 n2_8396_16401 8.317460e-02
R9641 n2_8396_16401 n2_8396_16434 2.095238e-02
R9642 n2_8396_16434 n2_8396_16617 1.161905e-01
R9643 n2_8396_16617 n2_8396_16650 2.095238e-02
R9644 n2_8396_16650 n2_8396_16833 1.161905e-01
R9645 n2_8396_16833 n2_8396_16866 2.095238e-02
R9646 n2_8396_16866 n2_8396_17049 1.161905e-01
R9647 n2_8396_17049 n2_8396_17082 2.095238e-02
R9648 n2_8396_17082 n2_8396_17096 8.888889e-03
R9649 n2_8396_17096 n2_8396_17119 1.460317e-02
R9650 n2_8396_17119 n2_8396_17265 9.269841e-02
R9651 n2_8396_17265 n2_8396_17298 2.095238e-02
R9652 n2_8396_17298 n2_8396_17299 6.349206e-04
R9653 n2_8396_17299 n2_8396_17312 8.253968e-03
R9654 n2_8396_17395 n2_8396_17481 5.460317e-02
R9655 n2_8396_17481 n2_8396_17514 2.095238e-02
R9656 n2_8396_17514 n2_8396_17697 1.161905e-01
R9657 n2_8396_17697 n2_8396_17730 2.095238e-02
R9658 n2_8396_17730 n2_8396_17913 1.161905e-01
R9659 n2_8396_17913 n2_8396_17946 2.095238e-02
R9660 n2_8396_17946 n2_8396_18129 1.161905e-01
R9661 n2_8396_18129 n2_8396_18162 2.095238e-02
R9662 n2_8396_18162 n2_8396_18345 1.161905e-01
R9663 n2_8396_18345 n2_8396_18378 2.095238e-02
R9664 n2_8396_18378 n2_8396_18392 8.888889e-03
R9665 n2_8396_18392 n2_8396_18421 1.841270e-02
R9666 n2_8396_18421 n2_8396_18424 1.904762e-03
R9667 n2_8396_18520 n2_8396_18561 2.603175e-02
R9668 n2_8396_18561 n2_8396_18594 2.095238e-02
R9669 n2_8396_18594 n2_8396_18608 8.888889e-03
R9670 n2_8396_18608 n2_8396_18777 1.073016e-01
R9671 n2_8396_18777 n2_8396_18810 2.095238e-02
R9672 n2_8396_18810 n2_8396_18993 1.161905e-01
R9673 n2_8396_18993 n2_8396_19026 2.095238e-02
R9674 n2_8396_19026 n2_8396_19209 1.161905e-01
R9675 n2_8396_19209 n2_8396_19242 2.095238e-02
R9676 n2_8396_19242 n2_8396_19256 8.888889e-03
R9677 n2_8396_19256 n2_8396_19279 1.460317e-02
R9678 n2_8396_19279 n2_8396_19425 9.269841e-02
R9679 n2_8396_19425 n2_8396_19458 2.095238e-02
R9680 n2_8396_19458 n2_8396_19549 5.777778e-02
R9681 n2_8396_19641 n2_8396_19645 2.539683e-03
R9682 n2_8396_19645 n2_8396_19674 1.841270e-02
R9683 n2_8396_19674 n2_8396_19857 1.161905e-01
R9684 n2_8396_19857 n2_8396_19890 2.095238e-02
R9685 n2_8396_19890 n2_8396_20073 1.161905e-01
R9686 n2_8396_20073 n2_8396_20106 2.095238e-02
R9687 n2_8396_20106 n2_8396_20289 1.161905e-01
R9688 n2_8396_20289 n2_8396_20322 2.095238e-02
R9689 n2_8396_20322 n2_8396_20505 1.161905e-01
R9690 n2_8396_20505 n2_8396_20538 2.095238e-02
R9691 n2_8396_20538 n2_8396_20674 8.634921e-02
R9692 n2_8396_20754 n2_8396_20770 1.015873e-02
R9693 n2_8396_20770 n2_8396_20937 1.060317e-01
R9694 n2_8396_20937 n2_8396_20970 2.095238e-02
R9695 n2_9241_9489 n2_9241_9522 2.095238e-02
R9696 n2_9241_9522 n2_9241_9705 1.161905e-01
R9697 n2_9241_9705 n2_9241_9738 2.095238e-02
R9698 n2_9241_9738 n2_9241_9921 1.161905e-01
R9699 n2_9241_9921 n2_9241_9954 2.095238e-02
R9700 n2_9241_9954 n2_9241_10034 5.079365e-02
R9701 n2_9241_10034 n2_9241_10137 6.539683e-02
R9702 n2_9241_10137 n2_9241_10170 2.095238e-02
R9703 n2_9241_10170 n2_9241_10353 1.161905e-01
R9704 n2_9241_10353 n2_9241_10386 2.095238e-02
R9705 n2_9241_10386 n2_9241_10549 1.034921e-01
R9706 n2_9241_10549 n2_9241_10569 1.269841e-02
R9707 n2_9241_10645 n2_9241_10785 8.888889e-02
R9708 n2_9241_10785 n2_9241_10818 2.095238e-02
R9709 n2_9241_10818 n2_9241_11001 1.161905e-01
R9710 n2_9241_11001 n2_9241_11034 2.095238e-02
R9711 n2_9241_11034 n2_9241_11160 8.000000e-02
R9712 n2_9241_11160 n2_9241_11217 3.619048e-02
R9713 n2_9241_11217 n2_9241_11250 2.095238e-02
R9714 n2_9241_11250 n2_9241_11433 1.161905e-01
R9715 n2_9241_11433 n2_9241_11466 2.095238e-02
R9716 n2_9241_11466 n2_9241_11649 1.161905e-01
R9717 n2_9241_11649 n2_9241_11682 2.095238e-02
R9718 n2_9241_10549 n2_9380_10549 8.825397e-02
R9719 n2_9380_10549 n2_9429_10549 3.111111e-02
R9720 n2_9241_10645 n2_9380_10645 8.825397e-02
R9721 n2_9380_10645 n2_9429_10645 3.111111e-02
R9722 n2_9429_9705 n2_9429_9738 2.095238e-02
R9723 n2_9429_9738 n2_9429_9921 1.161905e-01
R9724 n2_9429_9921 n2_9429_9954 2.095238e-02
R9725 n2_9429_9954 n2_9429_10137 1.161905e-01
R9726 n2_9429_10137 n2_9429_10170 2.095238e-02
R9727 n2_9429_10170 n2_9429_10353 1.161905e-01
R9728 n2_9429_10353 n2_9429_10386 2.095238e-02
R9729 n2_9429_10386 n2_9429_10549 1.034921e-01
R9730 n2_9429_10549 n2_9429_10569 1.269841e-02
R9731 n2_9429_10569 n2_9429_10602 2.095238e-02
R9732 n2_9429_10602 n2_9429_10645 2.730159e-02
R9733 n2_9429_10645 n2_9429_10785 8.888889e-02
R9734 n2_9429_10785 n2_9429_10818 2.095238e-02
R9735 n2_9429_10818 n2_9429_11001 1.161905e-01
R9736 n2_9429_11001 n2_9429_11034 2.095238e-02
R9737 n2_9429_11034 n2_9429_11217 1.161905e-01
R9738 n2_9429_11217 n2_9429_11250 2.095238e-02
R9739 n2_9429_11250 n2_9429_11433 1.161905e-01
R9740 n2_9429_11433 n2_9429_11466 2.095238e-02
R9741 n2_10366_201 n2_10366_234 2.095238e-02
R9742 n2_10366_234 n2_10366_417 1.161905e-01
R9743 n2_10366_417 n2_10366_424 4.444444e-03
R9744 n2_10366_424 n2_10366_450 1.650794e-02
R9745 n2_10366_520 n2_10366_633 7.174603e-02
R9746 n2_10366_633 n2_10366_666 2.095238e-02
R9747 n2_10366_666 n2_10366_849 1.161905e-01
R9748 n2_10366_849 n2_10366_882 2.095238e-02
R9749 n2_10366_882 n2_10366_1065 1.161905e-01
R9750 n2_10366_1065 n2_10366_1098 2.095238e-02
R9751 n2_10366_1098 n2_10366_1281 1.161905e-01
R9752 n2_10366_1281 n2_10366_1314 2.095238e-02
R9753 n2_10366_1314 n2_10366_1497 1.161905e-01
R9754 n2_10366_1497 n2_10366_1530 2.095238e-02
R9755 n2_10366_1530 n2_10366_1549 1.206349e-02
R9756 n2_10366_1645 n2_10366_1713 4.317460e-02
R9757 n2_10366_1713 n2_10366_1746 2.095238e-02
R9758 n2_10366_1746 n2_10366_1760 8.888889e-03
R9759 n2_10366_1760 n2_10366_1783 1.460317e-02
R9760 n2_10366_1783 n2_10366_1929 9.269841e-02
R9761 n2_10366_1929 n2_10366_1962 2.095238e-02
R9762 n2_10366_1962 n2_10366_2145 1.161905e-01
R9763 n2_10366_2145 n2_10366_2178 2.095238e-02
R9764 n2_10366_2178 n2_10366_2361 1.161905e-01
R9765 n2_10366_2361 n2_10366_2394 2.095238e-02
R9766 n2_10366_2394 n2_10366_2408 8.888889e-03
R9767 n2_10366_2408 n2_10366_2577 1.073016e-01
R9768 n2_10366_2577 n2_10366_2610 2.095238e-02
R9769 n2_10366_2610 n2_10366_2647 2.349206e-02
R9770 n2_10366_2647 n2_10366_2674 1.714286e-02
R9771 n2_10366_2770 n2_10366_2793 1.460317e-02
R9772 n2_10366_2793 n2_10366_2826 2.095238e-02
R9773 n2_10366_2826 n2_10366_2840 8.888889e-03
R9774 n2_10366_2840 n2_10366_2863 1.460317e-02
R9775 n2_10366_2863 n2_10366_3009 9.269841e-02
R9776 n2_10366_3009 n2_10366_3042 2.095238e-02
R9777 n2_10366_3042 n2_10366_3225 1.161905e-01
R9778 n2_10366_3225 n2_10366_3258 2.095238e-02
R9779 n2_10366_3258 n2_10366_3441 1.161905e-01
R9780 n2_10366_3441 n2_10366_3474 2.095238e-02
R9781 n2_10366_3474 n2_10366_3488 8.888889e-03
R9782 n2_10366_3488 n2_10366_3511 1.460317e-02
R9783 n2_10366_3511 n2_10366_3657 9.269841e-02
R9784 n2_10366_3657 n2_10366_3690 2.095238e-02
R9785 n2_10366_3690 n2_10366_3799 6.920635e-02
R9786 n2_10366_3873 n2_10366_3895 1.396825e-02
R9787 n2_10366_3895 n2_10366_3906 6.984127e-03
R9788 n2_10366_3906 n2_10366_4089 1.161905e-01
R9789 n2_10366_4089 n2_10366_4122 2.095238e-02
R9790 n2_10366_4122 n2_10366_4136 8.888889e-03
R9791 n2_10366_4136 n2_10366_4159 1.460317e-02
R9792 n2_10366_4159 n2_10366_4305 9.269841e-02
R9793 n2_10366_4305 n2_10366_4338 2.095238e-02
R9794 n2_10366_4338 n2_10366_4521 1.161905e-01
R9795 n2_10366_4521 n2_10366_4554 2.095238e-02
R9796 n2_10366_4554 n2_10366_4568 8.888889e-03
R9797 n2_10366_4568 n2_10366_4591 1.460317e-02
R9798 n2_10366_4591 n2_10366_4737 9.269841e-02
R9799 n2_10366_4737 n2_10366_4770 2.095238e-02
R9800 n2_10366_4770 n2_10366_4924 9.777778e-02
R9801 n2_10366_4924 n2_10366_4953 1.841270e-02
R9802 n2_10366_5020 n2_10366_5169 9.460317e-02
R9803 n2_10366_5169 n2_10366_5202 2.095238e-02
R9804 n2_10366_5202 n2_10366_5239 2.349206e-02
R9805 n2_10366_5239 n2_10366_5385 9.269841e-02
R9806 n2_10366_5385 n2_10366_5418 2.095238e-02
R9807 n2_10366_5418 n2_10366_5432 8.888889e-03
R9808 n2_10366_5432 n2_10366_5455 1.460317e-02
R9809 n2_10366_5455 n2_10366_5601 9.269841e-02
R9810 n2_10366_5601 n2_10366_5634 2.095238e-02
R9811 n2_10366_5634 n2_10366_5817 1.161905e-01
R9812 n2_10366_5817 n2_10366_5850 2.095238e-02
R9813 n2_10366_5850 n2_10366_6033 1.161905e-01
R9814 n2_10366_6033 n2_10366_6049 1.015873e-02
R9815 n2_10366_6049 n2_10366_6066 1.079365e-02
R9816 n2_10366_6145 n2_10366_6249 6.603175e-02
R9817 n2_10366_6249 n2_10366_6282 2.095238e-02
R9818 n2_10366_6282 n2_10366_6465 1.161905e-01
R9819 n2_10366_6465 n2_10366_6498 2.095238e-02
R9820 n2_10366_6498 n2_10366_6512 8.888889e-03
R9821 n2_10366_6512 n2_10366_6535 1.460317e-02
R9822 n2_10366_6535 n2_10366_6681 9.269841e-02
R9823 n2_10366_6681 n2_10366_6714 2.095238e-02
R9824 n2_10366_6714 n2_10366_6751 2.349206e-02
R9825 n2_10366_6751 n2_10366_6897 9.269841e-02
R9826 n2_10366_6897 n2_10366_6930 2.095238e-02
R9827 n2_10366_6930 n2_10366_6944 8.888889e-03
R9828 n2_10366_6944 n2_10366_6967 1.460317e-02
R9829 n2_10366_6967 n2_10366_7113 9.269841e-02
R9830 n2_10366_7113 n2_10366_7146 2.095238e-02
R9831 n2_10366_7146 n2_10366_7160 8.888889e-03
R9832 n2_10366_7160 n2_10366_7174 8.888889e-03
R9833 n2_10366_7174 n2_10366_7178 2.539683e-03
R9834 n2_10366_7270 n2_10366_7329 3.746032e-02
R9835 n2_10366_7329 n2_10366_7362 2.095238e-02
R9836 n2_10366_7362 n2_10366_7376 8.888889e-03
R9837 n2_10366_7376 n2_10366_7399 1.460317e-02
R9838 n2_10366_7399 n2_10366_7545 9.269841e-02
R9839 n2_10366_7545 n2_10366_7578 2.095238e-02
R9840 n2_10366_7578 n2_10366_7761 1.161905e-01
R9841 n2_10366_7761 n2_10366_7794 2.095238e-02
R9842 n2_10366_7794 n2_10366_7977 1.161905e-01
R9843 n2_10366_7977 n2_10366_8010 2.095238e-02
R9844 n2_10366_8010 n2_10366_8193 1.161905e-01
R9845 n2_10366_8193 n2_10366_8226 2.095238e-02
R9846 n2_10366_8226 n2_10366_8299 4.634921e-02
R9847 n2_10366_8395 n2_10366_8409 8.888889e-03
R9848 n2_10366_8409 n2_10366_8442 2.095238e-02
R9849 n2_10366_8442 n2_10366_8613 1.085714e-01
R9850 n2_10366_8613 n2_10366_8625 7.619048e-03
R9851 n2_10366_8625 n2_10366_8658 2.095238e-02
R9852 n2_10366_8658 n2_10366_8841 1.161905e-01
R9853 n2_10366_8841 n2_10366_8874 2.095238e-02
R9854 n2_10366_8874 n2_10366_9057 1.161905e-01
R9855 n2_10366_9057 n2_10366_9090 2.095238e-02
R9856 n2_10366_9090 n2_10366_9190 6.349206e-02
R9857 n2_10366_9190 n2_10366_9273 5.269841e-02
R9858 n2_10366_9273 n2_10366_9306 2.095238e-02
R9859 n2_10366_9306 n2_10366_9424 7.492063e-02
R9860 n2_10366_9489 n2_10366_9520 1.968254e-02
R9861 n2_10366_9520 n2_10366_9522 1.269841e-03
R9862 n2_10366_9522 n2_10366_9705 1.161905e-01
R9863 n2_10366_9705 n2_10366_9738 2.095238e-02
R9864 n2_10366_9738 n2_10366_9921 1.161905e-01
R9865 n2_10366_9921 n2_10366_9954 2.095238e-02
R9866 n2_10366_9954 n2_10366_10137 1.161905e-01
R9867 n2_10366_10137 n2_10366_10170 2.095238e-02
R9868 n2_10366_10170 n2_10366_10353 1.161905e-01
R9869 n2_10366_10353 n2_10366_10386 2.095238e-02
R9870 n2_10366_10386 n2_10366_10549 1.034921e-01
R9871 n2_10366_10549 n2_10366_10557 5.079365e-03
R9872 n2_10366_10557 n2_10366_10569 7.619048e-03
R9873 n2_10366_10645 n2_10366_10785 8.888889e-02
R9874 n2_10366_10785 n2_10366_10818 2.095238e-02
R9875 n2_10366_10818 n2_10366_11001 1.161905e-01
R9876 n2_10366_11001 n2_10366_11034 2.095238e-02
R9877 n2_10366_11034 n2_10366_11217 1.161905e-01
R9878 n2_10366_11217 n2_10366_11250 2.095238e-02
R9879 n2_10366_11250 n2_10366_11433 1.161905e-01
R9880 n2_10366_11433 n2_10366_11466 2.095238e-02
R9881 n2_10366_11466 n2_10366_11649 1.161905e-01
R9882 n2_10366_11649 n2_10366_11674 1.587302e-02
R9883 n2_10366_11674 n2_10366_11682 5.079365e-03
R9884 n2_10366_11770 n2_10366_11865 6.031746e-02
R9885 n2_10366_11865 n2_10366_11898 2.095238e-02
R9886 n2_10366_11898 n2_10366_12004 6.730159e-02
R9887 n2_10366_12004 n2_10366_12081 4.888889e-02
R9888 n2_10366_12081 n2_10366_12114 2.095238e-02
R9889 n2_10366_12114 n2_10366_12297 1.161905e-01
R9890 n2_10366_12297 n2_10366_12330 2.095238e-02
R9891 n2_10366_12330 n2_10366_12513 1.161905e-01
R9892 n2_10366_12513 n2_10366_12546 2.095238e-02
R9893 n2_10366_12546 n2_10366_12566 1.269841e-02
R9894 n2_10366_12566 n2_10366_12729 1.034921e-01
R9895 n2_10366_12729 n2_10366_12762 2.095238e-02
R9896 n2_10366_12762 n2_10366_12799 2.349206e-02
R9897 n2_10366_12895 n2_10366_12945 3.174603e-02
R9898 n2_10366_12945 n2_10366_12978 2.095238e-02
R9899 n2_10366_12978 n2_10366_13161 1.161905e-01
R9900 n2_10366_13161 n2_10366_13194 2.095238e-02
R9901 n2_10366_13194 n2_10366_13377 1.161905e-01
R9902 n2_10366_13377 n2_10366_13410 2.095238e-02
R9903 n2_10366_13410 n2_10366_13593 1.161905e-01
R9904 n2_10366_13593 n2_10366_13626 2.095238e-02
R9905 n2_10366_13626 n2_10366_13640 8.888889e-03
R9906 n2_10366_13640 n2_10366_13663 1.460317e-02
R9907 n2_10366_13663 n2_10366_13809 9.269841e-02
R9908 n2_10366_13809 n2_10366_13842 2.095238e-02
R9909 n2_10366_13842 n2_10366_13856 8.888889e-03
R9910 n2_10366_13856 n2_10366_13879 1.460317e-02
R9911 n2_10366_13879 n2_10366_13924 2.857143e-02
R9912 n2_10366_14020 n2_10366_14025 3.174603e-03
R9913 n2_10366_14025 n2_10366_14058 2.095238e-02
R9914 n2_10366_14058 n2_10366_14072 8.888889e-03
R9915 n2_10366_14072 n2_10366_14079 4.444444e-03
R9916 n2_10366_14079 n2_10366_14241 1.028571e-01
R9917 n2_10366_14241 n2_10366_14274 2.095238e-02
R9918 n2_10366_14274 n2_10366_14457 1.161905e-01
R9919 n2_10366_14457 n2_10366_14490 2.095238e-02
R9920 n2_10366_14490 n2_10366_14504 8.888889e-03
R9921 n2_10366_14504 n2_10366_14673 1.073016e-01
R9922 n2_10366_14673 n2_10366_14706 2.095238e-02
R9923 n2_10366_14706 n2_10366_14889 1.161905e-01
R9924 n2_10366_14889 n2_10366_14922 2.095238e-02
R9925 n2_10366_14922 n2_10366_15049 8.063492e-02
R9926 n2_10366_15138 n2_10366_15145 4.444444e-03
R9927 n2_10366_15145 n2_10366_15321 1.117460e-01
R9928 n2_10366_15321 n2_10366_15354 2.095238e-02
R9929 n2_10366_15354 n2_10366_15537 1.161905e-01
R9930 n2_10366_15537 n2_10366_15570 2.095238e-02
R9931 n2_10366_15570 n2_10366_15584 8.888889e-03
R9932 n2_10366_15584 n2_10366_15753 1.073016e-01
R9933 n2_10366_15753 n2_10366_15786 2.095238e-02
R9934 n2_10366_15786 n2_10366_15800 8.888889e-03
R9935 n2_10366_15800 n2_10366_15823 1.460317e-02
R9936 n2_10366_15823 n2_10366_15969 9.269841e-02
R9937 n2_10366_15969 n2_10366_16002 2.095238e-02
R9938 n2_10366_16002 n2_10366_16016 8.888889e-03
R9939 n2_10366_16016 n2_10366_16174 1.003175e-01
R9940 n2_10366_16174 n2_10366_16185 6.984127e-03
R9941 n2_10366_16270 n2_10366_16401 8.317460e-02
R9942 n2_10366_16401 n2_10366_16434 2.095238e-02
R9943 n2_10366_16434 n2_10366_16617 1.161905e-01
R9944 n2_10366_16617 n2_10366_16650 2.095238e-02
R9945 n2_10366_16650 n2_10366_16833 1.161905e-01
R9946 n2_10366_16833 n2_10366_16866 2.095238e-02
R9947 n2_10366_16866 n2_10366_17049 1.161905e-01
R9948 n2_10366_17049 n2_10366_17082 2.095238e-02
R9949 n2_10366_17082 n2_10366_17096 8.888889e-03
R9950 n2_10366_17096 n2_10366_17103 4.444444e-03
R9951 n2_10366_17103 n2_10366_17119 1.015873e-02
R9952 n2_10366_17119 n2_10366_17265 9.269841e-02
R9953 n2_10366_17265 n2_10366_17298 2.095238e-02
R9954 n2_10366_17298 n2_10366_17299 6.349206e-04
R9955 n2_10366_17299 n2_10366_17312 8.253968e-03
R9956 n2_10366_17395 n2_10366_17481 5.460317e-02
R9957 n2_10366_17481 n2_10366_17514 2.095238e-02
R9958 n2_10366_17514 n2_10366_17697 1.161905e-01
R9959 n2_10366_17697 n2_10366_17730 2.095238e-02
R9960 n2_10366_17730 n2_10366_17913 1.161905e-01
R9961 n2_10366_17913 n2_10366_17946 2.095238e-02
R9962 n2_10366_17946 n2_10366_18129 1.161905e-01
R9963 n2_10366_18129 n2_10366_18162 2.095238e-02
R9964 n2_10366_18162 n2_10366_18345 1.161905e-01
R9965 n2_10366_18345 n2_10366_18378 2.095238e-02
R9966 n2_10366_18378 n2_10366_18392 8.888889e-03
R9967 n2_10366_18392 n2_10366_18424 2.031746e-02
R9968 n2_10366_18520 n2_10366_18561 2.603175e-02
R9969 n2_10366_18561 n2_10366_18594 2.095238e-02
R9970 n2_10366_18594 n2_10366_18608 8.888889e-03
R9971 n2_10366_18608 n2_10366_18777 1.073016e-01
R9972 n2_10366_18777 n2_10366_18810 2.095238e-02
R9973 n2_10366_18810 n2_10366_18993 1.161905e-01
R9974 n2_10366_18993 n2_10366_19026 2.095238e-02
R9975 n2_10366_19026 n2_10366_19209 1.161905e-01
R9976 n2_10366_19209 n2_10366_19242 2.095238e-02
R9977 n2_10366_19242 n2_10366_19256 8.888889e-03
R9978 n2_10366_19256 n2_10366_19425 1.073016e-01
R9979 n2_10366_19425 n2_10366_19458 2.095238e-02
R9980 n2_10366_19458 n2_10366_19549 5.777778e-02
R9981 n2_10366_19641 n2_10366_19645 2.539683e-03
R9982 n2_10366_19645 n2_10366_19674 1.841270e-02
R9983 n2_10366_19674 n2_10366_19857 1.161905e-01
R9984 n2_10366_19857 n2_10366_19890 2.095238e-02
R9985 n2_10366_19890 n2_10366_20073 1.161905e-01
R9986 n2_10366_20073 n2_10366_20106 2.095238e-02
R9987 n2_10366_20106 n2_10366_20289 1.161905e-01
R9988 n2_10366_20289 n2_10366_20322 2.095238e-02
R9989 n2_10366_20322 n2_10366_20505 1.161905e-01
R9990 n2_10366_20505 n2_10366_20538 2.095238e-02
R9991 n2_10366_20538 n2_10366_20674 8.634921e-02
R9992 n2_10366_20754 n2_10366_20770 1.015873e-02
R9993 n2_10366_20770 n2_10366_20937 1.060317e-01
R9994 n2_10366_20937 n2_10366_20970 2.095238e-02
R9995 n2_10366_424 n2_10458_424 5.841270e-02
R9996 n2_10458_424 n2_10505_424 2.984127e-02
R9997 n2_10505_424 n2_10554_424 3.111111e-02
R9998 n2_10554_424 n2_10646_424 5.841270e-02
R9999 n2_10366_520 n2_10458_520 5.841270e-02
R10000 n2_10458_520 n2_10505_520 2.984127e-02
R10001 n2_10505_520 n2_10554_520 3.111111e-02
R10002 n2_10554_520 n2_10646_520 5.841270e-02
R10003 n2_10366_1549 n2_10458_1549 5.841270e-02
R10004 n2_10458_1549 n2_10505_1549 2.984127e-02
R10005 n2_10505_1549 n2_10554_1549 3.111111e-02
R10006 n2_10554_1549 n2_10646_1549 5.841270e-02
R10007 n2_10366_1645 n2_10458_1645 5.841270e-02
R10008 n2_10458_1645 n2_10505_1645 2.984127e-02
R10009 n2_10505_1645 n2_10554_1645 3.111111e-02
R10010 n2_10554_1645 n2_10646_1645 5.841270e-02
R10011 n2_10366_2674 n2_10458_2674 5.841270e-02
R10012 n2_10458_2674 n2_10505_2674 2.984127e-02
R10013 n2_10505_2674 n2_10554_2674 3.111111e-02
R10014 n2_10554_2674 n2_10646_2674 5.841270e-02
R10015 n2_10366_2770 n2_10458_2770 5.841270e-02
R10016 n2_10458_2770 n2_10505_2770 2.984127e-02
R10017 n2_10505_2770 n2_10554_2770 3.111111e-02
R10018 n2_10554_2770 n2_10646_2770 5.841270e-02
R10019 n2_10366_3799 n2_10458_3799 5.841270e-02
R10020 n2_10458_3799 n2_10505_3799 2.984127e-02
R10021 n2_10505_3799 n2_10554_3799 3.111111e-02
R10022 n2_10554_3799 n2_10646_3799 5.841270e-02
R10023 n2_10366_3895 n2_10458_3895 5.841270e-02
R10024 n2_10458_3895 n2_10505_3895 2.984127e-02
R10025 n2_10505_3895 n2_10554_3895 3.111111e-02
R10026 n2_10554_3895 n2_10646_3895 5.841270e-02
R10027 n2_10366_4924 n2_10458_4924 5.841270e-02
R10028 n2_10458_4924 n2_10505_4924 2.984127e-02
R10029 n2_10505_4924 n2_10554_4924 3.111111e-02
R10030 n2_10554_4924 n2_10646_4924 5.841270e-02
R10031 n2_10366_5020 n2_10458_5020 5.841270e-02
R10032 n2_10458_5020 n2_10505_5020 2.984127e-02
R10033 n2_10505_5020 n2_10554_5020 3.111111e-02
R10034 n2_10554_5020 n2_10646_5020 5.841270e-02
R10035 n2_10366_6049 n2_10458_6049 5.841270e-02
R10036 n2_10458_6049 n2_10505_6049 2.984127e-02
R10037 n2_10505_6049 n2_10554_6049 3.111111e-02
R10038 n2_10554_6049 n2_10646_6049 5.841270e-02
R10039 n2_10366_6145 n2_10458_6145 5.841270e-02
R10040 n2_10458_6145 n2_10505_6145 2.984127e-02
R10041 n2_10505_6145 n2_10554_6145 3.111111e-02
R10042 n2_10554_6145 n2_10646_6145 5.841270e-02
R10043 n2_10366_7174 n2_10458_7174 5.841270e-02
R10044 n2_10458_7174 n2_10505_7174 2.984127e-02
R10045 n2_10505_7174 n2_10554_7174 3.111111e-02
R10046 n2_10554_7174 n2_10646_7174 5.841270e-02
R10047 n2_10366_7270 n2_10458_7270 5.841270e-02
R10048 n2_10458_7270 n2_10505_7270 2.984127e-02
R10049 n2_10505_7270 n2_10554_7270 3.111111e-02
R10050 n2_10554_7270 n2_10646_7270 5.841270e-02
R10051 n2_10366_8299 n2_10458_8299 5.841270e-02
R10052 n2_10458_8299 n2_10505_8299 2.984127e-02
R10053 n2_10505_8299 n2_10554_8299 3.111111e-02
R10054 n2_10554_8299 n2_10646_8299 5.841270e-02
R10055 n2_10366_8395 n2_10458_8395 5.841270e-02
R10056 n2_10458_8395 n2_10505_8395 2.984127e-02
R10057 n2_10505_8395 n2_10554_8395 3.111111e-02
R10058 n2_10554_8395 n2_10646_8395 5.841270e-02
R10059 n2_10366_9424 n2_10458_9424 5.841270e-02
R10060 n2_10458_9424 n2_10505_9424 2.984127e-02
R10061 n2_10505_9424 n2_10554_9424 3.111111e-02
R10062 n2_10554_9424 n2_10646_9424 5.841270e-02
R10063 n2_10366_9520 n2_10458_9520 5.841270e-02
R10064 n2_10458_9520 n2_10505_9520 2.984127e-02
R10065 n2_10505_9520 n2_10554_9520 3.111111e-02
R10066 n2_10554_9520 n2_10646_9520 5.841270e-02
R10067 n2_10366_10549 n2_10458_10549 5.841270e-02
R10068 n2_10458_10549 n2_10505_10549 2.984127e-02
R10069 n2_10505_10549 n2_10554_10549 3.111111e-02
R10070 n2_10554_10549 n2_10646_10549 5.841270e-02
R10071 n2_10366_10645 n2_10458_10645 5.841270e-02
R10072 n2_10458_10645 n2_10505_10645 2.984127e-02
R10073 n2_10505_10645 n2_10554_10645 3.111111e-02
R10074 n2_10554_10645 n2_10646_10645 5.841270e-02
R10075 n2_10366_11674 n2_10458_11674 5.841270e-02
R10076 n2_10458_11674 n2_10505_11674 2.984127e-02
R10077 n2_10505_11674 n2_10554_11674 3.111111e-02
R10078 n2_10554_11674 n2_10646_11674 5.841270e-02
R10079 n2_10366_11770 n2_10458_11770 5.841270e-02
R10080 n2_10458_11770 n2_10505_11770 2.984127e-02
R10081 n2_10505_11770 n2_10554_11770 3.111111e-02
R10082 n2_10554_11770 n2_10646_11770 5.841270e-02
R10083 n2_10366_12799 n2_10458_12799 5.841270e-02
R10084 n2_10458_12799 n2_10505_12799 2.984127e-02
R10085 n2_10505_12799 n2_10554_12799 3.111111e-02
R10086 n2_10554_12799 n2_10646_12799 5.841270e-02
R10087 n2_10366_12895 n2_10458_12895 5.841270e-02
R10088 n2_10458_12895 n2_10505_12895 2.984127e-02
R10089 n2_10505_12895 n2_10554_12895 3.111111e-02
R10090 n2_10554_12895 n2_10646_12895 5.841270e-02
R10091 n2_10366_13924 n2_10458_13924 5.841270e-02
R10092 n2_10458_13924 n2_10505_13924 2.984127e-02
R10093 n2_10505_13924 n2_10554_13924 3.111111e-02
R10094 n2_10554_13924 n2_10646_13924 5.841270e-02
R10095 n2_10366_14020 n2_10458_14020 5.841270e-02
R10096 n2_10458_14020 n2_10505_14020 2.984127e-02
R10097 n2_10505_14020 n2_10554_14020 3.111111e-02
R10098 n2_10554_14020 n2_10646_14020 5.841270e-02
R10099 n2_10366_15049 n2_10458_15049 5.841270e-02
R10100 n2_10458_15049 n2_10505_15049 2.984127e-02
R10101 n2_10505_15049 n2_10554_15049 3.111111e-02
R10102 n2_10554_15049 n2_10646_15049 5.841270e-02
R10103 n2_10366_15145 n2_10458_15145 5.841270e-02
R10104 n2_10458_15145 n2_10505_15145 2.984127e-02
R10105 n2_10505_15145 n2_10554_15145 3.111111e-02
R10106 n2_10554_15145 n2_10646_15145 5.841270e-02
R10107 n2_10366_16174 n2_10458_16174 5.841270e-02
R10108 n2_10458_16174 n2_10505_16174 2.984127e-02
R10109 n2_10505_16174 n2_10554_16174 3.111111e-02
R10110 n2_10554_16174 n2_10646_16174 5.841270e-02
R10111 n2_10366_16270 n2_10458_16270 5.841270e-02
R10112 n2_10458_16270 n2_10505_16270 2.984127e-02
R10113 n2_10505_16270 n2_10554_16270 3.111111e-02
R10114 n2_10554_16270 n2_10646_16270 5.841270e-02
R10115 n2_10366_17299 n2_10458_17299 5.841270e-02
R10116 n2_10458_17299 n2_10505_17299 2.984127e-02
R10117 n2_10505_17299 n2_10554_17299 3.111111e-02
R10118 n2_10554_17299 n2_10646_17299 5.841270e-02
R10119 n2_10366_17395 n2_10458_17395 5.841270e-02
R10120 n2_10458_17395 n2_10505_17395 2.984127e-02
R10121 n2_10505_17395 n2_10554_17395 3.111111e-02
R10122 n2_10554_17395 n2_10646_17395 5.841270e-02
R10123 n2_10366_18424 n2_10458_18424 5.841270e-02
R10124 n2_10458_18424 n2_10505_18424 2.984127e-02
R10125 n2_10505_18424 n2_10554_18424 3.111111e-02
R10126 n2_10554_18424 n2_10646_18424 5.841270e-02
R10127 n2_10366_18520 n2_10458_18520 5.841270e-02
R10128 n2_10458_18520 n2_10505_18520 2.984127e-02
R10129 n2_10505_18520 n2_10554_18520 3.111111e-02
R10130 n2_10554_18520 n2_10646_18520 5.841270e-02
R10131 n2_10366_19549 n2_10458_19549 5.841270e-02
R10132 n2_10458_19549 n2_10505_19549 2.984127e-02
R10133 n2_10505_19549 n2_10554_19549 3.111111e-02
R10134 n2_10554_19549 n2_10646_19549 5.841270e-02
R10135 n2_10366_19645 n2_10458_19645 5.841270e-02
R10136 n2_10458_19645 n2_10505_19645 2.984127e-02
R10137 n2_10505_19645 n2_10554_19645 3.111111e-02
R10138 n2_10554_19645 n2_10646_19645 5.841270e-02
R10139 n2_10366_20674 n2_10458_20674 5.841270e-02
R10140 n2_10458_20674 n2_10505_20674 2.984127e-02
R10141 n2_10505_20674 n2_10554_20674 3.111111e-02
R10142 n2_10554_20674 n2_10646_20674 5.841270e-02
R10143 n2_10366_20770 n2_10458_20770 5.841270e-02
R10144 n2_10458_20770 n2_10505_20770 2.984127e-02
R10145 n2_10505_20770 n2_10554_20770 3.111111e-02
R10146 n2_10554_20770 n2_10646_20770 5.841270e-02
R10147 n2_10458_201 n2_10458_234 2.095238e-02
R10148 n2_10458_234 n2_10458_417 1.161905e-01
R10149 n2_10458_417 n2_10458_424 4.444444e-03
R10150 n2_10458_424 n2_10458_450 1.650794e-02
R10151 n2_10458_450 n2_10458_520 4.444444e-02
R10152 n2_10458_520 n2_10458_633 7.174603e-02
R10153 n2_10458_633 n2_10458_666 2.095238e-02
R10154 n2_10458_666 n2_10458_849 1.161905e-01
R10155 n2_10458_849 n2_10458_882 2.095238e-02
R10156 n2_10458_882 n2_10458_1065 1.161905e-01
R10157 n2_10458_1065 n2_10458_1098 2.095238e-02
R10158 n2_10458_1098 n2_10458_1281 1.161905e-01
R10159 n2_10458_1281 n2_10458_1314 2.095238e-02
R10160 n2_10458_1314 n2_10458_1497 1.161905e-01
R10161 n2_10458_1497 n2_10458_1530 2.095238e-02
R10162 n2_10458_1530 n2_10458_1549 1.206349e-02
R10163 n2_10458_1549 n2_10458_1645 6.095238e-02
R10164 n2_10458_1645 n2_10458_1713 4.317460e-02
R10165 n2_10458_1713 n2_10458_1746 2.095238e-02
R10166 n2_10458_1746 n2_10458_1760 8.888889e-03
R10167 n2_10458_1760 n2_10458_1783 1.460317e-02
R10168 n2_10458_1783 n2_10458_1929 9.269841e-02
R10169 n2_10458_1929 n2_10458_1962 2.095238e-02
R10170 n2_10458_1962 n2_10458_2145 1.161905e-01
R10171 n2_10458_2145 n2_10458_2178 2.095238e-02
R10172 n2_10458_2178 n2_10458_2361 1.161905e-01
R10173 n2_10458_2361 n2_10458_2394 2.095238e-02
R10174 n2_10458_2394 n2_10458_2408 8.888889e-03
R10175 n2_10458_2408 n2_10458_2577 1.073016e-01
R10176 n2_10458_2577 n2_10458_2610 2.095238e-02
R10177 n2_10458_2610 n2_10458_2647 2.349206e-02
R10178 n2_10458_2647 n2_10458_2674 1.714286e-02
R10179 n2_10458_2674 n2_10458_2770 6.095238e-02
R10180 n2_10458_2770 n2_10458_2793 1.460317e-02
R10181 n2_10458_2793 n2_10458_2826 2.095238e-02
R10182 n2_10458_2826 n2_10458_2840 8.888889e-03
R10183 n2_10458_2840 n2_10458_2863 1.460317e-02
R10184 n2_10458_2863 n2_10458_3009 9.269841e-02
R10185 n2_10458_3009 n2_10458_3042 2.095238e-02
R10186 n2_10458_3042 n2_10458_3225 1.161905e-01
R10187 n2_10458_3225 n2_10458_3258 2.095238e-02
R10188 n2_10458_3258 n2_10458_3441 1.161905e-01
R10189 n2_10458_3441 n2_10458_3474 2.095238e-02
R10190 n2_10458_3474 n2_10458_3488 8.888889e-03
R10191 n2_10458_3488 n2_10458_3511 1.460317e-02
R10192 n2_10458_3511 n2_10458_3657 9.269841e-02
R10193 n2_10458_3657 n2_10458_3690 2.095238e-02
R10194 n2_10458_3690 n2_10458_3799 6.920635e-02
R10195 n2_10458_3799 n2_10458_3873 4.698413e-02
R10196 n2_10458_3873 n2_10458_3895 1.396825e-02
R10197 n2_10458_3895 n2_10458_3906 6.984127e-03
R10198 n2_10458_3906 n2_10458_4089 1.161905e-01
R10199 n2_10458_4089 n2_10458_4122 2.095238e-02
R10200 n2_10458_4122 n2_10458_4136 8.888889e-03
R10201 n2_10458_4136 n2_10458_4159 1.460317e-02
R10202 n2_10458_4159 n2_10458_4305 9.269841e-02
R10203 n2_10458_4305 n2_10458_4338 2.095238e-02
R10204 n2_10458_4338 n2_10458_4521 1.161905e-01
R10205 n2_10458_4521 n2_10458_4554 2.095238e-02
R10206 n2_10458_4554 n2_10458_4568 8.888889e-03
R10207 n2_10458_4568 n2_10458_4591 1.460317e-02
R10208 n2_10458_4591 n2_10458_4737 9.269841e-02
R10209 n2_10458_4737 n2_10458_4770 2.095238e-02
R10210 n2_10458_4770 n2_10458_4924 9.777778e-02
R10211 n2_10458_4924 n2_10458_4953 1.841270e-02
R10212 n2_10458_4953 n2_10458_4986 2.095238e-02
R10213 n2_10458_4986 n2_10458_5020 2.158730e-02
R10214 n2_10458_5020 n2_10458_5169 9.460317e-02
R10215 n2_10458_5169 n2_10458_5202 2.095238e-02
R10216 n2_10458_5202 n2_10458_5239 2.349206e-02
R10217 n2_10458_5239 n2_10458_5385 9.269841e-02
R10218 n2_10458_5385 n2_10458_5418 2.095238e-02
R10219 n2_10458_5418 n2_10458_5432 8.888889e-03
R10220 n2_10458_5432 n2_10458_5455 1.460317e-02
R10221 n2_10458_5455 n2_10458_5601 9.269841e-02
R10222 n2_10458_5601 n2_10458_5634 2.095238e-02
R10223 n2_10458_5634 n2_10458_5817 1.161905e-01
R10224 n2_10458_5817 n2_10458_5850 2.095238e-02
R10225 n2_10458_5850 n2_10458_6033 1.161905e-01
R10226 n2_10458_6033 n2_10458_6049 1.015873e-02
R10227 n2_10458_6049 n2_10458_6066 1.079365e-02
R10228 n2_10458_6066 n2_10458_6145 5.015873e-02
R10229 n2_10458_6145 n2_10458_6249 6.603175e-02
R10230 n2_10458_6249 n2_10458_6282 2.095238e-02
R10231 n2_10458_6282 n2_10458_6465 1.161905e-01
R10232 n2_10458_6465 n2_10458_6498 2.095238e-02
R10233 n2_10458_6498 n2_10458_6512 8.888889e-03
R10234 n2_10458_6512 n2_10458_6535 1.460317e-02
R10235 n2_10458_6535 n2_10458_6681 9.269841e-02
R10236 n2_10458_6681 n2_10458_6714 2.095238e-02
R10237 n2_10458_6714 n2_10458_6751 2.349206e-02
R10238 n2_10458_6751 n2_10458_6897 9.269841e-02
R10239 n2_10458_6897 n2_10458_6930 2.095238e-02
R10240 n2_10458_6930 n2_10458_6944 8.888889e-03
R10241 n2_10458_6944 n2_10458_6967 1.460317e-02
R10242 n2_10458_6967 n2_10458_7113 9.269841e-02
R10243 n2_10458_7113 n2_10458_7146 2.095238e-02
R10244 n2_10458_7146 n2_10458_7160 8.888889e-03
R10245 n2_10458_7160 n2_10458_7174 8.888889e-03
R10246 n2_10458_7174 n2_10458_7178 2.539683e-03
R10247 n2_10458_7178 n2_10458_7270 5.841270e-02
R10248 n2_10458_7270 n2_10458_7329 3.746032e-02
R10249 n2_10458_7329 n2_10458_7362 2.095238e-02
R10250 n2_10458_7362 n2_10458_7376 8.888889e-03
R10251 n2_10458_7376 n2_10458_7399 1.460317e-02
R10252 n2_10458_7399 n2_10458_7545 9.269841e-02
R10253 n2_10458_7545 n2_10458_7578 2.095238e-02
R10254 n2_10458_7578 n2_10458_7761 1.161905e-01
R10255 n2_10458_7761 n2_10458_7794 2.095238e-02
R10256 n2_10458_7794 n2_10458_7977 1.161905e-01
R10257 n2_10458_7977 n2_10458_8010 2.095238e-02
R10258 n2_10458_8010 n2_10458_8193 1.161905e-01
R10259 n2_10458_8193 n2_10458_8226 2.095238e-02
R10260 n2_10458_8226 n2_10458_8299 4.634921e-02
R10261 n2_10458_8299 n2_10458_8395 6.095238e-02
R10262 n2_10458_8395 n2_10458_8409 8.888889e-03
R10263 n2_10458_8409 n2_10458_8442 2.095238e-02
R10264 n2_10458_8442 n2_10458_8625 1.161905e-01
R10265 n2_10458_8625 n2_10458_8658 2.095238e-02
R10266 n2_10458_8658 n2_10458_8841 1.161905e-01
R10267 n2_10458_8841 n2_10458_8874 2.095238e-02
R10268 n2_10458_8874 n2_10458_9057 1.161905e-01
R10269 n2_10458_9057 n2_10458_9090 2.095238e-02
R10270 n2_10458_9090 n2_10458_9273 1.161905e-01
R10271 n2_10458_9273 n2_10458_9306 2.095238e-02
R10272 n2_10458_9306 n2_10458_9424 7.492063e-02
R10273 n2_10458_9424 n2_10458_9489 4.126984e-02
R10274 n2_10458_9489 n2_10458_9520 1.968254e-02
R10275 n2_10458_9520 n2_10458_9522 1.269841e-03
R10276 n2_10458_9522 n2_10458_9705 1.161905e-01
R10277 n2_10458_9705 n2_10458_9738 2.095238e-02
R10278 n2_10458_9738 n2_10458_9921 1.161905e-01
R10279 n2_10458_9921 n2_10458_9954 2.095238e-02
R10280 n2_10458_9954 n2_10458_10137 1.161905e-01
R10281 n2_10458_10137 n2_10458_10170 2.095238e-02
R10282 n2_10458_10170 n2_10458_10353 1.161905e-01
R10283 n2_10458_10353 n2_10458_10386 2.095238e-02
R10284 n2_10458_10386 n2_10458_10549 1.034921e-01
R10285 n2_10458_10549 n2_10458_10569 1.269841e-02
R10286 n2_10458_10569 n2_10458_10602 2.095238e-02
R10287 n2_10458_10602 n2_10458_10645 2.730159e-02
R10288 n2_10458_10645 n2_10458_10785 8.888889e-02
R10289 n2_10458_10785 n2_10458_10818 2.095238e-02
R10290 n2_10458_10818 n2_10458_11001 1.161905e-01
R10291 n2_10458_11001 n2_10458_11034 2.095238e-02
R10292 n2_10458_11034 n2_10458_11217 1.161905e-01
R10293 n2_10458_11217 n2_10458_11250 2.095238e-02
R10294 n2_10458_11250 n2_10458_11433 1.161905e-01
R10295 n2_10458_11433 n2_10458_11466 2.095238e-02
R10296 n2_10458_11466 n2_10458_11649 1.161905e-01
R10297 n2_10458_11649 n2_10458_11674 1.587302e-02
R10298 n2_10458_11674 n2_10458_11682 5.079365e-03
R10299 n2_10458_11682 n2_10458_11770 5.587302e-02
R10300 n2_10458_11770 n2_10458_11865 6.031746e-02
R10301 n2_10458_11865 n2_10458_11898 2.095238e-02
R10302 n2_10458_11898 n2_10458_12081 1.161905e-01
R10303 n2_10458_12081 n2_10458_12114 2.095238e-02
R10304 n2_10458_12114 n2_10458_12297 1.161905e-01
R10305 n2_10458_12297 n2_10458_12330 2.095238e-02
R10306 n2_10458_12330 n2_10458_12513 1.161905e-01
R10307 n2_10458_12513 n2_10458_12546 2.095238e-02
R10308 n2_10458_12546 n2_10458_12729 1.161905e-01
R10309 n2_10458_12729 n2_10458_12762 2.095238e-02
R10310 n2_10458_12762 n2_10458_12799 2.349206e-02
R10311 n2_10458_12799 n2_10458_12895 6.095238e-02
R10312 n2_10458_12895 n2_10458_12945 3.174603e-02
R10313 n2_10458_12945 n2_10458_12978 2.095238e-02
R10314 n2_10458_12978 n2_10458_13161 1.161905e-01
R10315 n2_10458_13161 n2_10458_13194 2.095238e-02
R10316 n2_10458_13194 n2_10458_13377 1.161905e-01
R10317 n2_10458_13377 n2_10458_13410 2.095238e-02
R10318 n2_10458_13410 n2_10458_13593 1.161905e-01
R10319 n2_10458_13593 n2_10458_13626 2.095238e-02
R10320 n2_10458_13626 n2_10458_13640 8.888889e-03
R10321 n2_10458_13640 n2_10458_13663 1.460317e-02
R10322 n2_10458_13663 n2_10458_13809 9.269841e-02
R10323 n2_10458_13809 n2_10458_13842 2.095238e-02
R10324 n2_10458_13842 n2_10458_13856 8.888889e-03
R10325 n2_10458_13856 n2_10458_13879 1.460317e-02
R10326 n2_10458_13879 n2_10458_13924 2.857143e-02
R10327 n2_10458_13924 n2_10458_14020 6.095238e-02
R10328 n2_10458_14020 n2_10458_14025 3.174603e-03
R10329 n2_10458_14025 n2_10458_14058 2.095238e-02
R10330 n2_10458_14058 n2_10458_14072 8.888889e-03
R10331 n2_10458_14072 n2_10458_14079 4.444444e-03
R10332 n2_10458_14079 n2_10458_14241 1.028571e-01
R10333 n2_10458_14241 n2_10458_14274 2.095238e-02
R10334 n2_10458_14274 n2_10458_14457 1.161905e-01
R10335 n2_10458_14457 n2_10458_14490 2.095238e-02
R10336 n2_10458_14490 n2_10458_14504 8.888889e-03
R10337 n2_10458_14504 n2_10458_14673 1.073016e-01
R10338 n2_10458_14673 n2_10458_14706 2.095238e-02
R10339 n2_10458_14706 n2_10458_14889 1.161905e-01
R10340 n2_10458_14889 n2_10458_14922 2.095238e-02
R10341 n2_10458_14922 n2_10458_15049 8.063492e-02
R10342 n2_10458_15049 n2_10458_15105 3.555556e-02
R10343 n2_10458_15105 n2_10458_15138 2.095238e-02
R10344 n2_10458_15138 n2_10458_15145 4.444444e-03
R10345 n2_10458_15145 n2_10458_15321 1.117460e-01
R10346 n2_10458_15321 n2_10458_15354 2.095238e-02
R10347 n2_10458_15354 n2_10458_15537 1.161905e-01
R10348 n2_10458_15537 n2_10458_15570 2.095238e-02
R10349 n2_10458_15570 n2_10458_15584 8.888889e-03
R10350 n2_10458_15584 n2_10458_15753 1.073016e-01
R10351 n2_10458_15753 n2_10458_15786 2.095238e-02
R10352 n2_10458_15786 n2_10458_15800 8.888889e-03
R10353 n2_10458_15800 n2_10458_15823 1.460317e-02
R10354 n2_10458_15823 n2_10458_15969 9.269841e-02
R10355 n2_10458_15969 n2_10458_16002 2.095238e-02
R10356 n2_10458_16002 n2_10458_16016 8.888889e-03
R10357 n2_10458_16016 n2_10458_16174 1.003175e-01
R10358 n2_10458_16174 n2_10458_16185 6.984127e-03
R10359 n2_10458_16185 n2_10458_16218 2.095238e-02
R10360 n2_10458_16218 n2_10458_16270 3.301587e-02
R10361 n2_10458_16270 n2_10458_16401 8.317460e-02
R10362 n2_10458_16401 n2_10458_16434 2.095238e-02
R10363 n2_10458_16434 n2_10458_16617 1.161905e-01
R10364 n2_10458_16617 n2_10458_16650 2.095238e-02
R10365 n2_10458_16650 n2_10458_16833 1.161905e-01
R10366 n2_10458_16833 n2_10458_16866 2.095238e-02
R10367 n2_10458_16866 n2_10458_17049 1.161905e-01
R10368 n2_10458_17049 n2_10458_17082 2.095238e-02
R10369 n2_10458_17082 n2_10458_17096 8.888889e-03
R10370 n2_10458_17096 n2_10458_17103 4.444444e-03
R10371 n2_10458_17103 n2_10458_17119 1.015873e-02
R10372 n2_10458_17119 n2_10458_17265 9.269841e-02
R10373 n2_10458_17265 n2_10458_17298 2.095238e-02
R10374 n2_10458_17298 n2_10458_17299 6.349206e-04
R10375 n2_10458_17299 n2_10458_17312 8.253968e-03
R10376 n2_10458_17312 n2_10458_17395 5.269841e-02
R10377 n2_10458_17395 n2_10458_17481 5.460317e-02
R10378 n2_10458_17481 n2_10458_17514 2.095238e-02
R10379 n2_10458_17514 n2_10458_17697 1.161905e-01
R10380 n2_10458_17697 n2_10458_17730 2.095238e-02
R10381 n2_10458_17730 n2_10458_17913 1.161905e-01
R10382 n2_10458_17913 n2_10458_17946 2.095238e-02
R10383 n2_10458_17946 n2_10458_18129 1.161905e-01
R10384 n2_10458_18129 n2_10458_18162 2.095238e-02
R10385 n2_10458_18162 n2_10458_18345 1.161905e-01
R10386 n2_10458_18345 n2_10458_18378 2.095238e-02
R10387 n2_10458_18378 n2_10458_18392 8.888889e-03
R10388 n2_10458_18392 n2_10458_18424 2.031746e-02
R10389 n2_10458_18424 n2_10458_18520 6.095238e-02
R10390 n2_10458_18520 n2_10458_18561 2.603175e-02
R10391 n2_10458_18561 n2_10458_18594 2.095238e-02
R10392 n2_10458_18594 n2_10458_18608 8.888889e-03
R10393 n2_10458_18608 n2_10458_18777 1.073016e-01
R10394 n2_10458_18777 n2_10458_18810 2.095238e-02
R10395 n2_10458_18810 n2_10458_18993 1.161905e-01
R10396 n2_10458_18993 n2_10458_19026 2.095238e-02
R10397 n2_10458_19026 n2_10458_19209 1.161905e-01
R10398 n2_10458_19209 n2_10458_19242 2.095238e-02
R10399 n2_10458_19242 n2_10458_19256 8.888889e-03
R10400 n2_10458_19256 n2_10458_19425 1.073016e-01
R10401 n2_10458_19425 n2_10458_19458 2.095238e-02
R10402 n2_10458_19458 n2_10458_19549 5.777778e-02
R10403 n2_10458_19549 n2_10458_19641 5.841270e-02
R10404 n2_10458_19641 n2_10458_19645 2.539683e-03
R10405 n2_10458_19645 n2_10458_19674 1.841270e-02
R10406 n2_10458_19674 n2_10458_19857 1.161905e-01
R10407 n2_10458_19857 n2_10458_19890 2.095238e-02
R10408 n2_10458_19890 n2_10458_20073 1.161905e-01
R10409 n2_10458_20073 n2_10458_20106 2.095238e-02
R10410 n2_10458_20106 n2_10458_20289 1.161905e-01
R10411 n2_10458_20289 n2_10458_20322 2.095238e-02
R10412 n2_10458_20322 n2_10458_20505 1.161905e-01
R10413 n2_10458_20505 n2_10458_20538 2.095238e-02
R10414 n2_10458_20538 n2_10458_20674 8.634921e-02
R10415 n2_10458_20674 n2_10458_20721 2.984127e-02
R10416 n2_10458_20721 n2_10458_20754 2.095238e-02
R10417 n2_10458_20754 n2_10458_20770 1.015873e-02
R10418 n2_10458_20770 n2_10458_20937 1.060317e-01
R10419 n2_10458_20937 n2_10458_20970 2.095238e-02
R10420 n2_10554_201 n2_10554_234 2.095238e-02
R10421 n2_10554_234 n2_10554_417 1.161905e-01
R10422 n2_10554_417 n2_10554_424 4.444444e-03
R10423 n2_10554_424 n2_10554_450 1.650794e-02
R10424 n2_10554_450 n2_10554_520 4.444444e-02
R10425 n2_10554_520 n2_10554_633 7.174603e-02
R10426 n2_10554_633 n2_10554_666 2.095238e-02
R10427 n2_10554_666 n2_10554_849 1.161905e-01
R10428 n2_10554_849 n2_10554_882 2.095238e-02
R10429 n2_10554_882 n2_10554_1065 1.161905e-01
R10430 n2_10554_1065 n2_10554_1098 2.095238e-02
R10431 n2_10554_1098 n2_10554_1281 1.161905e-01
R10432 n2_10554_1281 n2_10554_1314 2.095238e-02
R10433 n2_10554_1314 n2_10554_1497 1.161905e-01
R10434 n2_10554_1497 n2_10554_1530 2.095238e-02
R10435 n2_10554_1530 n2_10554_1549 1.206349e-02
R10436 n2_10554_1549 n2_10554_1645 6.095238e-02
R10437 n2_10554_1645 n2_10554_1713 4.317460e-02
R10438 n2_10554_1713 n2_10554_1746 2.095238e-02
R10439 n2_10554_1746 n2_10554_1760 8.888889e-03
R10440 n2_10554_1760 n2_10554_1783 1.460317e-02
R10441 n2_10554_1783 n2_10554_1929 9.269841e-02
R10442 n2_10554_1929 n2_10554_1962 2.095238e-02
R10443 n2_10554_1962 n2_10554_2145 1.161905e-01
R10444 n2_10554_2145 n2_10554_2178 2.095238e-02
R10445 n2_10554_2178 n2_10554_2361 1.161905e-01
R10446 n2_10554_2361 n2_10554_2394 2.095238e-02
R10447 n2_10554_2394 n2_10554_2408 8.888889e-03
R10448 n2_10554_2408 n2_10554_2577 1.073016e-01
R10449 n2_10554_2577 n2_10554_2610 2.095238e-02
R10450 n2_10554_2610 n2_10554_2647 2.349206e-02
R10451 n2_10554_2647 n2_10554_2674 1.714286e-02
R10452 n2_10554_2674 n2_10554_2770 6.095238e-02
R10453 n2_10554_2770 n2_10554_2793 1.460317e-02
R10454 n2_10554_2793 n2_10554_2826 2.095238e-02
R10455 n2_10554_2826 n2_10554_2840 8.888889e-03
R10456 n2_10554_2840 n2_10554_2863 1.460317e-02
R10457 n2_10554_2863 n2_10554_3009 9.269841e-02
R10458 n2_10554_3009 n2_10554_3042 2.095238e-02
R10459 n2_10554_3042 n2_10554_3225 1.161905e-01
R10460 n2_10554_3225 n2_10554_3258 2.095238e-02
R10461 n2_10554_3258 n2_10554_3441 1.161905e-01
R10462 n2_10554_3441 n2_10554_3474 2.095238e-02
R10463 n2_10554_3474 n2_10554_3488 8.888889e-03
R10464 n2_10554_3488 n2_10554_3511 1.460317e-02
R10465 n2_10554_3511 n2_10554_3657 9.269841e-02
R10466 n2_10554_3657 n2_10554_3690 2.095238e-02
R10467 n2_10554_3690 n2_10554_3799 6.920635e-02
R10468 n2_10554_3799 n2_10554_3873 4.698413e-02
R10469 n2_10554_3873 n2_10554_3895 1.396825e-02
R10470 n2_10554_3895 n2_10554_3906 6.984127e-03
R10471 n2_10554_3906 n2_10554_4089 1.161905e-01
R10472 n2_10554_4089 n2_10554_4122 2.095238e-02
R10473 n2_10554_4122 n2_10554_4136 8.888889e-03
R10474 n2_10554_4136 n2_10554_4159 1.460317e-02
R10475 n2_10554_4159 n2_10554_4305 9.269841e-02
R10476 n2_10554_4305 n2_10554_4338 2.095238e-02
R10477 n2_10554_4338 n2_10554_4521 1.161905e-01
R10478 n2_10554_4521 n2_10554_4554 2.095238e-02
R10479 n2_10554_4554 n2_10554_4568 8.888889e-03
R10480 n2_10554_4568 n2_10554_4591 1.460317e-02
R10481 n2_10554_4591 n2_10554_4737 9.269841e-02
R10482 n2_10554_4737 n2_10554_4770 2.095238e-02
R10483 n2_10554_4770 n2_10554_4924 9.777778e-02
R10484 n2_10554_4924 n2_10554_4953 1.841270e-02
R10485 n2_10554_4953 n2_10554_4986 2.095238e-02
R10486 n2_10554_4986 n2_10554_5020 2.158730e-02
R10487 n2_10554_5020 n2_10554_5169 9.460317e-02
R10488 n2_10554_5169 n2_10554_5202 2.095238e-02
R10489 n2_10554_5202 n2_10554_5239 2.349206e-02
R10490 n2_10554_5239 n2_10554_5385 9.269841e-02
R10491 n2_10554_5385 n2_10554_5418 2.095238e-02
R10492 n2_10554_5418 n2_10554_5432 8.888889e-03
R10493 n2_10554_5432 n2_10554_5455 1.460317e-02
R10494 n2_10554_5455 n2_10554_5601 9.269841e-02
R10495 n2_10554_5601 n2_10554_5634 2.095238e-02
R10496 n2_10554_5634 n2_10554_5817 1.161905e-01
R10497 n2_10554_5817 n2_10554_5850 2.095238e-02
R10498 n2_10554_5850 n2_10554_6033 1.161905e-01
R10499 n2_10554_6033 n2_10554_6049 1.015873e-02
R10500 n2_10554_6049 n2_10554_6066 1.079365e-02
R10501 n2_10554_6066 n2_10554_6145 5.015873e-02
R10502 n2_10554_6145 n2_10554_6249 6.603175e-02
R10503 n2_10554_6249 n2_10554_6282 2.095238e-02
R10504 n2_10554_6282 n2_10554_6465 1.161905e-01
R10505 n2_10554_6465 n2_10554_6498 2.095238e-02
R10506 n2_10554_6498 n2_10554_6512 8.888889e-03
R10507 n2_10554_6512 n2_10554_6535 1.460317e-02
R10508 n2_10554_6535 n2_10554_6681 9.269841e-02
R10509 n2_10554_6681 n2_10554_6714 2.095238e-02
R10510 n2_10554_6714 n2_10554_6751 2.349206e-02
R10511 n2_10554_6751 n2_10554_6897 9.269841e-02
R10512 n2_10554_6897 n2_10554_6930 2.095238e-02
R10513 n2_10554_6930 n2_10554_6944 8.888889e-03
R10514 n2_10554_6944 n2_10554_6967 1.460317e-02
R10515 n2_10554_6967 n2_10554_7113 9.269841e-02
R10516 n2_10554_7113 n2_10554_7146 2.095238e-02
R10517 n2_10554_7146 n2_10554_7160 8.888889e-03
R10518 n2_10554_7160 n2_10554_7174 8.888889e-03
R10519 n2_10554_7174 n2_10554_7178 2.539683e-03
R10520 n2_10554_7178 n2_10554_7270 5.841270e-02
R10521 n2_10554_7270 n2_10554_7329 3.746032e-02
R10522 n2_10554_7329 n2_10554_7362 2.095238e-02
R10523 n2_10554_7362 n2_10554_7376 8.888889e-03
R10524 n2_10554_7376 n2_10554_7399 1.460317e-02
R10525 n2_10554_7399 n2_10554_7545 9.269841e-02
R10526 n2_10554_7545 n2_10554_7578 2.095238e-02
R10527 n2_10554_7578 n2_10554_7761 1.161905e-01
R10528 n2_10554_7761 n2_10554_7794 2.095238e-02
R10529 n2_10554_7794 n2_10554_7977 1.161905e-01
R10530 n2_10554_7977 n2_10554_8010 2.095238e-02
R10531 n2_10554_8010 n2_10554_8193 1.161905e-01
R10532 n2_10554_8193 n2_10554_8226 2.095238e-02
R10533 n2_10554_8226 n2_10554_8299 4.634921e-02
R10534 n2_10554_8299 n2_10554_8395 6.095238e-02
R10535 n2_10554_8395 n2_10554_8409 8.888889e-03
R10536 n2_10554_8409 n2_10554_8442 2.095238e-02
R10537 n2_10554_8442 n2_10554_8625 1.161905e-01
R10538 n2_10554_8625 n2_10554_8658 2.095238e-02
R10539 n2_10554_8658 n2_10554_8841 1.161905e-01
R10540 n2_10554_8841 n2_10554_8874 2.095238e-02
R10541 n2_10554_8874 n2_10554_9057 1.161905e-01
R10542 n2_10554_9057 n2_10554_9090 2.095238e-02
R10543 n2_10554_9090 n2_10554_9273 1.161905e-01
R10544 n2_10554_9273 n2_10554_9306 2.095238e-02
R10545 n2_10554_9306 n2_10554_9424 7.492063e-02
R10546 n2_10554_9424 n2_10554_9489 4.126984e-02
R10547 n2_10554_9489 n2_10554_9520 1.968254e-02
R10548 n2_10554_9520 n2_10554_9522 1.269841e-03
R10549 n2_10554_9522 n2_10554_9705 1.161905e-01
R10550 n2_10554_9705 n2_10554_9738 2.095238e-02
R10551 n2_10554_9738 n2_10554_9921 1.161905e-01
R10552 n2_10554_9921 n2_10554_9954 2.095238e-02
R10553 n2_10554_9954 n2_10554_10137 1.161905e-01
R10554 n2_10554_10137 n2_10554_10170 2.095238e-02
R10555 n2_10554_10170 n2_10554_10353 1.161905e-01
R10556 n2_10554_10353 n2_10554_10386 2.095238e-02
R10557 n2_10554_10386 n2_10554_10549 1.034921e-01
R10558 n2_10554_10549 n2_10554_10569 1.269841e-02
R10559 n2_10554_10569 n2_10554_10602 2.095238e-02
R10560 n2_10554_10602 n2_10554_10645 2.730159e-02
R10561 n2_10554_10645 n2_10554_10785 8.888889e-02
R10562 n2_10554_10785 n2_10554_10818 2.095238e-02
R10563 n2_10554_10818 n2_10554_11001 1.161905e-01
R10564 n2_10554_11001 n2_10554_11034 2.095238e-02
R10565 n2_10554_11034 n2_10554_11217 1.161905e-01
R10566 n2_10554_11217 n2_10554_11250 2.095238e-02
R10567 n2_10554_11250 n2_10554_11433 1.161905e-01
R10568 n2_10554_11433 n2_10554_11466 2.095238e-02
R10569 n2_10554_11466 n2_10554_11649 1.161905e-01
R10570 n2_10554_11649 n2_10554_11674 1.587302e-02
R10571 n2_10554_11674 n2_10554_11682 5.079365e-03
R10572 n2_10554_11682 n2_10554_11770 5.587302e-02
R10573 n2_10554_11770 n2_10554_11865 6.031746e-02
R10574 n2_10554_11865 n2_10554_11898 2.095238e-02
R10575 n2_10554_11898 n2_10554_12081 1.161905e-01
R10576 n2_10554_12081 n2_10554_12114 2.095238e-02
R10577 n2_10554_12114 n2_10554_12297 1.161905e-01
R10578 n2_10554_12297 n2_10554_12330 2.095238e-02
R10579 n2_10554_12330 n2_10554_12513 1.161905e-01
R10580 n2_10554_12513 n2_10554_12546 2.095238e-02
R10581 n2_10554_12546 n2_10554_12729 1.161905e-01
R10582 n2_10554_12729 n2_10554_12762 2.095238e-02
R10583 n2_10554_12762 n2_10554_12799 2.349206e-02
R10584 n2_10554_12799 n2_10554_12895 6.095238e-02
R10585 n2_10554_12895 n2_10554_12945 3.174603e-02
R10586 n2_10554_12945 n2_10554_12978 2.095238e-02
R10587 n2_10554_12978 n2_10554_13161 1.161905e-01
R10588 n2_10554_13161 n2_10554_13194 2.095238e-02
R10589 n2_10554_13194 n2_10554_13377 1.161905e-01
R10590 n2_10554_13377 n2_10554_13410 2.095238e-02
R10591 n2_10554_13410 n2_10554_13593 1.161905e-01
R10592 n2_10554_13593 n2_10554_13626 2.095238e-02
R10593 n2_10554_13626 n2_10554_13640 8.888889e-03
R10594 n2_10554_13640 n2_10554_13663 1.460317e-02
R10595 n2_10554_13663 n2_10554_13809 9.269841e-02
R10596 n2_10554_13809 n2_10554_13842 2.095238e-02
R10597 n2_10554_13842 n2_10554_13856 8.888889e-03
R10598 n2_10554_13856 n2_10554_13879 1.460317e-02
R10599 n2_10554_13879 n2_10554_13924 2.857143e-02
R10600 n2_10554_13924 n2_10554_14020 6.095238e-02
R10601 n2_10554_14020 n2_10554_14025 3.174603e-03
R10602 n2_10554_14025 n2_10554_14058 2.095238e-02
R10603 n2_10554_14058 n2_10554_14072 8.888889e-03
R10604 n2_10554_14072 n2_10554_14079 4.444444e-03
R10605 n2_10554_14079 n2_10554_14241 1.028571e-01
R10606 n2_10554_14241 n2_10554_14274 2.095238e-02
R10607 n2_10554_14274 n2_10554_14457 1.161905e-01
R10608 n2_10554_14457 n2_10554_14490 2.095238e-02
R10609 n2_10554_14490 n2_10554_14504 8.888889e-03
R10610 n2_10554_14504 n2_10554_14673 1.073016e-01
R10611 n2_10554_14673 n2_10554_14706 2.095238e-02
R10612 n2_10554_14706 n2_10554_14889 1.161905e-01
R10613 n2_10554_14889 n2_10554_14922 2.095238e-02
R10614 n2_10554_14922 n2_10554_15049 8.063492e-02
R10615 n2_10554_15049 n2_10554_15105 3.555556e-02
R10616 n2_10554_15105 n2_10554_15138 2.095238e-02
R10617 n2_10554_15138 n2_10554_15145 4.444444e-03
R10618 n2_10554_15145 n2_10554_15321 1.117460e-01
R10619 n2_10554_15321 n2_10554_15354 2.095238e-02
R10620 n2_10554_15354 n2_10554_15537 1.161905e-01
R10621 n2_10554_15537 n2_10554_15570 2.095238e-02
R10622 n2_10554_15570 n2_10554_15584 8.888889e-03
R10623 n2_10554_15584 n2_10554_15753 1.073016e-01
R10624 n2_10554_15753 n2_10554_15786 2.095238e-02
R10625 n2_10554_15786 n2_10554_15800 8.888889e-03
R10626 n2_10554_15800 n2_10554_15823 1.460317e-02
R10627 n2_10554_15823 n2_10554_15969 9.269841e-02
R10628 n2_10554_15969 n2_10554_16002 2.095238e-02
R10629 n2_10554_16002 n2_10554_16016 8.888889e-03
R10630 n2_10554_16016 n2_10554_16174 1.003175e-01
R10631 n2_10554_16174 n2_10554_16185 6.984127e-03
R10632 n2_10554_16185 n2_10554_16218 2.095238e-02
R10633 n2_10554_16218 n2_10554_16270 3.301587e-02
R10634 n2_10554_16270 n2_10554_16401 8.317460e-02
R10635 n2_10554_16401 n2_10554_16434 2.095238e-02
R10636 n2_10554_16434 n2_10554_16617 1.161905e-01
R10637 n2_10554_16617 n2_10554_16650 2.095238e-02
R10638 n2_10554_16650 n2_10554_16833 1.161905e-01
R10639 n2_10554_16833 n2_10554_16866 2.095238e-02
R10640 n2_10554_16866 n2_10554_17049 1.161905e-01
R10641 n2_10554_17049 n2_10554_17082 2.095238e-02
R10642 n2_10554_17082 n2_10554_17096 8.888889e-03
R10643 n2_10554_17096 n2_10554_17103 4.444444e-03
R10644 n2_10554_17103 n2_10554_17119 1.015873e-02
R10645 n2_10554_17119 n2_10554_17265 9.269841e-02
R10646 n2_10554_17265 n2_10554_17298 2.095238e-02
R10647 n2_10554_17298 n2_10554_17299 6.349206e-04
R10648 n2_10554_17299 n2_10554_17312 8.253968e-03
R10649 n2_10554_17312 n2_10554_17395 5.269841e-02
R10650 n2_10554_17395 n2_10554_17481 5.460317e-02
R10651 n2_10554_17481 n2_10554_17514 2.095238e-02
R10652 n2_10554_17514 n2_10554_17697 1.161905e-01
R10653 n2_10554_17697 n2_10554_17730 2.095238e-02
R10654 n2_10554_17730 n2_10554_17913 1.161905e-01
R10655 n2_10554_17913 n2_10554_17946 2.095238e-02
R10656 n2_10554_17946 n2_10554_18129 1.161905e-01
R10657 n2_10554_18129 n2_10554_18162 2.095238e-02
R10658 n2_10554_18162 n2_10554_18345 1.161905e-01
R10659 n2_10554_18345 n2_10554_18378 2.095238e-02
R10660 n2_10554_18378 n2_10554_18392 8.888889e-03
R10661 n2_10554_18392 n2_10554_18424 2.031746e-02
R10662 n2_10554_18424 n2_10554_18520 6.095238e-02
R10663 n2_10554_18520 n2_10554_18561 2.603175e-02
R10664 n2_10554_18561 n2_10554_18594 2.095238e-02
R10665 n2_10554_18594 n2_10554_18608 8.888889e-03
R10666 n2_10554_18608 n2_10554_18777 1.073016e-01
R10667 n2_10554_18777 n2_10554_18810 2.095238e-02
R10668 n2_10554_18810 n2_10554_18993 1.161905e-01
R10669 n2_10554_18993 n2_10554_19026 2.095238e-02
R10670 n2_10554_19026 n2_10554_19209 1.161905e-01
R10671 n2_10554_19209 n2_10554_19242 2.095238e-02
R10672 n2_10554_19242 n2_10554_19256 8.888889e-03
R10673 n2_10554_19256 n2_10554_19425 1.073016e-01
R10674 n2_10554_19425 n2_10554_19458 2.095238e-02
R10675 n2_10554_19458 n2_10554_19549 5.777778e-02
R10676 n2_10554_19549 n2_10554_19641 5.841270e-02
R10677 n2_10554_19641 n2_10554_19645 2.539683e-03
R10678 n2_10554_19645 n2_10554_19674 1.841270e-02
R10679 n2_10554_19674 n2_10554_19857 1.161905e-01
R10680 n2_10554_19857 n2_10554_19890 2.095238e-02
R10681 n2_10554_19890 n2_10554_20073 1.161905e-01
R10682 n2_10554_20073 n2_10554_20106 2.095238e-02
R10683 n2_10554_20106 n2_10554_20289 1.161905e-01
R10684 n2_10554_20289 n2_10554_20322 2.095238e-02
R10685 n2_10554_20322 n2_10554_20505 1.161905e-01
R10686 n2_10554_20505 n2_10554_20538 2.095238e-02
R10687 n2_10554_20538 n2_10554_20674 8.634921e-02
R10688 n2_10554_20674 n2_10554_20721 2.984127e-02
R10689 n2_10554_20721 n2_10554_20754 2.095238e-02
R10690 n2_10554_20754 n2_10554_20770 1.015873e-02
R10691 n2_10554_20770 n2_10554_20937 1.060317e-01
R10692 n2_10554_20937 n2_10554_20970 2.095238e-02
R10693 n2_10646_201 n2_10646_234 2.095238e-02
R10694 n2_10646_234 n2_10646_417 1.161905e-01
R10695 n2_10646_417 n2_10646_424 4.444444e-03
R10696 n2_10646_424 n2_10646_450 1.650794e-02
R10697 n2_10646_520 n2_10646_633 7.174603e-02
R10698 n2_10646_633 n2_10646_666 2.095238e-02
R10699 n2_10646_666 n2_10646_849 1.161905e-01
R10700 n2_10646_849 n2_10646_882 2.095238e-02
R10701 n2_10646_882 n2_10646_1065 1.161905e-01
R10702 n2_10646_1065 n2_10646_1098 2.095238e-02
R10703 n2_10646_1098 n2_10646_1281 1.161905e-01
R10704 n2_10646_1281 n2_10646_1314 2.095238e-02
R10705 n2_10646_1314 n2_10646_1497 1.161905e-01
R10706 n2_10646_1497 n2_10646_1530 2.095238e-02
R10707 n2_10646_1530 n2_10646_1549 1.206349e-02
R10708 n2_10646_1645 n2_10646_1713 4.317460e-02
R10709 n2_10646_1713 n2_10646_1746 2.095238e-02
R10710 n2_10646_1746 n2_10646_1760 8.888889e-03
R10711 n2_10646_1760 n2_10646_1783 1.460317e-02
R10712 n2_10646_1783 n2_10646_1929 9.269841e-02
R10713 n2_10646_1929 n2_10646_1962 2.095238e-02
R10714 n2_10646_1962 n2_10646_2145 1.161905e-01
R10715 n2_10646_2145 n2_10646_2178 2.095238e-02
R10716 n2_10646_2178 n2_10646_2361 1.161905e-01
R10717 n2_10646_2361 n2_10646_2394 2.095238e-02
R10718 n2_10646_2394 n2_10646_2408 8.888889e-03
R10719 n2_10646_2408 n2_10646_2577 1.073016e-01
R10720 n2_10646_2577 n2_10646_2610 2.095238e-02
R10721 n2_10646_2610 n2_10646_2647 2.349206e-02
R10722 n2_10646_2647 n2_10646_2674 1.714286e-02
R10723 n2_10646_2770 n2_10646_2793 1.460317e-02
R10724 n2_10646_2793 n2_10646_2826 2.095238e-02
R10725 n2_10646_2826 n2_10646_2840 8.888889e-03
R10726 n2_10646_2840 n2_10646_2863 1.460317e-02
R10727 n2_10646_2863 n2_10646_3009 9.269841e-02
R10728 n2_10646_3009 n2_10646_3042 2.095238e-02
R10729 n2_10646_3042 n2_10646_3225 1.161905e-01
R10730 n2_10646_3225 n2_10646_3258 2.095238e-02
R10731 n2_10646_3258 n2_10646_3441 1.161905e-01
R10732 n2_10646_3441 n2_10646_3474 2.095238e-02
R10733 n2_10646_3474 n2_10646_3488 8.888889e-03
R10734 n2_10646_3488 n2_10646_3511 1.460317e-02
R10735 n2_10646_3511 n2_10646_3657 9.269841e-02
R10736 n2_10646_3657 n2_10646_3690 2.095238e-02
R10737 n2_10646_3690 n2_10646_3799 6.920635e-02
R10738 n2_10646_3873 n2_10646_3895 1.396825e-02
R10739 n2_10646_3895 n2_10646_3906 6.984127e-03
R10740 n2_10646_3906 n2_10646_4089 1.161905e-01
R10741 n2_10646_4089 n2_10646_4122 2.095238e-02
R10742 n2_10646_4122 n2_10646_4136 8.888889e-03
R10743 n2_10646_4136 n2_10646_4159 1.460317e-02
R10744 n2_10646_4159 n2_10646_4305 9.269841e-02
R10745 n2_10646_4305 n2_10646_4338 2.095238e-02
R10746 n2_10646_4338 n2_10646_4521 1.161905e-01
R10747 n2_10646_4521 n2_10646_4554 2.095238e-02
R10748 n2_10646_4554 n2_10646_4568 8.888889e-03
R10749 n2_10646_4568 n2_10646_4591 1.460317e-02
R10750 n2_10646_4591 n2_10646_4737 9.269841e-02
R10751 n2_10646_4737 n2_10646_4770 2.095238e-02
R10752 n2_10646_4770 n2_10646_4924 9.777778e-02
R10753 n2_10646_4924 n2_10646_4953 1.841270e-02
R10754 n2_10646_5020 n2_10646_5169 9.460317e-02
R10755 n2_10646_5169 n2_10646_5202 2.095238e-02
R10756 n2_10646_5202 n2_10646_5239 2.349206e-02
R10757 n2_10646_5239 n2_10646_5385 9.269841e-02
R10758 n2_10646_5385 n2_10646_5418 2.095238e-02
R10759 n2_10646_5418 n2_10646_5432 8.888889e-03
R10760 n2_10646_5432 n2_10646_5455 1.460317e-02
R10761 n2_10646_5455 n2_10646_5601 9.269841e-02
R10762 n2_10646_5601 n2_10646_5634 2.095238e-02
R10763 n2_10646_5634 n2_10646_5817 1.161905e-01
R10764 n2_10646_5817 n2_10646_5850 2.095238e-02
R10765 n2_10646_5850 n2_10646_6033 1.161905e-01
R10766 n2_10646_6033 n2_10646_6049 1.015873e-02
R10767 n2_10646_6049 n2_10646_6066 1.079365e-02
R10768 n2_10646_6145 n2_10646_6249 6.603175e-02
R10769 n2_10646_6249 n2_10646_6282 2.095238e-02
R10770 n2_10646_6282 n2_10646_6465 1.161905e-01
R10771 n2_10646_6465 n2_10646_6498 2.095238e-02
R10772 n2_10646_6498 n2_10646_6512 8.888889e-03
R10773 n2_10646_6512 n2_10646_6535 1.460317e-02
R10774 n2_10646_6535 n2_10646_6681 9.269841e-02
R10775 n2_10646_6681 n2_10646_6714 2.095238e-02
R10776 n2_10646_6714 n2_10646_6751 2.349206e-02
R10777 n2_10646_6751 n2_10646_6897 9.269841e-02
R10778 n2_10646_6897 n2_10646_6930 2.095238e-02
R10779 n2_10646_6930 n2_10646_6944 8.888889e-03
R10780 n2_10646_6944 n2_10646_6967 1.460317e-02
R10781 n2_10646_6967 n2_10646_7113 9.269841e-02
R10782 n2_10646_7113 n2_10646_7146 2.095238e-02
R10783 n2_10646_7146 n2_10646_7160 8.888889e-03
R10784 n2_10646_7160 n2_10646_7174 8.888889e-03
R10785 n2_10646_7174 n2_10646_7178 2.539683e-03
R10786 n2_10646_7270 n2_10646_7329 3.746032e-02
R10787 n2_10646_7329 n2_10646_7362 2.095238e-02
R10788 n2_10646_7362 n2_10646_7376 8.888889e-03
R10789 n2_10646_7376 n2_10646_7399 1.460317e-02
R10790 n2_10646_7399 n2_10646_7545 9.269841e-02
R10791 n2_10646_7545 n2_10646_7578 2.095238e-02
R10792 n2_10646_7578 n2_10646_7761 1.161905e-01
R10793 n2_10646_7761 n2_10646_7794 2.095238e-02
R10794 n2_10646_7794 n2_10646_7977 1.161905e-01
R10795 n2_10646_7977 n2_10646_8010 2.095238e-02
R10796 n2_10646_8010 n2_10646_8193 1.161905e-01
R10797 n2_10646_8193 n2_10646_8226 2.095238e-02
R10798 n2_10646_8226 n2_10646_8299 4.634921e-02
R10799 n2_10646_8395 n2_10646_8409 8.888889e-03
R10800 n2_10646_8409 n2_10646_8442 2.095238e-02
R10801 n2_10646_8442 n2_10646_8613 1.085714e-01
R10802 n2_10646_8613 n2_10646_8625 7.619048e-03
R10803 n2_10646_8625 n2_10646_8658 2.095238e-02
R10804 n2_10646_8658 n2_10646_8841 1.161905e-01
R10805 n2_10646_8841 n2_10646_8874 2.095238e-02
R10806 n2_10646_8874 n2_10646_9057 1.161905e-01
R10807 n2_10646_9057 n2_10646_9090 2.095238e-02
R10808 n2_10646_9090 n2_10646_9190 6.349206e-02
R10809 n2_10646_9190 n2_10646_9273 5.269841e-02
R10810 n2_10646_9273 n2_10646_9306 2.095238e-02
R10811 n2_10646_9306 n2_10646_9424 7.492063e-02
R10812 n2_10646_9489 n2_10646_9520 1.968254e-02
R10813 n2_10646_9520 n2_10646_9522 1.269841e-03
R10814 n2_10646_9522 n2_10646_9705 1.161905e-01
R10815 n2_10646_9705 n2_10646_9738 2.095238e-02
R10816 n2_10646_9738 n2_10646_9921 1.161905e-01
R10817 n2_10646_9921 n2_10646_9954 2.095238e-02
R10818 n2_10646_9954 n2_10646_10137 1.161905e-01
R10819 n2_10646_10137 n2_10646_10170 2.095238e-02
R10820 n2_10646_10170 n2_10646_10353 1.161905e-01
R10821 n2_10646_10353 n2_10646_10386 2.095238e-02
R10822 n2_10646_10386 n2_10646_10549 1.034921e-01
R10823 n2_10646_10549 n2_10646_10569 1.269841e-02
R10824 n2_10646_10645 n2_10646_10785 8.888889e-02
R10825 n2_10646_10785 n2_10646_10818 2.095238e-02
R10826 n2_10646_10818 n2_10646_11001 1.161905e-01
R10827 n2_10646_11001 n2_10646_11034 2.095238e-02
R10828 n2_10646_11034 n2_10646_11217 1.161905e-01
R10829 n2_10646_11217 n2_10646_11250 2.095238e-02
R10830 n2_10646_11250 n2_10646_11433 1.161905e-01
R10831 n2_10646_11433 n2_10646_11466 2.095238e-02
R10832 n2_10646_11466 n2_10646_11649 1.161905e-01
R10833 n2_10646_11649 n2_10646_11674 1.587302e-02
R10834 n2_10646_11674 n2_10646_11682 5.079365e-03
R10835 n2_10646_11770 n2_10646_11865 6.031746e-02
R10836 n2_10646_11865 n2_10646_11898 2.095238e-02
R10837 n2_10646_11898 n2_10646_12004 6.730159e-02
R10838 n2_10646_12004 n2_10646_12081 4.888889e-02
R10839 n2_10646_12081 n2_10646_12114 2.095238e-02
R10840 n2_10646_12114 n2_10646_12297 1.161905e-01
R10841 n2_10646_12297 n2_10646_12330 2.095238e-02
R10842 n2_10646_12330 n2_10646_12513 1.161905e-01
R10843 n2_10646_12513 n2_10646_12546 2.095238e-02
R10844 n2_10646_12546 n2_10646_12566 1.269841e-02
R10845 n2_10646_12566 n2_10646_12729 1.034921e-01
R10846 n2_10646_12729 n2_10646_12762 2.095238e-02
R10847 n2_10646_12762 n2_10646_12799 2.349206e-02
R10848 n2_10646_12895 n2_10646_12945 3.174603e-02
R10849 n2_10646_12945 n2_10646_12978 2.095238e-02
R10850 n2_10646_12978 n2_10646_13161 1.161905e-01
R10851 n2_10646_13161 n2_10646_13194 2.095238e-02
R10852 n2_10646_13194 n2_10646_13377 1.161905e-01
R10853 n2_10646_13377 n2_10646_13410 2.095238e-02
R10854 n2_10646_13410 n2_10646_13593 1.161905e-01
R10855 n2_10646_13593 n2_10646_13626 2.095238e-02
R10856 n2_10646_13626 n2_10646_13640 8.888889e-03
R10857 n2_10646_13640 n2_10646_13663 1.460317e-02
R10858 n2_10646_13663 n2_10646_13809 9.269841e-02
R10859 n2_10646_13809 n2_10646_13842 2.095238e-02
R10860 n2_10646_13842 n2_10646_13856 8.888889e-03
R10861 n2_10646_13856 n2_10646_13879 1.460317e-02
R10862 n2_10646_13879 n2_10646_13924 2.857143e-02
R10863 n2_10646_14020 n2_10646_14025 3.174603e-03
R10864 n2_10646_14025 n2_10646_14058 2.095238e-02
R10865 n2_10646_14058 n2_10646_14072 8.888889e-03
R10866 n2_10646_14072 n2_10646_14079 4.444444e-03
R10867 n2_10646_14079 n2_10646_14241 1.028571e-01
R10868 n2_10646_14241 n2_10646_14274 2.095238e-02
R10869 n2_10646_14274 n2_10646_14457 1.161905e-01
R10870 n2_10646_14457 n2_10646_14490 2.095238e-02
R10871 n2_10646_14490 n2_10646_14504 8.888889e-03
R10872 n2_10646_14504 n2_10646_14673 1.073016e-01
R10873 n2_10646_14673 n2_10646_14706 2.095238e-02
R10874 n2_10646_14706 n2_10646_14889 1.161905e-01
R10875 n2_10646_14889 n2_10646_14922 2.095238e-02
R10876 n2_10646_14922 n2_10646_15049 8.063492e-02
R10877 n2_10646_15138 n2_10646_15145 4.444444e-03
R10878 n2_10646_15145 n2_10646_15321 1.117460e-01
R10879 n2_10646_15321 n2_10646_15354 2.095238e-02
R10880 n2_10646_15354 n2_10646_15537 1.161905e-01
R10881 n2_10646_15537 n2_10646_15570 2.095238e-02
R10882 n2_10646_15570 n2_10646_15584 8.888889e-03
R10883 n2_10646_15584 n2_10646_15753 1.073016e-01
R10884 n2_10646_15753 n2_10646_15786 2.095238e-02
R10885 n2_10646_15786 n2_10646_15800 8.888889e-03
R10886 n2_10646_15800 n2_10646_15823 1.460317e-02
R10887 n2_10646_15823 n2_10646_15969 9.269841e-02
R10888 n2_10646_15969 n2_10646_16002 2.095238e-02
R10889 n2_10646_16002 n2_10646_16016 8.888889e-03
R10890 n2_10646_16016 n2_10646_16174 1.003175e-01
R10891 n2_10646_16174 n2_10646_16185 6.984127e-03
R10892 n2_10646_16270 n2_10646_16401 8.317460e-02
R10893 n2_10646_16401 n2_10646_16434 2.095238e-02
R10894 n2_10646_16434 n2_10646_16617 1.161905e-01
R10895 n2_10646_16617 n2_10646_16650 2.095238e-02
R10896 n2_10646_16650 n2_10646_16833 1.161905e-01
R10897 n2_10646_16833 n2_10646_16866 2.095238e-02
R10898 n2_10646_16866 n2_10646_17049 1.161905e-01
R10899 n2_10646_17049 n2_10646_17082 2.095238e-02
R10900 n2_10646_17082 n2_10646_17096 8.888889e-03
R10901 n2_10646_17096 n2_10646_17103 4.444444e-03
R10902 n2_10646_17103 n2_10646_17119 1.015873e-02
R10903 n2_10646_17119 n2_10646_17265 9.269841e-02
R10904 n2_10646_17265 n2_10646_17298 2.095238e-02
R10905 n2_10646_17298 n2_10646_17299 6.349206e-04
R10906 n2_10646_17299 n2_10646_17312 8.253968e-03
R10907 n2_10646_17395 n2_10646_17481 5.460317e-02
R10908 n2_10646_17481 n2_10646_17514 2.095238e-02
R10909 n2_10646_17514 n2_10646_17697 1.161905e-01
R10910 n2_10646_17697 n2_10646_17730 2.095238e-02
R10911 n2_10646_17730 n2_10646_17913 1.161905e-01
R10912 n2_10646_17913 n2_10646_17946 2.095238e-02
R10913 n2_10646_17946 n2_10646_18129 1.161905e-01
R10914 n2_10646_18129 n2_10646_18162 2.095238e-02
R10915 n2_10646_18162 n2_10646_18345 1.161905e-01
R10916 n2_10646_18345 n2_10646_18378 2.095238e-02
R10917 n2_10646_18378 n2_10646_18392 8.888889e-03
R10918 n2_10646_18392 n2_10646_18424 2.031746e-02
R10919 n2_10646_18520 n2_10646_18561 2.603175e-02
R10920 n2_10646_18561 n2_10646_18594 2.095238e-02
R10921 n2_10646_18594 n2_10646_18608 8.888889e-03
R10922 n2_10646_18608 n2_10646_18777 1.073016e-01
R10923 n2_10646_18777 n2_10646_18810 2.095238e-02
R10924 n2_10646_18810 n2_10646_18993 1.161905e-01
R10925 n2_10646_18993 n2_10646_19026 2.095238e-02
R10926 n2_10646_19026 n2_10646_19209 1.161905e-01
R10927 n2_10646_19209 n2_10646_19242 2.095238e-02
R10928 n2_10646_19242 n2_10646_19256 8.888889e-03
R10929 n2_10646_19256 n2_10646_19425 1.073016e-01
R10930 n2_10646_19425 n2_10646_19458 2.095238e-02
R10931 n2_10646_19458 n2_10646_19549 5.777778e-02
R10932 n2_10646_19641 n2_10646_19645 2.539683e-03
R10933 n2_10646_19645 n2_10646_19674 1.841270e-02
R10934 n2_10646_19674 n2_10646_19857 1.161905e-01
R10935 n2_10646_19857 n2_10646_19890 2.095238e-02
R10936 n2_10646_19890 n2_10646_20073 1.161905e-01
R10937 n2_10646_20073 n2_10646_20106 2.095238e-02
R10938 n2_10646_20106 n2_10646_20289 1.161905e-01
R10939 n2_10646_20289 n2_10646_20322 2.095238e-02
R10940 n2_10646_20322 n2_10646_20505 1.161905e-01
R10941 n2_10646_20505 n2_10646_20538 2.095238e-02
R10942 n2_10646_20538 n2_10646_20674 8.634921e-02
R10943 n2_10646_20754 n2_10646_20770 1.015873e-02
R10944 n2_10646_20770 n2_10646_20937 1.060317e-01
R10945 n2_10646_20937 n2_10646_20970 2.095238e-02
R10946 n2_11491_9489 n2_11491_9522 2.095238e-02
R10947 n2_11491_9522 n2_11491_9705 1.161905e-01
R10948 n2_11491_9705 n2_11491_9738 2.095238e-02
R10949 n2_11491_9738 n2_11491_9921 1.161905e-01
R10950 n2_11491_9921 n2_11491_9954 2.095238e-02
R10951 n2_11491_9954 n2_11491_10137 1.161905e-01
R10952 n2_11491_10137 n2_11491_10170 2.095238e-02
R10953 n2_11491_10170 n2_11491_10353 1.161905e-01
R10954 n2_11491_10353 n2_11491_10386 2.095238e-02
R10955 n2_11491_10386 n2_11491_10549 1.034921e-01
R10956 n2_11491_10549 n2_11491_10569 1.269841e-02
R10957 n2_11491_10645 n2_11491_10785 8.888889e-02
R10958 n2_11491_10785 n2_11491_10818 2.095238e-02
R10959 n2_11491_10818 n2_11491_11001 1.161905e-01
R10960 n2_11491_11001 n2_11491_11034 2.095238e-02
R10961 n2_11491_11034 n2_11491_11217 1.161905e-01
R10962 n2_11491_11217 n2_11491_11250 2.095238e-02
R10963 n2_11491_11250 n2_11491_11433 1.161905e-01
R10964 n2_11491_11433 n2_11491_11466 2.095238e-02
R10965 n2_11491_11466 n2_11491_11649 1.161905e-01
R10966 n2_11491_11649 n2_11491_11682 2.095238e-02
R10967 n2_11491_10549 n2_11630_10549 8.825397e-02
R10968 n2_11630_10549 n2_11679_10549 3.111111e-02
R10969 n2_11491_10645 n2_11630_10645 8.825397e-02
R10970 n2_11630_10645 n2_11679_10645 3.111111e-02
R10971 n2_11679_9705 n2_11679_9738 2.095238e-02
R10972 n2_11679_9738 n2_11679_9921 1.161905e-01
R10973 n2_11679_9921 n2_11679_9954 2.095238e-02
R10974 n2_11679_9954 n2_11679_10034 5.079365e-02
R10975 n2_11679_10034 n2_11679_10137 6.539683e-02
R10976 n2_11679_10137 n2_11679_10170 2.095238e-02
R10977 n2_11679_10170 n2_11679_10353 1.161905e-01
R10978 n2_11679_10353 n2_11679_10386 2.095238e-02
R10979 n2_11679_10386 n2_11679_10549 1.034921e-01
R10980 n2_11679_10549 n2_11679_10569 1.269841e-02
R10981 n2_11679_10569 n2_11679_10602 2.095238e-02
R10982 n2_11679_10602 n2_11679_10645 2.730159e-02
R10983 n2_11679_10645 n2_11679_10785 8.888889e-02
R10984 n2_11679_10785 n2_11679_10818 2.095238e-02
R10985 n2_11679_10818 n2_11679_11001 1.161905e-01
R10986 n2_11679_11001 n2_11679_11034 2.095238e-02
R10987 n2_11679_11034 n2_11679_11160 8.000000e-02
R10988 n2_11679_11160 n2_11679_11217 3.619048e-02
R10989 n2_11679_11217 n2_11679_11250 2.095238e-02
R10990 n2_11679_11250 n2_11679_11433 1.161905e-01
R10991 n2_11679_11433 n2_11679_11466 2.095238e-02
R10992 n2_12616_201 n2_12616_234 2.095238e-02
R10993 n2_12616_234 n2_12616_417 1.161905e-01
R10994 n2_12616_417 n2_12616_424 4.444444e-03
R10995 n2_12616_424 n2_12616_450 1.650794e-02
R10996 n2_12616_520 n2_12616_633 7.174603e-02
R10997 n2_12616_633 n2_12616_666 2.095238e-02
R10998 n2_12616_666 n2_12616_849 1.161905e-01
R10999 n2_12616_849 n2_12616_882 2.095238e-02
R11000 n2_12616_882 n2_12616_1065 1.161905e-01
R11001 n2_12616_1065 n2_12616_1098 2.095238e-02
R11002 n2_12616_1098 n2_12616_1281 1.161905e-01
R11003 n2_12616_1281 n2_12616_1314 2.095238e-02
R11004 n2_12616_1314 n2_12616_1497 1.161905e-01
R11005 n2_12616_1497 n2_12616_1530 2.095238e-02
R11006 n2_12616_1530 n2_12616_1549 1.206349e-02
R11007 n2_12616_1645 n2_12616_1713 4.317460e-02
R11008 n2_12616_1713 n2_12616_1746 2.095238e-02
R11009 n2_12616_1746 n2_12616_1783 2.349206e-02
R11010 n2_12616_1783 n2_12616_1929 9.269841e-02
R11011 n2_12616_1929 n2_12616_1962 2.095238e-02
R11012 n2_12616_1962 n2_12616_2145 1.161905e-01
R11013 n2_12616_2145 n2_12616_2178 2.095238e-02
R11014 n2_12616_2178 n2_12616_2361 1.161905e-01
R11015 n2_12616_2361 n2_12616_2394 2.095238e-02
R11016 n2_12616_2394 n2_12616_2431 2.349206e-02
R11017 n2_12616_2431 n2_12616_2577 9.269841e-02
R11018 n2_12616_2577 n2_12616_2610 2.095238e-02
R11019 n2_12616_2610 n2_12616_2674 4.063492e-02
R11020 n2_12616_2770 n2_12616_2793 1.460317e-02
R11021 n2_12616_2793 n2_12616_2826 2.095238e-02
R11022 n2_12616_2826 n2_12616_2863 2.349206e-02
R11023 n2_12616_2863 n2_12616_3009 9.269841e-02
R11024 n2_12616_3009 n2_12616_3042 2.095238e-02
R11025 n2_12616_3042 n2_12616_3225 1.161905e-01
R11026 n2_12616_3225 n2_12616_3258 2.095238e-02
R11027 n2_12616_3258 n2_12616_3441 1.161905e-01
R11028 n2_12616_3441 n2_12616_3474 2.095238e-02
R11029 n2_12616_3474 n2_12616_3511 2.349206e-02
R11030 n2_12616_3511 n2_12616_3657 9.269841e-02
R11031 n2_12616_3657 n2_12616_3690 2.095238e-02
R11032 n2_12616_3690 n2_12616_3799 6.920635e-02
R11033 n2_12616_3873 n2_12616_3895 1.396825e-02
R11034 n2_12616_3895 n2_12616_3906 6.984127e-03
R11035 n2_12616_3906 n2_12616_3943 2.349206e-02
R11036 n2_12616_3943 n2_12616_4089 9.269841e-02
R11037 n2_12616_4089 n2_12616_4122 2.095238e-02
R11038 n2_12616_4122 n2_12616_4159 2.349206e-02
R11039 n2_12616_4159 n2_12616_4305 9.269841e-02
R11040 n2_12616_4305 n2_12616_4338 2.095238e-02
R11041 n2_12616_4338 n2_12616_4521 1.161905e-01
R11042 n2_12616_4521 n2_12616_4554 2.095238e-02
R11043 n2_12616_4554 n2_12616_4591 2.349206e-02
R11044 n2_12616_4591 n2_12616_4737 9.269841e-02
R11045 n2_12616_4737 n2_12616_4770 2.095238e-02
R11046 n2_12616_4770 n2_12616_4924 9.777778e-02
R11047 n2_12616_4924 n2_12616_4953 1.841270e-02
R11048 n2_12616_5020 n2_12616_5023 1.904762e-03
R11049 n2_12616_5023 n2_12616_5169 9.269841e-02
R11050 n2_12616_5169 n2_12616_5202 2.095238e-02
R11051 n2_12616_5202 n2_12616_5239 2.349206e-02
R11052 n2_12616_5239 n2_12616_5385 9.269841e-02
R11053 n2_12616_5385 n2_12616_5418 2.095238e-02
R11054 n2_12616_5418 n2_12616_5601 1.161905e-01
R11055 n2_12616_5601 n2_12616_5634 2.095238e-02
R11056 n2_12616_5634 n2_12616_5671 2.349206e-02
R11057 n2_12616_5671 n2_12616_5817 9.269841e-02
R11058 n2_12616_5817 n2_12616_5850 2.095238e-02
R11059 n2_12616_5850 n2_12616_6033 1.161905e-01
R11060 n2_12616_6033 n2_12616_6049 1.015873e-02
R11061 n2_12616_6049 n2_12616_6066 1.079365e-02
R11062 n2_12616_6145 n2_12616_6249 6.603175e-02
R11063 n2_12616_6249 n2_12616_6282 2.095238e-02
R11064 n2_12616_6282 n2_12616_6319 2.349206e-02
R11065 n2_12616_6319 n2_12616_6465 9.269841e-02
R11066 n2_12616_6465 n2_12616_6498 2.095238e-02
R11067 n2_12616_6498 n2_12616_6681 1.161905e-01
R11068 n2_12616_6681 n2_12616_6714 2.095238e-02
R11069 n2_12616_6714 n2_12616_6751 2.349206e-02
R11070 n2_12616_6751 n2_12616_6897 9.269841e-02
R11071 n2_12616_6897 n2_12616_6930 2.095238e-02
R11072 n2_12616_6930 n2_12616_6967 2.349206e-02
R11073 n2_12616_6967 n2_12616_7113 9.269841e-02
R11074 n2_12616_7113 n2_12616_7146 2.095238e-02
R11075 n2_12616_7146 n2_12616_7174 1.777778e-02
R11076 n2_12616_7174 n2_12616_7178 2.539683e-03
R11077 n2_12616_7270 n2_12616_7329 3.746032e-02
R11078 n2_12616_7329 n2_12616_7362 2.095238e-02
R11079 n2_12616_7362 n2_12616_7399 2.349206e-02
R11080 n2_12616_7399 n2_12616_7545 9.269841e-02
R11081 n2_12616_7545 n2_12616_7578 2.095238e-02
R11082 n2_12616_7578 n2_12616_7761 1.161905e-01
R11083 n2_12616_7761 n2_12616_7794 2.095238e-02
R11084 n2_12616_7794 n2_12616_7831 2.349206e-02
R11085 n2_12616_7831 n2_12616_7977 9.269841e-02
R11086 n2_12616_7977 n2_12616_8010 2.095238e-02
R11087 n2_12616_8010 n2_12616_8193 1.161905e-01
R11088 n2_12616_8193 n2_12616_8226 2.095238e-02
R11089 n2_12616_8226 n2_12616_8299 4.634921e-02
R11090 n2_12616_8395 n2_12616_8409 8.888889e-03
R11091 n2_12616_8409 n2_12616_8442 2.095238e-02
R11092 n2_12616_8442 n2_12616_8625 1.161905e-01
R11093 n2_12616_8625 n2_12616_8658 2.095238e-02
R11094 n2_12616_8658 n2_12616_8695 2.349206e-02
R11095 n2_12616_8695 n2_12616_8841 9.269841e-02
R11096 n2_12616_8841 n2_12616_8874 2.095238e-02
R11097 n2_12616_8874 n2_12616_8911 2.349206e-02
R11098 n2_12616_8911 n2_12616_8948 2.349206e-02
R11099 n2_12616_8948 n2_12616_9057 6.920635e-02
R11100 n2_12616_9057 n2_12616_9090 2.095238e-02
R11101 n2_12616_9090 n2_12616_9273 1.161905e-01
R11102 n2_12616_9273 n2_12616_9306 2.095238e-02
R11103 n2_12616_9306 n2_12616_9489 1.161905e-01
R11104 n2_12616_9489 n2_12616_9522 2.095238e-02
R11105 n2_12616_9522 n2_12616_9705 1.161905e-01
R11106 n2_12616_9705 n2_12616_9738 2.095238e-02
R11107 n2_12616_9738 n2_12616_9775 2.349206e-02
R11108 n2_12616_9775 n2_12616_9921 9.269841e-02
R11109 n2_12616_9921 n2_12616_9954 2.095238e-02
R11110 n2_12616_9954 n2_12616_9991 2.349206e-02
R11111 n2_12616_9991 n2_12616_10034 2.730159e-02
R11112 n2_12616_10034 n2_12616_10137 6.539683e-02
R11113 n2_12616_10137 n2_12616_10170 2.095238e-02
R11114 n2_12616_10170 n2_12616_10353 1.161905e-01
R11115 n2_12616_10353 n2_12616_10386 2.095238e-02
R11116 n2_12616_10386 n2_12616_10549 1.034921e-01
R11117 n2_12616_10549 n2_12616_10569 1.269841e-02
R11118 n2_12616_10645 n2_12616_10785 8.888889e-02
R11119 n2_12616_10785 n2_12616_10818 2.095238e-02
R11120 n2_12616_10818 n2_12616_10832 8.888889e-03
R11121 n2_12616_10832 n2_12616_11001 1.073016e-01
R11122 n2_12616_11001 n2_12616_11034 2.095238e-02
R11123 n2_12616_11034 n2_12616_11048 8.888889e-03
R11124 n2_12616_11048 n2_12616_11160 7.111111e-02
R11125 n2_12616_11160 n2_12616_11217 3.619048e-02
R11126 n2_12616_11217 n2_12616_11250 2.095238e-02
R11127 n2_12616_11250 n2_12616_11433 1.161905e-01
R11128 n2_12616_11433 n2_12616_11466 2.095238e-02
R11129 n2_12616_11466 n2_12616_11649 1.161905e-01
R11130 n2_12616_11649 n2_12616_11682 2.095238e-02
R11131 n2_12616_11682 n2_12616_11865 1.161905e-01
R11132 n2_12616_11865 n2_12616_11898 2.095238e-02
R11133 n2_12616_11898 n2_12616_11912 8.888889e-03
R11134 n2_12616_11912 n2_12616_12081 1.073016e-01
R11135 n2_12616_12081 n2_12616_12114 2.095238e-02
R11136 n2_12616_12114 n2_12616_12128 8.888889e-03
R11137 n2_12616_12128 n2_12616_12285 9.968254e-02
R11138 n2_12616_12285 n2_12616_12297 7.619048e-03
R11139 n2_12616_12297 n2_12616_12330 2.095238e-02
R11140 n2_12616_12330 n2_12616_12513 1.161905e-01
R11141 n2_12616_12513 n2_12616_12546 2.095238e-02
R11142 n2_12616_12546 n2_12616_12729 1.161905e-01
R11143 n2_12616_12729 n2_12616_12762 2.095238e-02
R11144 n2_12616_12762 n2_12616_12799 2.349206e-02
R11145 n2_12616_12895 n2_12616_12945 3.174603e-02
R11146 n2_12616_12945 n2_12616_12978 2.095238e-02
R11147 n2_12616_12978 n2_12616_13129 9.587302e-02
R11148 n2_12616_13129 n2_12616_13161 2.031746e-02
R11149 n2_12616_13161 n2_12616_13194 2.095238e-02
R11150 n2_12616_13194 n2_12616_13377 1.161905e-01
R11151 n2_12616_13377 n2_12616_13410 2.095238e-02
R11152 n2_12616_13410 n2_12616_13593 1.161905e-01
R11153 n2_12616_13593 n2_12616_13626 2.095238e-02
R11154 n2_12616_13626 n2_12616_13663 2.349206e-02
R11155 n2_12616_13663 n2_12616_13700 2.349206e-02
R11156 n2_12616_13700 n2_12616_13809 6.920635e-02
R11157 n2_12616_13809 n2_12616_13842 2.095238e-02
R11158 n2_12616_13842 n2_12616_13924 5.206349e-02
R11159 n2_12616_14020 n2_12616_14025 3.174603e-03
R11160 n2_12616_14025 n2_12616_14058 2.095238e-02
R11161 n2_12616_14058 n2_12616_14079 1.333333e-02
R11162 n2_12616_14079 n2_12616_14229 9.523810e-02
R11163 n2_12616_14229 n2_12616_14241 7.619048e-03
R11164 n2_12616_14241 n2_12616_14274 2.095238e-02
R11165 n2_12616_14274 n2_12616_14457 1.161905e-01
R11166 n2_12616_14457 n2_12616_14490 2.095238e-02
R11167 n2_12616_14490 n2_12616_14673 1.161905e-01
R11168 n2_12616_14673 n2_12616_14706 2.095238e-02
R11169 n2_12616_14706 n2_12616_14727 1.333333e-02
R11170 n2_12616_14727 n2_12616_14816 5.650794e-02
R11171 n2_12616_14816 n2_12616_14889 4.634921e-02
R11172 n2_12616_14889 n2_12616_14922 2.095238e-02
R11173 n2_12616_14922 n2_12616_15049 8.063492e-02
R11174 n2_12616_15138 n2_12616_15145 4.444444e-03
R11175 n2_12616_15145 n2_12616_15321 1.117460e-01
R11176 n2_12616_15321 n2_12616_15354 2.095238e-02
R11177 n2_12616_15354 n2_12616_15368 8.888889e-03
R11178 n2_12616_15368 n2_12616_15537 1.073016e-01
R11179 n2_12616_15537 n2_12616_15570 2.095238e-02
R11180 n2_12616_15570 n2_12616_15753 1.161905e-01
R11181 n2_12616_15753 n2_12616_15786 2.095238e-02
R11182 n2_12616_15786 n2_12616_15800 8.888889e-03
R11183 n2_12616_15800 n2_12616_15807 4.444444e-03
R11184 n2_12616_15807 n2_12616_15969 1.028571e-01
R11185 n2_12616_15969 n2_12616_16002 2.095238e-02
R11186 n2_12616_16002 n2_12616_16174 1.092063e-01
R11187 n2_12616_16174 n2_12616_16185 6.984127e-03
R11188 n2_12616_16270 n2_12616_16401 8.317460e-02
R11189 n2_12616_16401 n2_12616_16434 2.095238e-02
R11190 n2_12616_16434 n2_12616_16448 8.888889e-03
R11191 n2_12616_16448 n2_12616_16617 1.073016e-01
R11192 n2_12616_16617 n2_12616_16650 2.095238e-02
R11193 n2_12616_16650 n2_12616_16833 1.161905e-01
R11194 n2_12616_16833 n2_12616_16866 2.095238e-02
R11195 n2_12616_16866 n2_12616_17049 1.161905e-01
R11196 n2_12616_17049 n2_12616_17082 2.095238e-02
R11197 n2_12616_17082 n2_12616_17096 8.888889e-03
R11198 n2_12616_17096 n2_12616_17103 4.444444e-03
R11199 n2_12616_17103 n2_12616_17265 1.028571e-01
R11200 n2_12616_17265 n2_12616_17298 2.095238e-02
R11201 n2_12616_17298 n2_12616_17299 6.349206e-04
R11202 n2_12616_17395 n2_12616_17481 5.460317e-02
R11203 n2_12616_17481 n2_12616_17514 2.095238e-02
R11204 n2_12616_17514 n2_12616_17528 8.888889e-03
R11205 n2_12616_17528 n2_12616_17697 1.073016e-01
R11206 n2_12616_17697 n2_12616_17730 2.095238e-02
R11207 n2_12616_17730 n2_12616_17913 1.161905e-01
R11208 n2_12616_17913 n2_12616_17946 2.095238e-02
R11209 n2_12616_17946 n2_12616_17983 2.349206e-02
R11210 n2_12616_17983 n2_12616_18129 9.269841e-02
R11211 n2_12616_18129 n2_12616_18162 2.095238e-02
R11212 n2_12616_18162 n2_12616_18176 8.888889e-03
R11213 n2_12616_18176 n2_12616_18183 4.444444e-03
R11214 n2_12616_18183 n2_12616_18345 1.028571e-01
R11215 n2_12616_18345 n2_12616_18378 2.095238e-02
R11216 n2_12616_18378 n2_12616_18424 2.920635e-02
R11217 n2_12616_18520 n2_12616_18561 2.603175e-02
R11218 n2_12616_18561 n2_12616_18594 2.095238e-02
R11219 n2_12616_18594 n2_12616_18608 8.888889e-03
R11220 n2_12616_18608 n2_12616_18777 1.073016e-01
R11221 n2_12616_18777 n2_12616_18810 2.095238e-02
R11222 n2_12616_18810 n2_12616_18993 1.161905e-01
R11223 n2_12616_18993 n2_12616_19026 2.095238e-02
R11224 n2_12616_19026 n2_12616_19209 1.161905e-01
R11225 n2_12616_19209 n2_12616_19242 2.095238e-02
R11226 n2_12616_19242 n2_12616_19256 8.888889e-03
R11227 n2_12616_19256 n2_12616_19263 4.444444e-03
R11228 n2_12616_19263 n2_12616_19425 1.028571e-01
R11229 n2_12616_19425 n2_12616_19458 2.095238e-02
R11230 n2_12616_19458 n2_12616_19549 5.777778e-02
R11231 n2_12616_19641 n2_12616_19645 2.539683e-03
R11232 n2_12616_19645 n2_12616_19674 1.841270e-02
R11233 n2_12616_19674 n2_12616_19857 1.161905e-01
R11234 n2_12616_19857 n2_12616_19890 2.095238e-02
R11235 n2_12616_19890 n2_12616_20073 1.161905e-01
R11236 n2_12616_20073 n2_12616_20106 2.095238e-02
R11237 n2_12616_20106 n2_12616_20289 1.161905e-01
R11238 n2_12616_20289 n2_12616_20322 2.095238e-02
R11239 n2_12616_20322 n2_12616_20505 1.161905e-01
R11240 n2_12616_20505 n2_12616_20538 2.095238e-02
R11241 n2_12616_20538 n2_12616_20674 8.634921e-02
R11242 n2_12616_20754 n2_12616_20770 1.015873e-02
R11243 n2_12616_20770 n2_12616_20937 1.060317e-01
R11244 n2_12616_20937 n2_12616_20970 2.095238e-02
R11245 n2_12616_8395 n2_12708_8395 5.841270e-02
R11246 n2_12708_8395 n2_12755_8395 2.984127e-02
R11247 n2_12755_8395 n2_12804_8395 3.111111e-02
R11248 n2_12616_10549 n2_12755_10549 8.825397e-02
R11249 n2_12755_10549 n2_12804_10549 3.111111e-02
R11250 n2_12616_10645 n2_12755_10645 8.825397e-02
R11251 n2_12755_10645 n2_12804_10645 3.111111e-02
R11252 n2_12616_12799 n2_12708_12799 5.841270e-02
R11253 n2_12708_12799 n2_12755_12799 2.984127e-02
R11254 n2_12755_12799 n2_12804_12799 3.111111e-02
R11255 n2_12616_424 n2_12708_424 5.841270e-02
R11256 n2_12708_424 n2_12755_424 2.984127e-02
R11257 n2_12755_424 n2_12804_424 3.111111e-02
R11258 n2_12804_424 n2_12896_424 5.841270e-02
R11259 n2_12616_520 n2_12708_520 5.841270e-02
R11260 n2_12708_520 n2_12755_520 2.984127e-02
R11261 n2_12755_520 n2_12804_520 3.111111e-02
R11262 n2_12804_520 n2_12896_520 5.841270e-02
R11263 n2_12616_1549 n2_12708_1549 5.841270e-02
R11264 n2_12708_1549 n2_12755_1549 2.984127e-02
R11265 n2_12755_1549 n2_12804_1549 3.111111e-02
R11266 n2_12804_1549 n2_12896_1549 5.841270e-02
R11267 n2_12616_1645 n2_12708_1645 5.841270e-02
R11268 n2_12708_1645 n2_12755_1645 2.984127e-02
R11269 n2_12755_1645 n2_12804_1645 3.111111e-02
R11270 n2_12804_1645 n2_12896_1645 5.841270e-02
R11271 n2_12616_2674 n2_12708_2674 5.841270e-02
R11272 n2_12708_2674 n2_12755_2674 2.984127e-02
R11273 n2_12755_2674 n2_12804_2674 3.111111e-02
R11274 n2_12804_2674 n2_12896_2674 5.841270e-02
R11275 n2_12616_2770 n2_12708_2770 5.841270e-02
R11276 n2_12708_2770 n2_12755_2770 2.984127e-02
R11277 n2_12755_2770 n2_12804_2770 3.111111e-02
R11278 n2_12804_2770 n2_12896_2770 5.841270e-02
R11279 n2_12616_3799 n2_12708_3799 5.841270e-02
R11280 n2_12708_3799 n2_12755_3799 2.984127e-02
R11281 n2_12755_3799 n2_12804_3799 3.111111e-02
R11282 n2_12804_3799 n2_12896_3799 5.841270e-02
R11283 n2_12616_3895 n2_12708_3895 5.841270e-02
R11284 n2_12708_3895 n2_12755_3895 2.984127e-02
R11285 n2_12755_3895 n2_12804_3895 3.111111e-02
R11286 n2_12804_3895 n2_12896_3895 5.841270e-02
R11287 n2_12616_4924 n2_12708_4924 5.841270e-02
R11288 n2_12708_4924 n2_12755_4924 2.984127e-02
R11289 n2_12755_4924 n2_12804_4924 3.111111e-02
R11290 n2_12804_4924 n2_12896_4924 5.841270e-02
R11291 n2_12616_5020 n2_12708_5020 5.841270e-02
R11292 n2_12708_5020 n2_12755_5020 2.984127e-02
R11293 n2_12755_5020 n2_12804_5020 3.111111e-02
R11294 n2_12804_5020 n2_12896_5020 5.841270e-02
R11295 n2_12616_6049 n2_12708_6049 5.841270e-02
R11296 n2_12708_6049 n2_12755_6049 2.984127e-02
R11297 n2_12755_6049 n2_12804_6049 3.111111e-02
R11298 n2_12804_6049 n2_12896_6049 5.841270e-02
R11299 n2_12616_6145 n2_12708_6145 5.841270e-02
R11300 n2_12708_6145 n2_12755_6145 2.984127e-02
R11301 n2_12755_6145 n2_12804_6145 3.111111e-02
R11302 n2_12804_6145 n2_12896_6145 5.841270e-02
R11303 n2_12616_7174 n2_12708_7174 5.841270e-02
R11304 n2_12708_7174 n2_12755_7174 2.984127e-02
R11305 n2_12755_7174 n2_12804_7174 3.111111e-02
R11306 n2_12804_7174 n2_12896_7174 5.841270e-02
R11307 n2_12616_7270 n2_12708_7270 5.841270e-02
R11308 n2_12708_7270 n2_12755_7270 2.984127e-02
R11309 n2_12755_7270 n2_12804_7270 3.111111e-02
R11310 n2_12804_7270 n2_12896_7270 5.841270e-02
R11311 n2_12616_8299 n2_12708_8299 5.841270e-02
R11312 n2_12708_8299 n2_12755_8299 2.984127e-02
R11313 n2_12755_8299 n2_12804_8299 3.111111e-02
R11314 n2_12804_8299 n2_12896_8299 5.841270e-02
R11315 n2_12616_12895 n2_12708_12895 5.841270e-02
R11316 n2_12708_12895 n2_12755_12895 2.984127e-02
R11317 n2_12755_12895 n2_12804_12895 3.111111e-02
R11318 n2_12804_12895 n2_12896_12895 5.841270e-02
R11319 n2_12616_13924 n2_12708_13924 5.841270e-02
R11320 n2_12708_13924 n2_12755_13924 2.984127e-02
R11321 n2_12755_13924 n2_12804_13924 3.111111e-02
R11322 n2_12804_13924 n2_12896_13924 5.841270e-02
R11323 n2_12616_14020 n2_12708_14020 5.841270e-02
R11324 n2_12708_14020 n2_12755_14020 2.984127e-02
R11325 n2_12755_14020 n2_12804_14020 3.111111e-02
R11326 n2_12804_14020 n2_12896_14020 5.841270e-02
R11327 n2_12616_15049 n2_12708_15049 5.841270e-02
R11328 n2_12708_15049 n2_12755_15049 2.984127e-02
R11329 n2_12755_15049 n2_12804_15049 3.111111e-02
R11330 n2_12804_15049 n2_12896_15049 5.841270e-02
R11331 n2_12616_15145 n2_12708_15145 5.841270e-02
R11332 n2_12708_15145 n2_12755_15145 2.984127e-02
R11333 n2_12755_15145 n2_12804_15145 3.111111e-02
R11334 n2_12804_15145 n2_12896_15145 5.841270e-02
R11335 n2_12616_16174 n2_12708_16174 5.841270e-02
R11336 n2_12708_16174 n2_12755_16174 2.984127e-02
R11337 n2_12755_16174 n2_12804_16174 3.111111e-02
R11338 n2_12804_16174 n2_12896_16174 5.841270e-02
R11339 n2_12616_16270 n2_12708_16270 5.841270e-02
R11340 n2_12708_16270 n2_12755_16270 2.984127e-02
R11341 n2_12755_16270 n2_12804_16270 3.111111e-02
R11342 n2_12804_16270 n2_12896_16270 5.841270e-02
R11343 n2_12616_17299 n2_12708_17299 5.841270e-02
R11344 n2_12708_17299 n2_12755_17299 2.984127e-02
R11345 n2_12755_17299 n2_12804_17299 3.111111e-02
R11346 n2_12804_17299 n2_12896_17299 5.841270e-02
R11347 n2_12616_17395 n2_12708_17395 5.841270e-02
R11348 n2_12708_17395 n2_12755_17395 2.984127e-02
R11349 n2_12755_17395 n2_12804_17395 3.111111e-02
R11350 n2_12804_17395 n2_12896_17395 5.841270e-02
R11351 n2_12616_18424 n2_12708_18424 5.841270e-02
R11352 n2_12708_18424 n2_12755_18424 2.984127e-02
R11353 n2_12755_18424 n2_12804_18424 3.111111e-02
R11354 n2_12804_18424 n2_12896_18424 5.841270e-02
R11355 n2_12616_18520 n2_12708_18520 5.841270e-02
R11356 n2_12708_18520 n2_12755_18520 2.984127e-02
R11357 n2_12755_18520 n2_12804_18520 3.111111e-02
R11358 n2_12804_18520 n2_12896_18520 5.841270e-02
R11359 n2_12616_19549 n2_12708_19549 5.841270e-02
R11360 n2_12708_19549 n2_12755_19549 2.984127e-02
R11361 n2_12755_19549 n2_12804_19549 3.111111e-02
R11362 n2_12804_19549 n2_12896_19549 5.841270e-02
R11363 n2_12616_19645 n2_12708_19645 5.841270e-02
R11364 n2_12708_19645 n2_12755_19645 2.984127e-02
R11365 n2_12755_19645 n2_12804_19645 3.111111e-02
R11366 n2_12804_19645 n2_12896_19645 5.841270e-02
R11367 n2_12616_20674 n2_12708_20674 5.841270e-02
R11368 n2_12708_20674 n2_12755_20674 2.984127e-02
R11369 n2_12755_20674 n2_12804_20674 3.111111e-02
R11370 n2_12804_20674 n2_12896_20674 5.841270e-02
R11371 n2_12616_20770 n2_12708_20770 5.841270e-02
R11372 n2_12708_20770 n2_12755_20770 2.984127e-02
R11373 n2_12755_20770 n2_12804_20770 3.111111e-02
R11374 n2_12804_20770 n2_12896_20770 5.841270e-02
R11375 n2_12708_201 n2_12708_234 2.095238e-02
R11376 n2_12708_234 n2_12708_417 1.161905e-01
R11377 n2_12708_417 n2_12708_424 4.444444e-03
R11378 n2_12708_424 n2_12708_450 1.650794e-02
R11379 n2_12708_450 n2_12708_520 4.444444e-02
R11380 n2_12708_520 n2_12708_633 7.174603e-02
R11381 n2_12708_633 n2_12708_666 2.095238e-02
R11382 n2_12708_666 n2_12708_849 1.161905e-01
R11383 n2_12708_849 n2_12708_882 2.095238e-02
R11384 n2_12708_882 n2_12708_1065 1.161905e-01
R11385 n2_12708_1065 n2_12708_1098 2.095238e-02
R11386 n2_12708_1098 n2_12708_1281 1.161905e-01
R11387 n2_12708_1281 n2_12708_1314 2.095238e-02
R11388 n2_12708_1314 n2_12708_1497 1.161905e-01
R11389 n2_12708_1497 n2_12708_1530 2.095238e-02
R11390 n2_12708_1530 n2_12708_1549 1.206349e-02
R11391 n2_12708_1549 n2_12708_1645 6.095238e-02
R11392 n2_12708_1645 n2_12708_1713 4.317460e-02
R11393 n2_12708_1713 n2_12708_1746 2.095238e-02
R11394 n2_12708_1746 n2_12708_1783 2.349206e-02
R11395 n2_12708_1783 n2_12708_1929 9.269841e-02
R11396 n2_12708_1929 n2_12708_1962 2.095238e-02
R11397 n2_12708_1962 n2_12708_2145 1.161905e-01
R11398 n2_12708_2145 n2_12708_2178 2.095238e-02
R11399 n2_12708_2178 n2_12708_2361 1.161905e-01
R11400 n2_12708_2361 n2_12708_2394 2.095238e-02
R11401 n2_12708_2394 n2_12708_2431 2.349206e-02
R11402 n2_12708_2431 n2_12708_2577 9.269841e-02
R11403 n2_12708_2577 n2_12708_2610 2.095238e-02
R11404 n2_12708_2610 n2_12708_2674 4.063492e-02
R11405 n2_12708_2674 n2_12708_2770 6.095238e-02
R11406 n2_12708_2770 n2_12708_2793 1.460317e-02
R11407 n2_12708_2793 n2_12708_2826 2.095238e-02
R11408 n2_12708_2826 n2_12708_2863 2.349206e-02
R11409 n2_12708_2863 n2_12708_3009 9.269841e-02
R11410 n2_12708_3009 n2_12708_3042 2.095238e-02
R11411 n2_12708_3042 n2_12708_3225 1.161905e-01
R11412 n2_12708_3225 n2_12708_3258 2.095238e-02
R11413 n2_12708_3258 n2_12708_3441 1.161905e-01
R11414 n2_12708_3441 n2_12708_3474 2.095238e-02
R11415 n2_12708_3474 n2_12708_3511 2.349206e-02
R11416 n2_12708_3511 n2_12708_3657 9.269841e-02
R11417 n2_12708_3657 n2_12708_3690 2.095238e-02
R11418 n2_12708_3690 n2_12708_3799 6.920635e-02
R11419 n2_12708_3799 n2_12708_3873 4.698413e-02
R11420 n2_12708_3873 n2_12708_3895 1.396825e-02
R11421 n2_12708_3895 n2_12708_3906 6.984127e-03
R11422 n2_12708_3906 n2_12708_3943 2.349206e-02
R11423 n2_12708_3943 n2_12708_4089 9.269841e-02
R11424 n2_12708_4089 n2_12708_4122 2.095238e-02
R11425 n2_12708_4122 n2_12708_4159 2.349206e-02
R11426 n2_12708_4159 n2_12708_4305 9.269841e-02
R11427 n2_12708_4305 n2_12708_4338 2.095238e-02
R11428 n2_12708_4338 n2_12708_4521 1.161905e-01
R11429 n2_12708_4521 n2_12708_4554 2.095238e-02
R11430 n2_12708_4554 n2_12708_4591 2.349206e-02
R11431 n2_12708_4591 n2_12708_4737 9.269841e-02
R11432 n2_12708_4737 n2_12708_4770 2.095238e-02
R11433 n2_12708_4770 n2_12708_4924 9.777778e-02
R11434 n2_12708_4924 n2_12708_4953 1.841270e-02
R11435 n2_12708_4953 n2_12708_4986 2.095238e-02
R11436 n2_12708_4986 n2_12708_5020 2.158730e-02
R11437 n2_12708_5020 n2_12708_5023 1.904762e-03
R11438 n2_12708_5023 n2_12708_5169 9.269841e-02
R11439 n2_12708_5169 n2_12708_5202 2.095238e-02
R11440 n2_12708_5202 n2_12708_5239 2.349206e-02
R11441 n2_12708_5239 n2_12708_5385 9.269841e-02
R11442 n2_12708_5385 n2_12708_5418 2.095238e-02
R11443 n2_12708_5418 n2_12708_5601 1.161905e-01
R11444 n2_12708_5601 n2_12708_5634 2.095238e-02
R11445 n2_12708_5634 n2_12708_5671 2.349206e-02
R11446 n2_12708_5671 n2_12708_5817 9.269841e-02
R11447 n2_12708_5817 n2_12708_5850 2.095238e-02
R11448 n2_12708_5850 n2_12708_6033 1.161905e-01
R11449 n2_12708_6033 n2_12708_6049 1.015873e-02
R11450 n2_12708_6049 n2_12708_6066 1.079365e-02
R11451 n2_12708_6066 n2_12708_6145 5.015873e-02
R11452 n2_12708_6145 n2_12708_6249 6.603175e-02
R11453 n2_12708_6249 n2_12708_6282 2.095238e-02
R11454 n2_12708_6282 n2_12708_6319 2.349206e-02
R11455 n2_12708_6319 n2_12708_6465 9.269841e-02
R11456 n2_12708_6465 n2_12708_6498 2.095238e-02
R11457 n2_12708_6498 n2_12708_6681 1.161905e-01
R11458 n2_12708_6681 n2_12708_6714 2.095238e-02
R11459 n2_12708_6714 n2_12708_6751 2.349206e-02
R11460 n2_12708_6751 n2_12708_6897 9.269841e-02
R11461 n2_12708_6897 n2_12708_6930 2.095238e-02
R11462 n2_12708_6930 n2_12708_6967 2.349206e-02
R11463 n2_12708_6967 n2_12708_7113 9.269841e-02
R11464 n2_12708_7113 n2_12708_7146 2.095238e-02
R11465 n2_12708_7146 n2_12708_7174 1.777778e-02
R11466 n2_12708_7174 n2_12708_7178 2.539683e-03
R11467 n2_12708_7178 n2_12708_7270 5.841270e-02
R11468 n2_12708_7270 n2_12708_7329 3.746032e-02
R11469 n2_12708_7329 n2_12708_7362 2.095238e-02
R11470 n2_12708_7362 n2_12708_7399 2.349206e-02
R11471 n2_12708_7399 n2_12708_7545 9.269841e-02
R11472 n2_12708_7545 n2_12708_7578 2.095238e-02
R11473 n2_12708_7578 n2_12708_7761 1.161905e-01
R11474 n2_12708_7761 n2_12708_7794 2.095238e-02
R11475 n2_12708_7794 n2_12708_7831 2.349206e-02
R11476 n2_12708_7831 n2_12708_7977 9.269841e-02
R11477 n2_12708_7977 n2_12708_8010 2.095238e-02
R11478 n2_12708_8010 n2_12708_8193 1.161905e-01
R11479 n2_12708_8193 n2_12708_8226 2.095238e-02
R11480 n2_12708_8226 n2_12708_8299 4.634921e-02
R11481 n2_12708_8299 n2_12708_8395 6.095238e-02
R11482 n2_12708_8395 n2_12708_8409 8.888889e-03
R11483 n2_12708_8409 n2_12708_8442 2.095238e-02
R11484 n2_12708_12762 n2_12708_12799 2.349206e-02
R11485 n2_12708_12799 n2_12708_12895 6.095238e-02
R11486 n2_12708_12895 n2_12708_12945 3.174603e-02
R11487 n2_12708_12945 n2_12708_12978 2.095238e-02
R11488 n2_12708_12978 n2_12708_13161 1.161905e-01
R11489 n2_12708_13161 n2_12708_13194 2.095238e-02
R11490 n2_12708_13194 n2_12708_13377 1.161905e-01
R11491 n2_12708_13377 n2_12708_13410 2.095238e-02
R11492 n2_12708_13410 n2_12708_13593 1.161905e-01
R11493 n2_12708_13593 n2_12708_13626 2.095238e-02
R11494 n2_12708_13626 n2_12708_13663 2.349206e-02
R11495 n2_12708_13663 n2_12708_13809 9.269841e-02
R11496 n2_12708_13809 n2_12708_13842 2.095238e-02
R11497 n2_12708_13842 n2_12708_13924 5.206349e-02
R11498 n2_12708_13924 n2_12708_14020 6.095238e-02
R11499 n2_12708_14020 n2_12708_14025 3.174603e-03
R11500 n2_12708_14025 n2_12708_14058 2.095238e-02
R11501 n2_12708_14058 n2_12708_14079 1.333333e-02
R11502 n2_12708_14079 n2_12708_14241 1.028571e-01
R11503 n2_12708_14241 n2_12708_14274 2.095238e-02
R11504 n2_12708_14274 n2_12708_14457 1.161905e-01
R11505 n2_12708_14457 n2_12708_14490 2.095238e-02
R11506 n2_12708_14490 n2_12708_14673 1.161905e-01
R11507 n2_12708_14673 n2_12708_14706 2.095238e-02
R11508 n2_12708_14706 n2_12708_14727 1.333333e-02
R11509 n2_12708_14727 n2_12708_14889 1.028571e-01
R11510 n2_12708_14889 n2_12708_14922 2.095238e-02
R11511 n2_12708_14922 n2_12708_15049 8.063492e-02
R11512 n2_12708_15049 n2_12708_15105 3.555556e-02
R11513 n2_12708_15105 n2_12708_15138 2.095238e-02
R11514 n2_12708_15138 n2_12708_15145 4.444444e-03
R11515 n2_12708_15145 n2_12708_15321 1.117460e-01
R11516 n2_12708_15321 n2_12708_15354 2.095238e-02
R11517 n2_12708_15354 n2_12708_15368 8.888889e-03
R11518 n2_12708_15368 n2_12708_15537 1.073016e-01
R11519 n2_12708_15537 n2_12708_15570 2.095238e-02
R11520 n2_12708_15570 n2_12708_15753 1.161905e-01
R11521 n2_12708_15753 n2_12708_15786 2.095238e-02
R11522 n2_12708_15786 n2_12708_15800 8.888889e-03
R11523 n2_12708_15800 n2_12708_15807 4.444444e-03
R11524 n2_12708_15807 n2_12708_15969 1.028571e-01
R11525 n2_12708_15969 n2_12708_16002 2.095238e-02
R11526 n2_12708_16002 n2_12708_16174 1.092063e-01
R11527 n2_12708_16174 n2_12708_16185 6.984127e-03
R11528 n2_12708_16185 n2_12708_16218 2.095238e-02
R11529 n2_12708_16218 n2_12708_16270 3.301587e-02
R11530 n2_12708_16270 n2_12708_16401 8.317460e-02
R11531 n2_12708_16401 n2_12708_16434 2.095238e-02
R11532 n2_12708_16434 n2_12708_16448 8.888889e-03
R11533 n2_12708_16448 n2_12708_16617 1.073016e-01
R11534 n2_12708_16617 n2_12708_16650 2.095238e-02
R11535 n2_12708_16650 n2_12708_16833 1.161905e-01
R11536 n2_12708_16833 n2_12708_16866 2.095238e-02
R11537 n2_12708_16866 n2_12708_17049 1.161905e-01
R11538 n2_12708_17049 n2_12708_17082 2.095238e-02
R11539 n2_12708_17082 n2_12708_17096 8.888889e-03
R11540 n2_12708_17096 n2_12708_17103 4.444444e-03
R11541 n2_12708_17103 n2_12708_17265 1.028571e-01
R11542 n2_12708_17265 n2_12708_17298 2.095238e-02
R11543 n2_12708_17298 n2_12708_17299 6.349206e-04
R11544 n2_12708_17299 n2_12708_17395 6.095238e-02
R11545 n2_12708_17395 n2_12708_17481 5.460317e-02
R11546 n2_12708_17481 n2_12708_17514 2.095238e-02
R11547 n2_12708_17514 n2_12708_17528 8.888889e-03
R11548 n2_12708_17528 n2_12708_17697 1.073016e-01
R11549 n2_12708_17697 n2_12708_17730 2.095238e-02
R11550 n2_12708_17730 n2_12708_17913 1.161905e-01
R11551 n2_12708_17913 n2_12708_17946 2.095238e-02
R11552 n2_12708_17946 n2_12708_17983 2.349206e-02
R11553 n2_12708_17983 n2_12708_18129 9.269841e-02
R11554 n2_12708_18129 n2_12708_18162 2.095238e-02
R11555 n2_12708_18162 n2_12708_18176 8.888889e-03
R11556 n2_12708_18176 n2_12708_18183 4.444444e-03
R11557 n2_12708_18183 n2_12708_18345 1.028571e-01
R11558 n2_12708_18345 n2_12708_18378 2.095238e-02
R11559 n2_12708_18378 n2_12708_18424 2.920635e-02
R11560 n2_12708_18424 n2_12708_18520 6.095238e-02
R11561 n2_12708_18520 n2_12708_18561 2.603175e-02
R11562 n2_12708_18561 n2_12708_18594 2.095238e-02
R11563 n2_12708_18594 n2_12708_18608 8.888889e-03
R11564 n2_12708_18608 n2_12708_18777 1.073016e-01
R11565 n2_12708_18777 n2_12708_18810 2.095238e-02
R11566 n2_12708_18810 n2_12708_18993 1.161905e-01
R11567 n2_12708_18993 n2_12708_19026 2.095238e-02
R11568 n2_12708_19026 n2_12708_19209 1.161905e-01
R11569 n2_12708_19209 n2_12708_19242 2.095238e-02
R11570 n2_12708_19242 n2_12708_19256 8.888889e-03
R11571 n2_12708_19256 n2_12708_19263 4.444444e-03
R11572 n2_12708_19263 n2_12708_19425 1.028571e-01
R11573 n2_12708_19425 n2_12708_19458 2.095238e-02
R11574 n2_12708_19458 n2_12708_19549 5.777778e-02
R11575 n2_12708_19549 n2_12708_19641 5.841270e-02
R11576 n2_12708_19641 n2_12708_19645 2.539683e-03
R11577 n2_12708_19645 n2_12708_19674 1.841270e-02
R11578 n2_12708_19674 n2_12708_19857 1.161905e-01
R11579 n2_12708_19857 n2_12708_19890 2.095238e-02
R11580 n2_12708_19890 n2_12708_20073 1.161905e-01
R11581 n2_12708_20073 n2_12708_20106 2.095238e-02
R11582 n2_12708_20106 n2_12708_20289 1.161905e-01
R11583 n2_12708_20289 n2_12708_20322 2.095238e-02
R11584 n2_12708_20322 n2_12708_20505 1.161905e-01
R11585 n2_12708_20505 n2_12708_20538 2.095238e-02
R11586 n2_12708_20538 n2_12708_20674 8.634921e-02
R11587 n2_12708_20674 n2_12708_20721 2.984127e-02
R11588 n2_12708_20721 n2_12708_20754 2.095238e-02
R11589 n2_12708_20754 n2_12708_20770 1.015873e-02
R11590 n2_12708_20770 n2_12708_20937 1.060317e-01
R11591 n2_12708_20937 n2_12708_20970 2.095238e-02
R11592 n2_12804_201 n2_12804_234 2.095238e-02
R11593 n2_12804_234 n2_12804_417 1.161905e-01
R11594 n2_12804_417 n2_12804_424 4.444444e-03
R11595 n2_12804_424 n2_12804_450 1.650794e-02
R11596 n2_12804_450 n2_12804_520 4.444444e-02
R11597 n2_12804_520 n2_12804_633 7.174603e-02
R11598 n2_12804_633 n2_12804_666 2.095238e-02
R11599 n2_12804_666 n2_12804_849 1.161905e-01
R11600 n2_12804_849 n2_12804_882 2.095238e-02
R11601 n2_12804_882 n2_12804_1065 1.161905e-01
R11602 n2_12804_1065 n2_12804_1098 2.095238e-02
R11603 n2_12804_1098 n2_12804_1281 1.161905e-01
R11604 n2_12804_1281 n2_12804_1314 2.095238e-02
R11605 n2_12804_1314 n2_12804_1497 1.161905e-01
R11606 n2_12804_1497 n2_12804_1530 2.095238e-02
R11607 n2_12804_1530 n2_12804_1549 1.206349e-02
R11608 n2_12804_1549 n2_12804_1645 6.095238e-02
R11609 n2_12804_1645 n2_12804_1713 4.317460e-02
R11610 n2_12804_1713 n2_12804_1746 2.095238e-02
R11611 n2_12804_1746 n2_12804_1783 2.349206e-02
R11612 n2_12804_1783 n2_12804_1929 9.269841e-02
R11613 n2_12804_1929 n2_12804_1962 2.095238e-02
R11614 n2_12804_1962 n2_12804_2145 1.161905e-01
R11615 n2_12804_2145 n2_12804_2178 2.095238e-02
R11616 n2_12804_2178 n2_12804_2361 1.161905e-01
R11617 n2_12804_2361 n2_12804_2394 2.095238e-02
R11618 n2_12804_2394 n2_12804_2431 2.349206e-02
R11619 n2_12804_2431 n2_12804_2577 9.269841e-02
R11620 n2_12804_2577 n2_12804_2610 2.095238e-02
R11621 n2_12804_2610 n2_12804_2674 4.063492e-02
R11622 n2_12804_2674 n2_12804_2770 6.095238e-02
R11623 n2_12804_2770 n2_12804_2793 1.460317e-02
R11624 n2_12804_2793 n2_12804_2826 2.095238e-02
R11625 n2_12804_2826 n2_12804_2863 2.349206e-02
R11626 n2_12804_2863 n2_12804_3009 9.269841e-02
R11627 n2_12804_3009 n2_12804_3042 2.095238e-02
R11628 n2_12804_3042 n2_12804_3225 1.161905e-01
R11629 n2_12804_3225 n2_12804_3258 2.095238e-02
R11630 n2_12804_3258 n2_12804_3441 1.161905e-01
R11631 n2_12804_3441 n2_12804_3474 2.095238e-02
R11632 n2_12804_3474 n2_12804_3511 2.349206e-02
R11633 n2_12804_3511 n2_12804_3657 9.269841e-02
R11634 n2_12804_3657 n2_12804_3690 2.095238e-02
R11635 n2_12804_3690 n2_12804_3799 6.920635e-02
R11636 n2_12804_3799 n2_12804_3873 4.698413e-02
R11637 n2_12804_3873 n2_12804_3895 1.396825e-02
R11638 n2_12804_3895 n2_12804_3906 6.984127e-03
R11639 n2_12804_3906 n2_12804_3943 2.349206e-02
R11640 n2_12804_3943 n2_12804_4089 9.269841e-02
R11641 n2_12804_4089 n2_12804_4122 2.095238e-02
R11642 n2_12804_4122 n2_12804_4159 2.349206e-02
R11643 n2_12804_4159 n2_12804_4305 9.269841e-02
R11644 n2_12804_4305 n2_12804_4338 2.095238e-02
R11645 n2_12804_4338 n2_12804_4521 1.161905e-01
R11646 n2_12804_4521 n2_12804_4554 2.095238e-02
R11647 n2_12804_4554 n2_12804_4591 2.349206e-02
R11648 n2_12804_4591 n2_12804_4737 9.269841e-02
R11649 n2_12804_4737 n2_12804_4770 2.095238e-02
R11650 n2_12804_4770 n2_12804_4924 9.777778e-02
R11651 n2_12804_4924 n2_12804_4953 1.841270e-02
R11652 n2_12804_4953 n2_12804_4986 2.095238e-02
R11653 n2_12804_4986 n2_12804_5020 2.158730e-02
R11654 n2_12804_5020 n2_12804_5023 1.904762e-03
R11655 n2_12804_5023 n2_12804_5169 9.269841e-02
R11656 n2_12804_5169 n2_12804_5202 2.095238e-02
R11657 n2_12804_5202 n2_12804_5239 2.349206e-02
R11658 n2_12804_5239 n2_12804_5385 9.269841e-02
R11659 n2_12804_5385 n2_12804_5418 2.095238e-02
R11660 n2_12804_5418 n2_12804_5601 1.161905e-01
R11661 n2_12804_5601 n2_12804_5634 2.095238e-02
R11662 n2_12804_5634 n2_12804_5671 2.349206e-02
R11663 n2_12804_5671 n2_12804_5817 9.269841e-02
R11664 n2_12804_5817 n2_12804_5850 2.095238e-02
R11665 n2_12804_5850 n2_12804_6033 1.161905e-01
R11666 n2_12804_6033 n2_12804_6049 1.015873e-02
R11667 n2_12804_6049 n2_12804_6066 1.079365e-02
R11668 n2_12804_6066 n2_12804_6145 5.015873e-02
R11669 n2_12804_6145 n2_12804_6249 6.603175e-02
R11670 n2_12804_6249 n2_12804_6282 2.095238e-02
R11671 n2_12804_6282 n2_12804_6319 2.349206e-02
R11672 n2_12804_6319 n2_12804_6465 9.269841e-02
R11673 n2_12804_6465 n2_12804_6498 2.095238e-02
R11674 n2_12804_6498 n2_12804_6681 1.161905e-01
R11675 n2_12804_6681 n2_12804_6714 2.095238e-02
R11676 n2_12804_6714 n2_12804_6751 2.349206e-02
R11677 n2_12804_6751 n2_12804_6897 9.269841e-02
R11678 n2_12804_6897 n2_12804_6930 2.095238e-02
R11679 n2_12804_6930 n2_12804_6967 2.349206e-02
R11680 n2_12804_6967 n2_12804_7113 9.269841e-02
R11681 n2_12804_7113 n2_12804_7146 2.095238e-02
R11682 n2_12804_7146 n2_12804_7174 1.777778e-02
R11683 n2_12804_7174 n2_12804_7178 2.539683e-03
R11684 n2_12804_7178 n2_12804_7270 5.841270e-02
R11685 n2_12804_7270 n2_12804_7329 3.746032e-02
R11686 n2_12804_7329 n2_12804_7362 2.095238e-02
R11687 n2_12804_7362 n2_12804_7399 2.349206e-02
R11688 n2_12804_7399 n2_12804_7545 9.269841e-02
R11689 n2_12804_7545 n2_12804_7578 2.095238e-02
R11690 n2_12804_7578 n2_12804_7761 1.161905e-01
R11691 n2_12804_7761 n2_12804_7794 2.095238e-02
R11692 n2_12804_7794 n2_12804_7831 2.349206e-02
R11693 n2_12804_7831 n2_12804_7977 9.269841e-02
R11694 n2_12804_7977 n2_12804_8010 2.095238e-02
R11695 n2_12804_8010 n2_12804_8193 1.161905e-01
R11696 n2_12804_8193 n2_12804_8226 2.095238e-02
R11697 n2_12804_8226 n2_12804_8299 4.634921e-02
R11698 n2_12804_8299 n2_12804_8395 6.095238e-02
R11699 n2_12804_8395 n2_12804_8409 8.888889e-03
R11700 n2_12804_8409 n2_12804_8442 2.095238e-02
R11701 n2_12804_8442 n2_12804_8625 1.161905e-01
R11702 n2_12804_8625 n2_12804_8658 2.095238e-02
R11703 n2_12804_8658 n2_12804_8695 2.349206e-02
R11704 n2_12804_8695 n2_12804_8841 9.269841e-02
R11705 n2_12804_8841 n2_12804_8874 2.095238e-02
R11706 n2_12804_8874 n2_12804_8911 2.349206e-02
R11707 n2_12804_8911 n2_12804_9057 9.269841e-02
R11708 n2_12804_9057 n2_12804_9090 2.095238e-02
R11709 n2_12804_9090 n2_12804_9273 1.161905e-01
R11710 n2_12804_9273 n2_12804_9306 2.095238e-02
R11711 n2_12804_9705 n2_12804_9738 2.095238e-02
R11712 n2_12804_9738 n2_12804_9775 2.349206e-02
R11713 n2_12804_9775 n2_12804_9921 9.269841e-02
R11714 n2_12804_9921 n2_12804_9954 2.095238e-02
R11715 n2_12804_9954 n2_12804_9991 2.349206e-02
R11716 n2_12804_9991 n2_12804_10137 9.269841e-02
R11717 n2_12804_10137 n2_12804_10170 2.095238e-02
R11718 n2_12804_10170 n2_12804_10353 1.161905e-01
R11719 n2_12804_10353 n2_12804_10386 2.095238e-02
R11720 n2_12804_10386 n2_12804_10549 1.034921e-01
R11721 n2_12804_10549 n2_12804_10569 1.269841e-02
R11722 n2_12804_10569 n2_12804_10602 2.095238e-02
R11723 n2_12804_10602 n2_12804_10645 2.730159e-02
R11724 n2_12804_10645 n2_12804_10785 8.888889e-02
R11725 n2_12804_10785 n2_12804_10818 2.095238e-02
R11726 n2_12804_10818 n2_12804_10832 8.888889e-03
R11727 n2_12804_10832 n2_12804_11001 1.073016e-01
R11728 n2_12804_11001 n2_12804_11034 2.095238e-02
R11729 n2_12804_11034 n2_12804_11048 8.888889e-03
R11730 n2_12804_11048 n2_12804_11217 1.073016e-01
R11731 n2_12804_11217 n2_12804_11250 2.095238e-02
R11732 n2_12804_11250 n2_12804_11433 1.161905e-01
R11733 n2_12804_11433 n2_12804_11466 2.095238e-02
R11734 n2_12804_11865 n2_12804_11898 2.095238e-02
R11735 n2_12804_11898 n2_12804_11912 8.888889e-03
R11736 n2_12804_11912 n2_12804_12081 1.073016e-01
R11737 n2_12804_12081 n2_12804_12114 2.095238e-02
R11738 n2_12804_12114 n2_12804_12128 8.888889e-03
R11739 n2_12804_12128 n2_12804_12297 1.073016e-01
R11740 n2_12804_12297 n2_12804_12330 2.095238e-02
R11741 n2_12804_12330 n2_12804_12513 1.161905e-01
R11742 n2_12804_12513 n2_12804_12546 2.095238e-02
R11743 n2_12804_12546 n2_12804_12729 1.161905e-01
R11744 n2_12804_12729 n2_12804_12762 2.095238e-02
R11745 n2_12804_12762 n2_12804_12799 2.349206e-02
R11746 n2_12804_12799 n2_12804_12895 6.095238e-02
R11747 n2_12804_12895 n2_12804_12945 3.174603e-02
R11748 n2_12804_12945 n2_12804_12978 2.095238e-02
R11749 n2_12804_12978 n2_12804_13161 1.161905e-01
R11750 n2_12804_13161 n2_12804_13194 2.095238e-02
R11751 n2_12804_13194 n2_12804_13377 1.161905e-01
R11752 n2_12804_13377 n2_12804_13410 2.095238e-02
R11753 n2_12804_13410 n2_12804_13593 1.161905e-01
R11754 n2_12804_13593 n2_12804_13626 2.095238e-02
R11755 n2_12804_13626 n2_12804_13663 2.349206e-02
R11756 n2_12804_13663 n2_12804_13809 9.269841e-02
R11757 n2_12804_13809 n2_12804_13842 2.095238e-02
R11758 n2_12804_13842 n2_12804_13924 5.206349e-02
R11759 n2_12804_13924 n2_12804_14020 6.095238e-02
R11760 n2_12804_14020 n2_12804_14025 3.174603e-03
R11761 n2_12804_14025 n2_12804_14058 2.095238e-02
R11762 n2_12804_14058 n2_12804_14079 1.333333e-02
R11763 n2_12804_14079 n2_12804_14241 1.028571e-01
R11764 n2_12804_14241 n2_12804_14274 2.095238e-02
R11765 n2_12804_14274 n2_12804_14457 1.161905e-01
R11766 n2_12804_14457 n2_12804_14490 2.095238e-02
R11767 n2_12804_14490 n2_12804_14673 1.161905e-01
R11768 n2_12804_14673 n2_12804_14706 2.095238e-02
R11769 n2_12804_14706 n2_12804_14727 1.333333e-02
R11770 n2_12804_14727 n2_12804_14889 1.028571e-01
R11771 n2_12804_14889 n2_12804_14922 2.095238e-02
R11772 n2_12804_14922 n2_12804_15049 8.063492e-02
R11773 n2_12804_15049 n2_12804_15105 3.555556e-02
R11774 n2_12804_15105 n2_12804_15138 2.095238e-02
R11775 n2_12804_15138 n2_12804_15145 4.444444e-03
R11776 n2_12804_15145 n2_12804_15321 1.117460e-01
R11777 n2_12804_15321 n2_12804_15354 2.095238e-02
R11778 n2_12804_15354 n2_12804_15368 8.888889e-03
R11779 n2_12804_15368 n2_12804_15537 1.073016e-01
R11780 n2_12804_15537 n2_12804_15570 2.095238e-02
R11781 n2_12804_15570 n2_12804_15753 1.161905e-01
R11782 n2_12804_15753 n2_12804_15786 2.095238e-02
R11783 n2_12804_15786 n2_12804_15800 8.888889e-03
R11784 n2_12804_15800 n2_12804_15807 4.444444e-03
R11785 n2_12804_15807 n2_12804_15969 1.028571e-01
R11786 n2_12804_15969 n2_12804_16002 2.095238e-02
R11787 n2_12804_16002 n2_12804_16174 1.092063e-01
R11788 n2_12804_16174 n2_12804_16185 6.984127e-03
R11789 n2_12804_16185 n2_12804_16218 2.095238e-02
R11790 n2_12804_16218 n2_12804_16270 3.301587e-02
R11791 n2_12804_16270 n2_12804_16401 8.317460e-02
R11792 n2_12804_16401 n2_12804_16434 2.095238e-02
R11793 n2_12804_16434 n2_12804_16448 8.888889e-03
R11794 n2_12804_16448 n2_12804_16617 1.073016e-01
R11795 n2_12804_16617 n2_12804_16650 2.095238e-02
R11796 n2_12804_16650 n2_12804_16833 1.161905e-01
R11797 n2_12804_16833 n2_12804_16866 2.095238e-02
R11798 n2_12804_16866 n2_12804_17049 1.161905e-01
R11799 n2_12804_17049 n2_12804_17082 2.095238e-02
R11800 n2_12804_17082 n2_12804_17096 8.888889e-03
R11801 n2_12804_17096 n2_12804_17103 4.444444e-03
R11802 n2_12804_17103 n2_12804_17265 1.028571e-01
R11803 n2_12804_17265 n2_12804_17298 2.095238e-02
R11804 n2_12804_17298 n2_12804_17299 6.349206e-04
R11805 n2_12804_17299 n2_12804_17395 6.095238e-02
R11806 n2_12804_17395 n2_12804_17481 5.460317e-02
R11807 n2_12804_17481 n2_12804_17514 2.095238e-02
R11808 n2_12804_17514 n2_12804_17528 8.888889e-03
R11809 n2_12804_17528 n2_12804_17697 1.073016e-01
R11810 n2_12804_17697 n2_12804_17730 2.095238e-02
R11811 n2_12804_17730 n2_12804_17913 1.161905e-01
R11812 n2_12804_17913 n2_12804_17946 2.095238e-02
R11813 n2_12804_17946 n2_12804_17983 2.349206e-02
R11814 n2_12804_17983 n2_12804_18129 9.269841e-02
R11815 n2_12804_18129 n2_12804_18162 2.095238e-02
R11816 n2_12804_18162 n2_12804_18176 8.888889e-03
R11817 n2_12804_18176 n2_12804_18183 4.444444e-03
R11818 n2_12804_18183 n2_12804_18345 1.028571e-01
R11819 n2_12804_18345 n2_12804_18378 2.095238e-02
R11820 n2_12804_18378 n2_12804_18424 2.920635e-02
R11821 n2_12804_18424 n2_12804_18520 6.095238e-02
R11822 n2_12804_18520 n2_12804_18561 2.603175e-02
R11823 n2_12804_18561 n2_12804_18594 2.095238e-02
R11824 n2_12804_18594 n2_12804_18608 8.888889e-03
R11825 n2_12804_18608 n2_12804_18777 1.073016e-01
R11826 n2_12804_18777 n2_12804_18810 2.095238e-02
R11827 n2_12804_18810 n2_12804_18993 1.161905e-01
R11828 n2_12804_18993 n2_12804_19026 2.095238e-02
R11829 n2_12804_19026 n2_12804_19209 1.161905e-01
R11830 n2_12804_19209 n2_12804_19242 2.095238e-02
R11831 n2_12804_19242 n2_12804_19256 8.888889e-03
R11832 n2_12804_19256 n2_12804_19263 4.444444e-03
R11833 n2_12804_19263 n2_12804_19425 1.028571e-01
R11834 n2_12804_19425 n2_12804_19458 2.095238e-02
R11835 n2_12804_19458 n2_12804_19549 5.777778e-02
R11836 n2_12804_19549 n2_12804_19641 5.841270e-02
R11837 n2_12804_19641 n2_12804_19645 2.539683e-03
R11838 n2_12804_19645 n2_12804_19674 1.841270e-02
R11839 n2_12804_19674 n2_12804_19857 1.161905e-01
R11840 n2_12804_19857 n2_12804_19890 2.095238e-02
R11841 n2_12804_19890 n2_12804_20073 1.161905e-01
R11842 n2_12804_20073 n2_12804_20106 2.095238e-02
R11843 n2_12804_20106 n2_12804_20289 1.161905e-01
R11844 n2_12804_20289 n2_12804_20322 2.095238e-02
R11845 n2_12804_20322 n2_12804_20505 1.161905e-01
R11846 n2_12804_20505 n2_12804_20538 2.095238e-02
R11847 n2_12804_20538 n2_12804_20674 8.634921e-02
R11848 n2_12804_20674 n2_12804_20721 2.984127e-02
R11849 n2_12804_20721 n2_12804_20754 2.095238e-02
R11850 n2_12804_20754 n2_12804_20770 1.015873e-02
R11851 n2_12804_20770 n2_12804_20937 1.060317e-01
R11852 n2_12804_20937 n2_12804_20970 2.095238e-02
R11853 n2_12896_201 n2_12896_234 2.095238e-02
R11854 n2_12896_234 n2_12896_417 1.161905e-01
R11855 n2_12896_417 n2_12896_424 4.444444e-03
R11856 n2_12896_424 n2_12896_450 1.650794e-02
R11857 n2_12896_520 n2_12896_633 7.174603e-02
R11858 n2_12896_633 n2_12896_666 2.095238e-02
R11859 n2_12896_666 n2_12896_849 1.161905e-01
R11860 n2_12896_849 n2_12896_882 2.095238e-02
R11861 n2_12896_882 n2_12896_1065 1.161905e-01
R11862 n2_12896_1065 n2_12896_1098 2.095238e-02
R11863 n2_12896_1098 n2_12896_1281 1.161905e-01
R11864 n2_12896_1281 n2_12896_1314 2.095238e-02
R11865 n2_12896_1314 n2_12896_1497 1.161905e-01
R11866 n2_12896_1497 n2_12896_1530 2.095238e-02
R11867 n2_12896_1530 n2_12896_1549 1.206349e-02
R11868 n2_12896_1645 n2_12896_1713 4.317460e-02
R11869 n2_12896_1713 n2_12896_1746 2.095238e-02
R11870 n2_12896_1746 n2_12896_1783 2.349206e-02
R11871 n2_12896_1783 n2_12896_1929 9.269841e-02
R11872 n2_12896_1929 n2_12896_1962 2.095238e-02
R11873 n2_12896_1962 n2_12896_2145 1.161905e-01
R11874 n2_12896_2145 n2_12896_2178 2.095238e-02
R11875 n2_12896_2178 n2_12896_2361 1.161905e-01
R11876 n2_12896_2361 n2_12896_2394 2.095238e-02
R11877 n2_12896_2394 n2_12896_2431 2.349206e-02
R11878 n2_12896_2431 n2_12896_2577 9.269841e-02
R11879 n2_12896_2577 n2_12896_2610 2.095238e-02
R11880 n2_12896_2610 n2_12896_2674 4.063492e-02
R11881 n2_12896_2770 n2_12896_2793 1.460317e-02
R11882 n2_12896_2793 n2_12896_2826 2.095238e-02
R11883 n2_12896_2826 n2_12896_2863 2.349206e-02
R11884 n2_12896_2863 n2_12896_3009 9.269841e-02
R11885 n2_12896_3009 n2_12896_3042 2.095238e-02
R11886 n2_12896_3042 n2_12896_3225 1.161905e-01
R11887 n2_12896_3225 n2_12896_3258 2.095238e-02
R11888 n2_12896_3258 n2_12896_3441 1.161905e-01
R11889 n2_12896_3441 n2_12896_3474 2.095238e-02
R11890 n2_12896_3474 n2_12896_3511 2.349206e-02
R11891 n2_12896_3511 n2_12896_3657 9.269841e-02
R11892 n2_12896_3657 n2_12896_3690 2.095238e-02
R11893 n2_12896_3690 n2_12896_3799 6.920635e-02
R11894 n2_12896_3873 n2_12896_3895 1.396825e-02
R11895 n2_12896_3895 n2_12896_3906 6.984127e-03
R11896 n2_12896_3906 n2_12896_3943 2.349206e-02
R11897 n2_12896_3943 n2_12896_4089 9.269841e-02
R11898 n2_12896_4089 n2_12896_4122 2.095238e-02
R11899 n2_12896_4122 n2_12896_4159 2.349206e-02
R11900 n2_12896_4159 n2_12896_4305 9.269841e-02
R11901 n2_12896_4305 n2_12896_4338 2.095238e-02
R11902 n2_12896_4338 n2_12896_4521 1.161905e-01
R11903 n2_12896_4521 n2_12896_4554 2.095238e-02
R11904 n2_12896_4554 n2_12896_4591 2.349206e-02
R11905 n2_12896_4591 n2_12896_4737 9.269841e-02
R11906 n2_12896_4737 n2_12896_4770 2.095238e-02
R11907 n2_12896_4770 n2_12896_4924 9.777778e-02
R11908 n2_12896_4924 n2_12896_4953 1.841270e-02
R11909 n2_12896_5020 n2_12896_5023 1.904762e-03
R11910 n2_12896_5023 n2_12896_5169 9.269841e-02
R11911 n2_12896_5169 n2_12896_5202 2.095238e-02
R11912 n2_12896_5202 n2_12896_5239 2.349206e-02
R11913 n2_12896_5239 n2_12896_5385 9.269841e-02
R11914 n2_12896_5385 n2_12896_5418 2.095238e-02
R11915 n2_12896_5418 n2_12896_5601 1.161905e-01
R11916 n2_12896_5601 n2_12896_5634 2.095238e-02
R11917 n2_12896_5634 n2_12896_5671 2.349206e-02
R11918 n2_12896_5671 n2_12896_5817 9.269841e-02
R11919 n2_12896_5817 n2_12896_5850 2.095238e-02
R11920 n2_12896_5850 n2_12896_6033 1.161905e-01
R11921 n2_12896_6033 n2_12896_6049 1.015873e-02
R11922 n2_12896_6049 n2_12896_6066 1.079365e-02
R11923 n2_12896_6145 n2_12896_6249 6.603175e-02
R11924 n2_12896_6249 n2_12896_6282 2.095238e-02
R11925 n2_12896_6282 n2_12896_6319 2.349206e-02
R11926 n2_12896_6319 n2_12896_6465 9.269841e-02
R11927 n2_12896_6465 n2_12896_6498 2.095238e-02
R11928 n2_12896_6498 n2_12896_6681 1.161905e-01
R11929 n2_12896_6681 n2_12896_6714 2.095238e-02
R11930 n2_12896_6714 n2_12896_6751 2.349206e-02
R11931 n2_12896_6751 n2_12896_6897 9.269841e-02
R11932 n2_12896_6897 n2_12896_6930 2.095238e-02
R11933 n2_12896_6930 n2_12896_6967 2.349206e-02
R11934 n2_12896_6967 n2_12896_7113 9.269841e-02
R11935 n2_12896_7113 n2_12896_7146 2.095238e-02
R11936 n2_12896_7146 n2_12896_7174 1.777778e-02
R11937 n2_12896_7174 n2_12896_7178 2.539683e-03
R11938 n2_12896_7270 n2_12896_7329 3.746032e-02
R11939 n2_12896_7329 n2_12896_7362 2.095238e-02
R11940 n2_12896_7362 n2_12896_7399 2.349206e-02
R11941 n2_12896_7399 n2_12896_7545 9.269841e-02
R11942 n2_12896_7545 n2_12896_7578 2.095238e-02
R11943 n2_12896_7578 n2_12896_7761 1.161905e-01
R11944 n2_12896_7761 n2_12896_7794 2.095238e-02
R11945 n2_12896_7794 n2_12896_7831 2.349206e-02
R11946 n2_12896_7831 n2_12896_7977 9.269841e-02
R11947 n2_12896_7977 n2_12896_8010 2.095238e-02
R11948 n2_12896_8010 n2_12896_8193 1.161905e-01
R11949 n2_12896_8193 n2_12896_8226 2.095238e-02
R11950 n2_12896_8226 n2_12896_8299 4.634921e-02
R11951 n2_12896_12895 n2_12896_12945 3.174603e-02
R11952 n2_12896_12945 n2_12896_12978 2.095238e-02
R11953 n2_12896_12978 n2_12896_13161 1.161905e-01
R11954 n2_12896_13161 n2_12896_13194 2.095238e-02
R11955 n2_12896_13194 n2_12896_13377 1.161905e-01
R11956 n2_12896_13377 n2_12896_13410 2.095238e-02
R11957 n2_12896_13410 n2_12896_13593 1.161905e-01
R11958 n2_12896_13593 n2_12896_13626 2.095238e-02
R11959 n2_12896_13626 n2_12896_13663 2.349206e-02
R11960 n2_12896_13663 n2_12896_13809 9.269841e-02
R11961 n2_12896_13809 n2_12896_13842 2.095238e-02
R11962 n2_12896_13842 n2_12896_13924 5.206349e-02
R11963 n2_12896_14020 n2_12896_14025 3.174603e-03
R11964 n2_12896_14025 n2_12896_14058 2.095238e-02
R11965 n2_12896_14058 n2_12896_14079 1.333333e-02
R11966 n2_12896_14079 n2_12896_14241 1.028571e-01
R11967 n2_12896_14241 n2_12896_14274 2.095238e-02
R11968 n2_12896_14274 n2_12896_14457 1.161905e-01
R11969 n2_12896_14457 n2_12896_14490 2.095238e-02
R11970 n2_12896_14490 n2_12896_14673 1.161905e-01
R11971 n2_12896_14673 n2_12896_14706 2.095238e-02
R11972 n2_12896_14706 n2_12896_14727 1.333333e-02
R11973 n2_12896_14727 n2_12896_14889 1.028571e-01
R11974 n2_12896_14889 n2_12896_14922 2.095238e-02
R11975 n2_12896_14922 n2_12896_15049 8.063492e-02
R11976 n2_12896_15138 n2_12896_15145 4.444444e-03
R11977 n2_12896_15145 n2_12896_15321 1.117460e-01
R11978 n2_12896_15321 n2_12896_15354 2.095238e-02
R11979 n2_12896_15354 n2_12896_15368 8.888889e-03
R11980 n2_12896_15368 n2_12896_15537 1.073016e-01
R11981 n2_12896_15537 n2_12896_15570 2.095238e-02
R11982 n2_12896_15570 n2_12896_15753 1.161905e-01
R11983 n2_12896_15753 n2_12896_15786 2.095238e-02
R11984 n2_12896_15786 n2_12896_15800 8.888889e-03
R11985 n2_12896_15800 n2_12896_15807 4.444444e-03
R11986 n2_12896_15807 n2_12896_15969 1.028571e-01
R11987 n2_12896_15969 n2_12896_16002 2.095238e-02
R11988 n2_12896_16002 n2_12896_16174 1.092063e-01
R11989 n2_12896_16174 n2_12896_16185 6.984127e-03
R11990 n2_12896_16270 n2_12896_16401 8.317460e-02
R11991 n2_12896_16401 n2_12896_16434 2.095238e-02
R11992 n2_12896_16434 n2_12896_16448 8.888889e-03
R11993 n2_12896_16448 n2_12896_16617 1.073016e-01
R11994 n2_12896_16617 n2_12896_16650 2.095238e-02
R11995 n2_12896_16650 n2_12896_16833 1.161905e-01
R11996 n2_12896_16833 n2_12896_16866 2.095238e-02
R11997 n2_12896_16866 n2_12896_17049 1.161905e-01
R11998 n2_12896_17049 n2_12896_17082 2.095238e-02
R11999 n2_12896_17082 n2_12896_17096 8.888889e-03
R12000 n2_12896_17096 n2_12896_17103 4.444444e-03
R12001 n2_12896_17103 n2_12896_17265 1.028571e-01
R12002 n2_12896_17265 n2_12896_17298 2.095238e-02
R12003 n2_12896_17298 n2_12896_17299 6.349206e-04
R12004 n2_12896_17395 n2_12896_17481 5.460317e-02
R12005 n2_12896_17481 n2_12896_17514 2.095238e-02
R12006 n2_12896_17514 n2_12896_17528 8.888889e-03
R12007 n2_12896_17528 n2_12896_17697 1.073016e-01
R12008 n2_12896_17697 n2_12896_17730 2.095238e-02
R12009 n2_12896_17730 n2_12896_17913 1.161905e-01
R12010 n2_12896_17913 n2_12896_17946 2.095238e-02
R12011 n2_12896_17946 n2_12896_17983 2.349206e-02
R12012 n2_12896_17983 n2_12896_18129 9.269841e-02
R12013 n2_12896_18129 n2_12896_18162 2.095238e-02
R12014 n2_12896_18162 n2_12896_18176 8.888889e-03
R12015 n2_12896_18176 n2_12896_18183 4.444444e-03
R12016 n2_12896_18183 n2_12896_18345 1.028571e-01
R12017 n2_12896_18345 n2_12896_18378 2.095238e-02
R12018 n2_12896_18378 n2_12896_18424 2.920635e-02
R12019 n2_12896_18520 n2_12896_18561 2.603175e-02
R12020 n2_12896_18561 n2_12896_18594 2.095238e-02
R12021 n2_12896_18594 n2_12896_18608 8.888889e-03
R12022 n2_12896_18608 n2_12896_18777 1.073016e-01
R12023 n2_12896_18777 n2_12896_18810 2.095238e-02
R12024 n2_12896_18810 n2_12896_18993 1.161905e-01
R12025 n2_12896_18993 n2_12896_19026 2.095238e-02
R12026 n2_12896_19026 n2_12896_19209 1.161905e-01
R12027 n2_12896_19209 n2_12896_19242 2.095238e-02
R12028 n2_12896_19242 n2_12896_19256 8.888889e-03
R12029 n2_12896_19256 n2_12896_19263 4.444444e-03
R12030 n2_12896_19263 n2_12896_19425 1.028571e-01
R12031 n2_12896_19425 n2_12896_19458 2.095238e-02
R12032 n2_12896_19458 n2_12896_19549 5.777778e-02
R12033 n2_12896_19641 n2_12896_19645 2.539683e-03
R12034 n2_12896_19645 n2_12896_19674 1.841270e-02
R12035 n2_12896_19674 n2_12896_19857 1.161905e-01
R12036 n2_12896_19857 n2_12896_19890 2.095238e-02
R12037 n2_12896_19890 n2_12896_20073 1.161905e-01
R12038 n2_12896_20073 n2_12896_20106 2.095238e-02
R12039 n2_12896_20106 n2_12896_20289 1.161905e-01
R12040 n2_12896_20289 n2_12896_20322 2.095238e-02
R12041 n2_12896_20322 n2_12896_20505 1.161905e-01
R12042 n2_12896_20505 n2_12896_20538 2.095238e-02
R12043 n2_12896_20538 n2_12896_20674 8.634921e-02
R12044 n2_12896_20754 n2_12896_20770 1.015873e-02
R12045 n2_12896_20770 n2_12896_20937 1.060317e-01
R12046 n2_12896_20937 n2_12896_20970 2.095238e-02
R12047 n2_13741_7329 n2_13741_7362 2.095238e-02
R12048 n2_13741_7362 n2_13741_7545 1.161905e-01
R12049 n2_13741_7545 n2_13741_7578 2.095238e-02
R12050 n2_13741_7578 n2_13741_7761 1.161905e-01
R12051 n2_13741_7761 n2_13741_7794 2.095238e-02
R12052 n2_13741_7794 n2_13741_7831 2.349206e-02
R12053 n2_13741_7831 n2_13741_7977 9.269841e-02
R12054 n2_13741_7977 n2_13741_8010 2.095238e-02
R12055 n2_13741_8010 n2_13741_8193 1.161905e-01
R12056 n2_13741_8193 n2_13741_8226 2.095238e-02
R12057 n2_13741_8226 n2_13741_8299 4.634921e-02
R12058 n2_13741_8395 n2_13741_8409 8.888889e-03
R12059 n2_13741_8409 n2_13741_8442 2.095238e-02
R12060 n2_13741_8442 n2_13741_8625 1.161905e-01
R12061 n2_13741_8625 n2_13741_8658 2.095238e-02
R12062 n2_13741_8658 n2_13741_8695 2.349206e-02
R12063 n2_13741_8695 n2_13741_8841 9.269841e-02
R12064 n2_13741_8841 n2_13741_8874 2.095238e-02
R12065 n2_13741_8874 n2_13741_8911 2.349206e-02
R12066 n2_13741_8911 n2_13741_9057 9.269841e-02
R12067 n2_13741_9057 n2_13741_9090 2.095238e-02
R12068 n2_13741_9090 n2_13741_9273 1.161905e-01
R12069 n2_13741_9273 n2_13741_9306 2.095238e-02
R12070 n2_13741_9306 n2_13741_9489 1.161905e-01
R12071 n2_13741_9489 n2_13741_9522 2.095238e-02
R12072 n2_13741_9522 n2_13741_9705 1.161905e-01
R12073 n2_13741_9705 n2_13741_9738 2.095238e-02
R12074 n2_13741_9738 n2_13741_9775 2.349206e-02
R12075 n2_13741_9775 n2_13741_9921 9.269841e-02
R12076 n2_13741_9921 n2_13741_9954 2.095238e-02
R12077 n2_13741_9954 n2_13741_9991 2.349206e-02
R12078 n2_13741_9991 n2_13741_10137 9.269841e-02
R12079 n2_13741_10137 n2_13741_10170 2.095238e-02
R12080 n2_13741_10170 n2_13741_10353 1.161905e-01
R12081 n2_13741_10353 n2_13741_10386 2.095238e-02
R12082 n2_13741_10386 n2_13741_10549 1.034921e-01
R12083 n2_13741_10549 n2_13741_10569 1.269841e-02
R12084 n2_13741_10645 n2_13741_10785 8.888889e-02
R12085 n2_13741_10785 n2_13741_10818 2.095238e-02
R12086 n2_13741_10818 n2_13741_10832 8.888889e-03
R12087 n2_13741_10832 n2_13741_11001 1.073016e-01
R12088 n2_13741_11001 n2_13741_11034 2.095238e-02
R12089 n2_13741_11034 n2_13741_11048 8.888889e-03
R12090 n2_13741_11048 n2_13741_11217 1.073016e-01
R12091 n2_13741_11217 n2_13741_11250 2.095238e-02
R12092 n2_13741_11250 n2_13741_11433 1.161905e-01
R12093 n2_13741_11433 n2_13741_11466 2.095238e-02
R12094 n2_13741_11466 n2_13741_11649 1.161905e-01
R12095 n2_13741_11649 n2_13741_11682 2.095238e-02
R12096 n2_13741_11682 n2_13741_11865 1.161905e-01
R12097 n2_13741_11865 n2_13741_11898 2.095238e-02
R12098 n2_13741_11898 n2_13741_11912 8.888889e-03
R12099 n2_13741_11912 n2_13741_12081 1.073016e-01
R12100 n2_13741_12081 n2_13741_12114 2.095238e-02
R12101 n2_13741_12114 n2_13741_12128 8.888889e-03
R12102 n2_13741_12128 n2_13741_12297 1.073016e-01
R12103 n2_13741_12297 n2_13741_12330 2.095238e-02
R12104 n2_13741_12330 n2_13741_12513 1.161905e-01
R12105 n2_13741_12513 n2_13741_12546 2.095238e-02
R12106 n2_13741_12546 n2_13741_12729 1.161905e-01
R12107 n2_13741_12729 n2_13741_12762 2.095238e-02
R12108 n2_13741_12762 n2_13741_12776 8.888889e-03
R12109 n2_13741_12776 n2_13741_12799 1.460317e-02
R12110 n2_13741_12895 n2_13741_12945 3.174603e-02
R12111 n2_13741_12945 n2_13741_12978 2.095238e-02
R12112 n2_13741_12978 n2_13741_12992 8.888889e-03
R12113 n2_13741_12992 n2_13741_13161 1.073016e-01
R12114 n2_13741_13161 n2_13741_13194 2.095238e-02
R12115 n2_13741_13194 n2_13741_13377 1.161905e-01
R12116 n2_13741_13377 n2_13741_13410 2.095238e-02
R12117 n2_13741_13410 n2_13741_13423 8.253968e-03
R12118 n2_13741_13423 n2_13741_13593 1.079365e-01
R12119 n2_13741_13593 n2_13741_13626 2.095238e-02
R12120 n2_13741_13626 n2_13741_13809 1.161905e-01
R12121 n2_13741_13809 n2_13741_13842 2.095238e-02
R12122 n2_13741_8299 n2_13880_8299 8.825397e-02
R12123 n2_13880_8299 n2_13929_8299 3.111111e-02
R12124 n2_13741_8395 n2_13880_8395 8.825397e-02
R12125 n2_13880_8395 n2_13929_8395 3.111111e-02
R12126 n2_13741_10549 n2_13880_10549 8.825397e-02
R12127 n2_13880_10549 n2_13929_10549 3.111111e-02
R12128 n2_13741_10645 n2_13880_10645 8.825397e-02
R12129 n2_13880_10645 n2_13929_10645 3.111111e-02
R12130 n2_13741_12799 n2_13880_12799 8.825397e-02
R12131 n2_13880_12799 n2_13929_12799 3.111111e-02
R12132 n2_13741_12895 n2_13880_12895 8.825397e-02
R12133 n2_13880_12895 n2_13929_12895 3.111111e-02
R12134 n2_13929_7329 n2_13929_7362 2.095238e-02
R12135 n2_13929_7362 n2_13929_7545 1.161905e-01
R12136 n2_13929_7545 n2_13929_7578 2.095238e-02
R12137 n2_13929_7578 n2_13929_7761 1.161905e-01
R12138 n2_13929_7761 n2_13929_7794 2.095238e-02
R12139 n2_13929_7794 n2_13929_7831 2.349206e-02
R12140 n2_13929_7831 n2_13929_7977 9.269841e-02
R12141 n2_13929_7977 n2_13929_8010 2.095238e-02
R12142 n2_13929_8010 n2_13929_8193 1.161905e-01
R12143 n2_13929_8193 n2_13929_8226 2.095238e-02
R12144 n2_13929_8226 n2_13929_8299 4.634921e-02
R12145 n2_13929_8299 n2_13929_8395 6.095238e-02
R12146 n2_13929_8395 n2_13929_8409 8.888889e-03
R12147 n2_13929_8409 n2_13929_8442 2.095238e-02
R12148 n2_13929_8442 n2_13929_8625 1.161905e-01
R12149 n2_13929_8625 n2_13929_8658 2.095238e-02
R12150 n2_13929_8658 n2_13929_8695 2.349206e-02
R12151 n2_13929_8695 n2_13929_8841 9.269841e-02
R12152 n2_13929_8841 n2_13929_8874 2.095238e-02
R12153 n2_13929_8874 n2_13929_8911 2.349206e-02
R12154 n2_13929_8911 n2_13929_9057 9.269841e-02
R12155 n2_13929_9057 n2_13929_9090 2.095238e-02
R12156 n2_13929_9090 n2_13929_9273 1.161905e-01
R12157 n2_13929_9273 n2_13929_9306 2.095238e-02
R12158 n2_13929_9705 n2_13929_9738 2.095238e-02
R12159 n2_13929_9738 n2_13929_9775 2.349206e-02
R12160 n2_13929_9775 n2_13929_9921 9.269841e-02
R12161 n2_13929_9921 n2_13929_9954 2.095238e-02
R12162 n2_13929_9954 n2_13929_9991 2.349206e-02
R12163 n2_13929_9991 n2_13929_10137 9.269841e-02
R12164 n2_13929_10137 n2_13929_10170 2.095238e-02
R12165 n2_13929_10170 n2_13929_10353 1.161905e-01
R12166 n2_13929_10353 n2_13929_10386 2.095238e-02
R12167 n2_13929_10386 n2_13929_10549 1.034921e-01
R12168 n2_13929_10549 n2_13929_10569 1.269841e-02
R12169 n2_13929_10569 n2_13929_10602 2.095238e-02
R12170 n2_13929_10602 n2_13929_10645 2.730159e-02
R12171 n2_13929_10645 n2_13929_10785 8.888889e-02
R12172 n2_13929_10785 n2_13929_10818 2.095238e-02
R12173 n2_13929_10818 n2_13929_10832 8.888889e-03
R12174 n2_13929_10832 n2_13929_11001 1.073016e-01
R12175 n2_13929_11001 n2_13929_11034 2.095238e-02
R12176 n2_13929_11034 n2_13929_11048 8.888889e-03
R12177 n2_13929_11048 n2_13929_11217 1.073016e-01
R12178 n2_13929_11217 n2_13929_11250 2.095238e-02
R12179 n2_13929_11250 n2_13929_11433 1.161905e-01
R12180 n2_13929_11433 n2_13929_11466 2.095238e-02
R12181 n2_13929_11865 n2_13929_11898 2.095238e-02
R12182 n2_13929_11898 n2_13929_11912 8.888889e-03
R12183 n2_13929_11912 n2_13929_12081 1.073016e-01
R12184 n2_13929_12081 n2_13929_12114 2.095238e-02
R12185 n2_13929_12114 n2_13929_12128 8.888889e-03
R12186 n2_13929_12128 n2_13929_12297 1.073016e-01
R12187 n2_13929_12297 n2_13929_12330 2.095238e-02
R12188 n2_13929_12330 n2_13929_12513 1.161905e-01
R12189 n2_13929_12513 n2_13929_12546 2.095238e-02
R12190 n2_13929_12546 n2_13929_12729 1.161905e-01
R12191 n2_13929_12729 n2_13929_12762 2.095238e-02
R12192 n2_13929_12762 n2_13929_12776 8.888889e-03
R12193 n2_13929_12776 n2_13929_12799 1.460317e-02
R12194 n2_13929_12799 n2_13929_12895 6.095238e-02
R12195 n2_13929_12895 n2_13929_12945 3.174603e-02
R12196 n2_13929_12945 n2_13929_12978 2.095238e-02
R12197 n2_13929_12978 n2_13929_12992 8.888889e-03
R12198 n2_13929_12992 n2_13929_13161 1.073016e-01
R12199 n2_13929_13161 n2_13929_13194 2.095238e-02
R12200 n2_13929_13194 n2_13929_13377 1.161905e-01
R12201 n2_13929_13377 n2_13929_13410 2.095238e-02
R12202 n2_13929_13410 n2_13929_13423 8.253968e-03
R12203 n2_13929_13423 n2_13929_13593 1.079365e-01
R12204 n2_13929_13593 n2_13929_13626 2.095238e-02
R12205 n2_13929_13626 n2_13929_13809 1.161905e-01
R12206 n2_13929_13809 n2_13929_13842 2.095238e-02
R12207 n2_14866_201 n2_14866_234 2.095238e-02
R12208 n2_14866_234 n2_14866_417 1.161905e-01
R12209 n2_14866_417 n2_14866_424 4.444444e-03
R12210 n2_14866_424 n2_14866_450 1.650794e-02
R12211 n2_14866_520 n2_14866_633 7.174603e-02
R12212 n2_14866_633 n2_14866_666 2.095238e-02
R12213 n2_14866_666 n2_14866_849 1.161905e-01
R12214 n2_14866_849 n2_14866_882 2.095238e-02
R12215 n2_14866_882 n2_14866_1065 1.161905e-01
R12216 n2_14866_1065 n2_14866_1098 2.095238e-02
R12217 n2_14866_1098 n2_14866_1281 1.161905e-01
R12218 n2_14866_1281 n2_14866_1314 2.095238e-02
R12219 n2_14866_1314 n2_14866_1497 1.161905e-01
R12220 n2_14866_1497 n2_14866_1530 2.095238e-02
R12221 n2_14866_1530 n2_14866_1549 1.206349e-02
R12222 n2_14866_1645 n2_14866_1713 4.317460e-02
R12223 n2_14866_1713 n2_14866_1746 2.095238e-02
R12224 n2_14866_1746 n2_14866_1783 2.349206e-02
R12225 n2_14866_1783 n2_14866_1929 9.269841e-02
R12226 n2_14866_1929 n2_14866_1962 2.095238e-02
R12227 n2_14866_1962 n2_14866_2145 1.161905e-01
R12228 n2_14866_2145 n2_14866_2178 2.095238e-02
R12229 n2_14866_2178 n2_14866_2361 1.161905e-01
R12230 n2_14866_2361 n2_14866_2394 2.095238e-02
R12231 n2_14866_2394 n2_14866_2431 2.349206e-02
R12232 n2_14866_2431 n2_14866_2577 9.269841e-02
R12233 n2_14866_2577 n2_14866_2610 2.095238e-02
R12234 n2_14866_2610 n2_14866_2674 4.063492e-02
R12235 n2_14866_2770 n2_14866_2793 1.460317e-02
R12236 n2_14866_2793 n2_14866_2826 2.095238e-02
R12237 n2_14866_2826 n2_14866_2863 2.349206e-02
R12238 n2_14866_2863 n2_14866_3009 9.269841e-02
R12239 n2_14866_3009 n2_14866_3042 2.095238e-02
R12240 n2_14866_3042 n2_14866_3225 1.161905e-01
R12241 n2_14866_3225 n2_14866_3258 2.095238e-02
R12242 n2_14866_3258 n2_14866_3295 2.349206e-02
R12243 n2_14866_3295 n2_14866_3441 9.269841e-02
R12244 n2_14866_3441 n2_14866_3474 2.095238e-02
R12245 n2_14866_3474 n2_14866_3511 2.349206e-02
R12246 n2_14866_3511 n2_14866_3657 9.269841e-02
R12247 n2_14866_3657 n2_14866_3690 2.095238e-02
R12248 n2_14866_3690 n2_14866_3799 6.920635e-02
R12249 n2_14866_3873 n2_14866_3895 1.396825e-02
R12250 n2_14866_3895 n2_14866_3906 6.984127e-03
R12251 n2_14866_3906 n2_14866_3943 2.349206e-02
R12252 n2_14866_3943 n2_14866_4089 9.269841e-02
R12253 n2_14866_4089 n2_14866_4122 2.095238e-02
R12254 n2_14866_4122 n2_14866_4159 2.349206e-02
R12255 n2_14866_4159 n2_14866_4305 9.269841e-02
R12256 n2_14866_4305 n2_14866_4338 2.095238e-02
R12257 n2_14866_4338 n2_14866_4375 2.349206e-02
R12258 n2_14866_4375 n2_14866_4521 9.269841e-02
R12259 n2_14866_4521 n2_14866_4554 2.095238e-02
R12260 n2_14866_4554 n2_14866_4591 2.349206e-02
R12261 n2_14866_4591 n2_14866_4737 9.269841e-02
R12262 n2_14866_4737 n2_14866_4770 2.095238e-02
R12263 n2_14866_4770 n2_14866_4807 2.349206e-02
R12264 n2_14866_4807 n2_14866_4924 7.428571e-02
R12265 n2_14866_4924 n2_14866_4953 1.841270e-02
R12266 n2_14866_5020 n2_14866_5169 9.460317e-02
R12267 n2_14866_5169 n2_14866_5202 2.095238e-02
R12268 n2_14866_5202 n2_14866_5239 2.349206e-02
R12269 n2_14866_5239 n2_14866_5385 9.269841e-02
R12270 n2_14866_5385 n2_14866_5418 2.095238e-02
R12271 n2_14866_5418 n2_14866_5455 2.349206e-02
R12272 n2_14866_5455 n2_14866_5601 9.269841e-02
R12273 n2_14866_5601 n2_14866_5634 2.095238e-02
R12274 n2_14866_5634 n2_14866_5671 2.349206e-02
R12275 n2_14866_5671 n2_14866_5817 9.269841e-02
R12276 n2_14866_5817 n2_14866_5850 2.095238e-02
R12277 n2_14866_5850 n2_14866_6033 1.161905e-01
R12278 n2_14866_6033 n2_14866_6049 1.015873e-02
R12279 n2_14866_6049 n2_14866_6066 1.079365e-02
R12280 n2_14866_6145 n2_14866_6249 6.603175e-02
R12281 n2_14866_6249 n2_14866_6282 2.095238e-02
R12282 n2_14866_6282 n2_14866_6319 2.349206e-02
R12283 n2_14866_6319 n2_14866_6465 9.269841e-02
R12284 n2_14866_6465 n2_14866_6498 2.095238e-02
R12285 n2_14866_6498 n2_14866_6535 2.349206e-02
R12286 n2_14866_6535 n2_14866_6681 9.269841e-02
R12287 n2_14866_6681 n2_14866_6714 2.095238e-02
R12288 n2_14866_6714 n2_14866_6897 1.161905e-01
R12289 n2_14866_6897 n2_14866_6930 2.095238e-02
R12290 n2_14866_6930 n2_14866_7113 1.161905e-01
R12291 n2_14866_7113 n2_14866_7146 2.095238e-02
R12292 n2_14866_7146 n2_14866_7329 1.161905e-01
R12293 n2_14866_7329 n2_14866_7362 2.095238e-02
R12294 n2_14866_7362 n2_14866_7545 1.161905e-01
R12295 n2_14866_7545 n2_14866_7578 2.095238e-02
R12296 n2_14866_7578 n2_14866_7761 1.161905e-01
R12297 n2_14866_7761 n2_14866_7794 2.095238e-02
R12298 n2_14866_7794 n2_14866_7831 2.349206e-02
R12299 n2_14866_7831 n2_14866_7977 9.269841e-02
R12300 n2_14866_7977 n2_14866_8010 2.095238e-02
R12301 n2_14866_8010 n2_14866_8193 1.161905e-01
R12302 n2_14866_8193 n2_14866_8226 2.095238e-02
R12303 n2_14866_8226 n2_14866_8299 4.634921e-02
R12304 n2_14866_8395 n2_14866_8409 8.888889e-03
R12305 n2_14866_8409 n2_14866_8442 2.095238e-02
R12306 n2_14866_8442 n2_14866_8625 1.161905e-01
R12307 n2_14866_8625 n2_14866_8658 2.095238e-02
R12308 n2_14866_8658 n2_14866_8841 1.161905e-01
R12309 n2_14866_8841 n2_14866_8874 2.095238e-02
R12310 n2_14866_8874 n2_14866_8911 2.349206e-02
R12311 n2_14866_8911 n2_14866_9057 9.269841e-02
R12312 n2_14866_9057 n2_14866_9090 2.095238e-02
R12313 n2_14866_9090 n2_14866_9273 1.161905e-01
R12314 n2_14866_9273 n2_14866_9306 2.095238e-02
R12315 n2_14866_9306 n2_14866_9489 1.161905e-01
R12316 n2_14866_9489 n2_14866_9522 2.095238e-02
R12317 n2_14866_9522 n2_14866_9705 1.161905e-01
R12318 n2_14866_9705 n2_14866_9738 2.095238e-02
R12319 n2_14866_9738 n2_14866_9921 1.161905e-01
R12320 n2_14866_9921 n2_14866_9954 2.095238e-02
R12321 n2_14866_9954 n2_14866_9991 2.349206e-02
R12322 n2_14866_9991 n2_14866_10137 9.269841e-02
R12323 n2_14866_10137 n2_14866_10170 2.095238e-02
R12324 n2_14866_10170 n2_14866_10353 1.161905e-01
R12325 n2_14866_10353 n2_14866_10386 2.095238e-02
R12326 n2_14866_10386 n2_14866_10549 1.034921e-01
R12327 n2_14866_10549 n2_14866_10569 1.269841e-02
R12328 n2_14866_10645 n2_14866_10785 8.888889e-02
R12329 n2_14866_10785 n2_14866_10818 2.095238e-02
R12330 n2_14866_10818 n2_14866_11001 1.161905e-01
R12331 n2_14866_11001 n2_14866_11034 2.095238e-02
R12332 n2_14866_11034 n2_14866_11048 8.888889e-03
R12333 n2_14866_11048 n2_14866_11217 1.073016e-01
R12334 n2_14866_11217 n2_14866_11250 2.095238e-02
R12335 n2_14866_11250 n2_14866_11433 1.161905e-01
R12336 n2_14866_11433 n2_14866_11466 2.095238e-02
R12337 n2_14866_11466 n2_14866_11649 1.161905e-01
R12338 n2_14866_11649 n2_14866_11682 2.095238e-02
R12339 n2_14866_11682 n2_14866_11865 1.161905e-01
R12340 n2_14866_11865 n2_14866_11898 2.095238e-02
R12341 n2_14866_11898 n2_14866_12081 1.161905e-01
R12342 n2_14866_12081 n2_14866_12114 2.095238e-02
R12343 n2_14866_12114 n2_14866_12128 8.888889e-03
R12344 n2_14866_12128 n2_14866_12135 4.444444e-03
R12345 n2_14866_12135 n2_14866_12297 1.028571e-01
R12346 n2_14866_12297 n2_14866_12330 2.095238e-02
R12347 n2_14866_12330 n2_14866_12513 1.161905e-01
R12348 n2_14866_12513 n2_14866_12546 2.095238e-02
R12349 n2_14866_12546 n2_14866_12729 1.161905e-01
R12350 n2_14866_12729 n2_14866_12762 2.095238e-02
R12351 n2_14866_12762 n2_14866_12776 8.888889e-03
R12352 n2_14866_12776 n2_14866_12799 1.460317e-02
R12353 n2_14866_12895 n2_14866_12945 3.174603e-02
R12354 n2_14866_12945 n2_14866_12978 2.095238e-02
R12355 n2_14866_12978 n2_14866_12992 8.888889e-03
R12356 n2_14866_12992 n2_14866_13161 1.073016e-01
R12357 n2_14866_13161 n2_14866_13194 2.095238e-02
R12358 n2_14866_13194 n2_14866_13377 1.161905e-01
R12359 n2_14866_13377 n2_14866_13410 2.095238e-02
R12360 n2_14866_13410 n2_14866_13423 8.253968e-03
R12361 n2_14866_13423 n2_14866_13593 1.079365e-01
R12362 n2_14866_13593 n2_14866_13626 2.095238e-02
R12363 n2_14866_13626 n2_14866_13809 1.161905e-01
R12364 n2_14866_13809 n2_14866_13842 2.095238e-02
R12365 n2_14866_13842 n2_14866_14025 1.161905e-01
R12366 n2_14866_14025 n2_14866_14058 2.095238e-02
R12367 n2_14866_14058 n2_14866_14241 1.161905e-01
R12368 n2_14866_14241 n2_14866_14274 2.095238e-02
R12369 n2_14866_14274 n2_14866_14457 1.161905e-01
R12370 n2_14866_14457 n2_14866_14490 2.095238e-02
R12371 n2_14866_14490 n2_14866_14511 1.333333e-02
R12372 n2_14866_14511 n2_14866_14673 1.028571e-01
R12373 n2_14866_14673 n2_14866_14706 2.095238e-02
R12374 n2_14866_14706 n2_14866_14889 1.161905e-01
R12375 n2_14866_14889 n2_14866_14922 2.095238e-02
R12376 n2_14866_14922 n2_14866_14943 1.333333e-02
R12377 n2_14866_14943 n2_14866_15049 6.730159e-02
R12378 n2_14866_15138 n2_14866_15145 4.444444e-03
R12379 n2_14866_15145 n2_14866_15159 8.888889e-03
R12380 n2_14866_15159 n2_14866_15321 1.028571e-01
R12381 n2_14866_15321 n2_14866_15354 2.095238e-02
R12382 n2_14866_15354 n2_14866_15368 8.888889e-03
R12383 n2_14866_15368 n2_14866_15537 1.073016e-01
R12384 n2_14866_15537 n2_14866_15570 2.095238e-02
R12385 n2_14866_15570 n2_14866_15584 8.888889e-03
R12386 n2_14866_15584 n2_14866_15753 1.073016e-01
R12387 n2_14866_15753 n2_14866_15786 2.095238e-02
R12388 n2_14866_15786 n2_14866_15800 8.888889e-03
R12389 n2_14866_15800 n2_14866_15969 1.073016e-01
R12390 n2_14866_15969 n2_14866_16002 2.095238e-02
R12391 n2_14866_16002 n2_14866_16174 1.092063e-01
R12392 n2_14866_16174 n2_14866_16185 6.984127e-03
R12393 n2_14866_16270 n2_14866_16401 8.317460e-02
R12394 n2_14866_16401 n2_14866_16434 2.095238e-02
R12395 n2_14866_16434 n2_14866_16448 8.888889e-03
R12396 n2_14866_16448 n2_14866_16617 1.073016e-01
R12397 n2_14866_16617 n2_14866_16650 2.095238e-02
R12398 n2_14866_16650 n2_14866_16687 2.349206e-02
R12399 n2_14866_16687 n2_14866_16833 9.269841e-02
R12400 n2_14866_16833 n2_14866_16866 2.095238e-02
R12401 n2_14866_16866 n2_14866_17049 1.161905e-01
R12402 n2_14866_17049 n2_14866_17082 2.095238e-02
R12403 n2_14866_17082 n2_14866_17096 8.888889e-03
R12404 n2_14866_17096 n2_14866_17265 1.073016e-01
R12405 n2_14866_17265 n2_14866_17298 2.095238e-02
R12406 n2_14866_17298 n2_14866_17299 6.349206e-04
R12407 n2_14866_17395 n2_14866_17481 5.460317e-02
R12408 n2_14866_17481 n2_14866_17514 2.095238e-02
R12409 n2_14866_17514 n2_14866_17528 8.888889e-03
R12410 n2_14866_17528 n2_14866_17697 1.073016e-01
R12411 n2_14866_17697 n2_14866_17730 2.095238e-02
R12412 n2_14866_17730 n2_14866_17913 1.161905e-01
R12413 n2_14866_17913 n2_14866_17946 2.095238e-02
R12414 n2_14866_17946 n2_14866_17983 2.349206e-02
R12415 n2_14866_17983 n2_14866_18129 9.269841e-02
R12416 n2_14866_18129 n2_14866_18162 2.095238e-02
R12417 n2_14866_18162 n2_14866_18176 8.888889e-03
R12418 n2_14866_18176 n2_14866_18345 1.073016e-01
R12419 n2_14866_18345 n2_14866_18378 2.095238e-02
R12420 n2_14866_18378 n2_14866_18424 2.920635e-02
R12421 n2_14866_18520 n2_14866_18561 2.603175e-02
R12422 n2_14866_18561 n2_14866_18594 2.095238e-02
R12423 n2_14866_18594 n2_14866_18608 8.888889e-03
R12424 n2_14866_18608 n2_14866_18777 1.073016e-01
R12425 n2_14866_18777 n2_14866_18810 2.095238e-02
R12426 n2_14866_18810 n2_14866_18993 1.161905e-01
R12427 n2_14866_18993 n2_14866_19026 2.095238e-02
R12428 n2_14866_19026 n2_14866_19209 1.161905e-01
R12429 n2_14866_19209 n2_14866_19242 2.095238e-02
R12430 n2_14866_19242 n2_14866_19256 8.888889e-03
R12431 n2_14866_19256 n2_14866_19263 4.444444e-03
R12432 n2_14866_19263 n2_14866_19425 1.028571e-01
R12433 n2_14866_19425 n2_14866_19458 2.095238e-02
R12434 n2_14866_19458 n2_14866_19549 5.777778e-02
R12435 n2_14866_19641 n2_14866_19645 2.539683e-03
R12436 n2_14866_19645 n2_14866_19674 1.841270e-02
R12437 n2_14866_19674 n2_14866_19857 1.161905e-01
R12438 n2_14866_19857 n2_14866_19890 2.095238e-02
R12439 n2_14866_19890 n2_14866_20073 1.161905e-01
R12440 n2_14866_20073 n2_14866_20106 2.095238e-02
R12441 n2_14866_20106 n2_14866_20289 1.161905e-01
R12442 n2_14866_20289 n2_14866_20322 2.095238e-02
R12443 n2_14866_20322 n2_14866_20505 1.161905e-01
R12444 n2_14866_20505 n2_14866_20538 2.095238e-02
R12445 n2_14866_20538 n2_14866_20674 8.634921e-02
R12446 n2_14866_20754 n2_14866_20770 1.015873e-02
R12447 n2_14866_20770 n2_14866_20937 1.060317e-01
R12448 n2_14866_20937 n2_14866_20970 2.095238e-02
R12449 n2_14866_6145 n2_14958_6145 5.841270e-02
R12450 n2_14958_6145 n2_15005_6145 2.984127e-02
R12451 n2_15005_6145 n2_15054_6145 3.111111e-02
R12452 n2_14866_8299 n2_15005_8299 8.825397e-02
R12453 n2_15005_8299 n2_15054_8299 3.111111e-02
R12454 n2_14866_8395 n2_15005_8395 8.825397e-02
R12455 n2_15005_8395 n2_15054_8395 3.111111e-02
R12456 n2_14866_10549 n2_15005_10549 8.825397e-02
R12457 n2_15005_10549 n2_15054_10549 3.111111e-02
R12458 n2_14866_10645 n2_15005_10645 8.825397e-02
R12459 n2_15005_10645 n2_15054_10645 3.111111e-02
R12460 n2_14866_12799 n2_15005_12799 8.825397e-02
R12461 n2_15005_12799 n2_15054_12799 3.111111e-02
R12462 n2_14866_12895 n2_15005_12895 8.825397e-02
R12463 n2_15005_12895 n2_15054_12895 3.111111e-02
R12464 n2_14866_15049 n2_14958_15049 5.841270e-02
R12465 n2_14958_15049 n2_15005_15049 2.984127e-02
R12466 n2_15005_15049 n2_15054_15049 3.111111e-02
R12467 n2_14866_424 n2_14958_424 5.841270e-02
R12468 n2_14958_424 n2_15005_424 2.984127e-02
R12469 n2_15005_424 n2_15054_424 3.111111e-02
R12470 n2_15054_424 n2_15146_424 5.841270e-02
R12471 n2_14866_520 n2_14958_520 5.841270e-02
R12472 n2_14958_520 n2_15005_520 2.984127e-02
R12473 n2_15005_520 n2_15054_520 3.111111e-02
R12474 n2_15054_520 n2_15146_520 5.841270e-02
R12475 n2_14866_1549 n2_14958_1549 5.841270e-02
R12476 n2_14958_1549 n2_15005_1549 2.984127e-02
R12477 n2_15005_1549 n2_15054_1549 3.111111e-02
R12478 n2_15054_1549 n2_15146_1549 5.841270e-02
R12479 n2_14866_1645 n2_14958_1645 5.841270e-02
R12480 n2_14958_1645 n2_15005_1645 2.984127e-02
R12481 n2_15005_1645 n2_15054_1645 3.111111e-02
R12482 n2_15054_1645 n2_15146_1645 5.841270e-02
R12483 n2_14866_2674 n2_14958_2674 5.841270e-02
R12484 n2_14958_2674 n2_15005_2674 2.984127e-02
R12485 n2_15005_2674 n2_15054_2674 3.111111e-02
R12486 n2_15054_2674 n2_15146_2674 5.841270e-02
R12487 n2_14866_2770 n2_14958_2770 5.841270e-02
R12488 n2_14958_2770 n2_15005_2770 2.984127e-02
R12489 n2_15005_2770 n2_15054_2770 3.111111e-02
R12490 n2_15054_2770 n2_15146_2770 5.841270e-02
R12491 n2_14866_3799 n2_14958_3799 5.841270e-02
R12492 n2_14958_3799 n2_15005_3799 2.984127e-02
R12493 n2_15005_3799 n2_15054_3799 3.111111e-02
R12494 n2_15054_3799 n2_15146_3799 5.841270e-02
R12495 n2_14866_3895 n2_14958_3895 5.841270e-02
R12496 n2_14958_3895 n2_15005_3895 2.984127e-02
R12497 n2_15005_3895 n2_15054_3895 3.111111e-02
R12498 n2_15054_3895 n2_15146_3895 5.841270e-02
R12499 n2_14866_4924 n2_14958_4924 5.841270e-02
R12500 n2_14958_4924 n2_15005_4924 2.984127e-02
R12501 n2_15005_4924 n2_15054_4924 3.111111e-02
R12502 n2_15054_4924 n2_15146_4924 5.841270e-02
R12503 n2_14866_5020 n2_14958_5020 5.841270e-02
R12504 n2_14958_5020 n2_15005_5020 2.984127e-02
R12505 n2_15005_5020 n2_15054_5020 3.111111e-02
R12506 n2_15054_5020 n2_15146_5020 5.841270e-02
R12507 n2_14866_6049 n2_14958_6049 5.841270e-02
R12508 n2_14958_6049 n2_15005_6049 2.984127e-02
R12509 n2_15005_6049 n2_15054_6049 3.111111e-02
R12510 n2_15054_6049 n2_15146_6049 5.841270e-02
R12511 n2_14866_15145 n2_14958_15145 5.841270e-02
R12512 n2_14958_15145 n2_15005_15145 2.984127e-02
R12513 n2_15005_15145 n2_15054_15145 3.111111e-02
R12514 n2_15054_15145 n2_15146_15145 5.841270e-02
R12515 n2_14866_16174 n2_14958_16174 5.841270e-02
R12516 n2_14958_16174 n2_15005_16174 2.984127e-02
R12517 n2_15005_16174 n2_15054_16174 3.111111e-02
R12518 n2_15054_16174 n2_15146_16174 5.841270e-02
R12519 n2_14866_16270 n2_14958_16270 5.841270e-02
R12520 n2_14958_16270 n2_15005_16270 2.984127e-02
R12521 n2_15005_16270 n2_15054_16270 3.111111e-02
R12522 n2_15054_16270 n2_15146_16270 5.841270e-02
R12523 n2_14866_17299 n2_14958_17299 5.841270e-02
R12524 n2_14958_17299 n2_15005_17299 2.984127e-02
R12525 n2_15005_17299 n2_15054_17299 3.111111e-02
R12526 n2_15054_17299 n2_15146_17299 5.841270e-02
R12527 n2_14866_17395 n2_14958_17395 5.841270e-02
R12528 n2_14958_17395 n2_15005_17395 2.984127e-02
R12529 n2_15005_17395 n2_15054_17395 3.111111e-02
R12530 n2_15054_17395 n2_15146_17395 5.841270e-02
R12531 n2_14866_18424 n2_14958_18424 5.841270e-02
R12532 n2_14958_18424 n2_15005_18424 2.984127e-02
R12533 n2_15005_18424 n2_15054_18424 3.111111e-02
R12534 n2_15054_18424 n2_15146_18424 5.841270e-02
R12535 n2_14866_18520 n2_14958_18520 5.841270e-02
R12536 n2_14958_18520 n2_15005_18520 2.984127e-02
R12537 n2_15005_18520 n2_15054_18520 3.111111e-02
R12538 n2_15054_18520 n2_15146_18520 5.841270e-02
R12539 n2_14866_19549 n2_14958_19549 5.841270e-02
R12540 n2_14958_19549 n2_15005_19549 2.984127e-02
R12541 n2_15005_19549 n2_15054_19549 3.111111e-02
R12542 n2_15054_19549 n2_15146_19549 5.841270e-02
R12543 n2_14866_19645 n2_14958_19645 5.841270e-02
R12544 n2_14958_19645 n2_15005_19645 2.984127e-02
R12545 n2_15005_19645 n2_15054_19645 3.111111e-02
R12546 n2_15054_19645 n2_15146_19645 5.841270e-02
R12547 n2_14866_20674 n2_14958_20674 5.841270e-02
R12548 n2_14958_20674 n2_15005_20674 2.984127e-02
R12549 n2_15005_20674 n2_15054_20674 3.111111e-02
R12550 n2_15054_20674 n2_15146_20674 5.841270e-02
R12551 n2_14866_20770 n2_14958_20770 5.841270e-02
R12552 n2_14958_20770 n2_15005_20770 2.984127e-02
R12553 n2_15005_20770 n2_15054_20770 3.111111e-02
R12554 n2_15054_20770 n2_15146_20770 5.841270e-02
R12555 n2_14958_201 n2_14958_234 2.095238e-02
R12556 n2_14958_234 n2_14958_417 1.161905e-01
R12557 n2_14958_417 n2_14958_424 4.444444e-03
R12558 n2_14958_424 n2_14958_450 1.650794e-02
R12559 n2_14958_450 n2_14958_520 4.444444e-02
R12560 n2_14958_520 n2_14958_633 7.174603e-02
R12561 n2_14958_633 n2_14958_666 2.095238e-02
R12562 n2_14958_666 n2_14958_849 1.161905e-01
R12563 n2_14958_849 n2_14958_882 2.095238e-02
R12564 n2_14958_882 n2_14958_1065 1.161905e-01
R12565 n2_14958_1065 n2_14958_1098 2.095238e-02
R12566 n2_14958_1098 n2_14958_1281 1.161905e-01
R12567 n2_14958_1281 n2_14958_1314 2.095238e-02
R12568 n2_14958_1314 n2_14958_1497 1.161905e-01
R12569 n2_14958_1497 n2_14958_1530 2.095238e-02
R12570 n2_14958_1530 n2_14958_1549 1.206349e-02
R12571 n2_14958_1549 n2_14958_1645 6.095238e-02
R12572 n2_14958_1645 n2_14958_1713 4.317460e-02
R12573 n2_14958_1713 n2_14958_1746 2.095238e-02
R12574 n2_14958_1746 n2_14958_1783 2.349206e-02
R12575 n2_14958_1783 n2_14958_1929 9.269841e-02
R12576 n2_14958_1929 n2_14958_1962 2.095238e-02
R12577 n2_14958_1962 n2_14958_2145 1.161905e-01
R12578 n2_14958_2145 n2_14958_2178 2.095238e-02
R12579 n2_14958_2178 n2_14958_2361 1.161905e-01
R12580 n2_14958_2361 n2_14958_2394 2.095238e-02
R12581 n2_14958_2394 n2_14958_2431 2.349206e-02
R12582 n2_14958_2431 n2_14958_2577 9.269841e-02
R12583 n2_14958_2577 n2_14958_2610 2.095238e-02
R12584 n2_14958_2610 n2_14958_2674 4.063492e-02
R12585 n2_14958_2674 n2_14958_2770 6.095238e-02
R12586 n2_14958_2770 n2_14958_2793 1.460317e-02
R12587 n2_14958_2793 n2_14958_2826 2.095238e-02
R12588 n2_14958_2826 n2_14958_2863 2.349206e-02
R12589 n2_14958_2863 n2_14958_3009 9.269841e-02
R12590 n2_14958_3009 n2_14958_3042 2.095238e-02
R12591 n2_14958_3042 n2_14958_3225 1.161905e-01
R12592 n2_14958_3225 n2_14958_3258 2.095238e-02
R12593 n2_14958_3258 n2_14958_3295 2.349206e-02
R12594 n2_14958_3295 n2_14958_3441 9.269841e-02
R12595 n2_14958_3441 n2_14958_3474 2.095238e-02
R12596 n2_14958_3474 n2_14958_3511 2.349206e-02
R12597 n2_14958_3511 n2_14958_3657 9.269841e-02
R12598 n2_14958_3657 n2_14958_3690 2.095238e-02
R12599 n2_14958_3690 n2_14958_3799 6.920635e-02
R12600 n2_14958_3799 n2_14958_3873 4.698413e-02
R12601 n2_14958_3873 n2_14958_3895 1.396825e-02
R12602 n2_14958_3895 n2_14958_3906 6.984127e-03
R12603 n2_14958_3906 n2_14958_3943 2.349206e-02
R12604 n2_14958_3943 n2_14958_4089 9.269841e-02
R12605 n2_14958_4089 n2_14958_4122 2.095238e-02
R12606 n2_14958_4122 n2_14958_4159 2.349206e-02
R12607 n2_14958_4159 n2_14958_4305 9.269841e-02
R12608 n2_14958_4305 n2_14958_4338 2.095238e-02
R12609 n2_14958_4338 n2_14958_4375 2.349206e-02
R12610 n2_14958_4375 n2_14958_4521 9.269841e-02
R12611 n2_14958_4521 n2_14958_4554 2.095238e-02
R12612 n2_14958_4554 n2_14958_4591 2.349206e-02
R12613 n2_14958_4591 n2_14958_4737 9.269841e-02
R12614 n2_14958_4737 n2_14958_4770 2.095238e-02
R12615 n2_14958_4770 n2_14958_4807 2.349206e-02
R12616 n2_14958_4807 n2_14958_4924 7.428571e-02
R12617 n2_14958_4924 n2_14958_4953 1.841270e-02
R12618 n2_14958_4953 n2_14958_4986 2.095238e-02
R12619 n2_14958_4986 n2_14958_5020 2.158730e-02
R12620 n2_14958_5020 n2_14958_5169 9.460317e-02
R12621 n2_14958_5169 n2_14958_5202 2.095238e-02
R12622 n2_14958_5202 n2_14958_5239 2.349206e-02
R12623 n2_14958_5239 n2_14958_5385 9.269841e-02
R12624 n2_14958_5385 n2_14958_5418 2.095238e-02
R12625 n2_14958_5418 n2_14958_5455 2.349206e-02
R12626 n2_14958_5455 n2_14958_5601 9.269841e-02
R12627 n2_14958_5601 n2_14958_5634 2.095238e-02
R12628 n2_14958_5634 n2_14958_5671 2.349206e-02
R12629 n2_14958_5671 n2_14958_5817 9.269841e-02
R12630 n2_14958_5817 n2_14958_5850 2.095238e-02
R12631 n2_14958_5850 n2_14958_6033 1.161905e-01
R12632 n2_14958_6033 n2_14958_6049 1.015873e-02
R12633 n2_14958_6049 n2_14958_6066 1.079365e-02
R12634 n2_14958_6066 n2_14958_6145 5.015873e-02
R12635 n2_14958_15049 n2_14958_15105 3.555556e-02
R12636 n2_14958_15105 n2_14958_15138 2.095238e-02
R12637 n2_14958_15138 n2_14958_15145 4.444444e-03
R12638 n2_14958_15145 n2_14958_15159 8.888889e-03
R12639 n2_14958_15159 n2_14958_15321 1.028571e-01
R12640 n2_14958_15321 n2_14958_15354 2.095238e-02
R12641 n2_14958_15354 n2_14958_15368 8.888889e-03
R12642 n2_14958_15368 n2_14958_15537 1.073016e-01
R12643 n2_14958_15537 n2_14958_15570 2.095238e-02
R12644 n2_14958_15570 n2_14958_15584 8.888889e-03
R12645 n2_14958_15584 n2_14958_15753 1.073016e-01
R12646 n2_14958_15753 n2_14958_15786 2.095238e-02
R12647 n2_14958_15786 n2_14958_15800 8.888889e-03
R12648 n2_14958_15800 n2_14958_15969 1.073016e-01
R12649 n2_14958_15969 n2_14958_16002 2.095238e-02
R12650 n2_14958_16002 n2_14958_16174 1.092063e-01
R12651 n2_14958_16174 n2_14958_16185 6.984127e-03
R12652 n2_14958_16185 n2_14958_16218 2.095238e-02
R12653 n2_14958_16218 n2_14958_16270 3.301587e-02
R12654 n2_14958_16270 n2_14958_16401 8.317460e-02
R12655 n2_14958_16401 n2_14958_16434 2.095238e-02
R12656 n2_14958_16434 n2_14958_16448 8.888889e-03
R12657 n2_14958_16448 n2_14958_16617 1.073016e-01
R12658 n2_14958_16617 n2_14958_16650 2.095238e-02
R12659 n2_14958_16650 n2_14958_16687 2.349206e-02
R12660 n2_14958_16687 n2_14958_16833 9.269841e-02
R12661 n2_14958_16833 n2_14958_16866 2.095238e-02
R12662 n2_14958_16866 n2_14958_17049 1.161905e-01
R12663 n2_14958_17049 n2_14958_17082 2.095238e-02
R12664 n2_14958_17082 n2_14958_17096 8.888889e-03
R12665 n2_14958_17096 n2_14958_17265 1.073016e-01
R12666 n2_14958_17265 n2_14958_17298 2.095238e-02
R12667 n2_14958_17298 n2_14958_17299 6.349206e-04
R12668 n2_14958_17299 n2_14958_17395 6.095238e-02
R12669 n2_14958_17395 n2_14958_17481 5.460317e-02
R12670 n2_14958_17481 n2_14958_17514 2.095238e-02
R12671 n2_14958_17514 n2_14958_17528 8.888889e-03
R12672 n2_14958_17528 n2_14958_17697 1.073016e-01
R12673 n2_14958_17697 n2_14958_17730 2.095238e-02
R12674 n2_14958_17730 n2_14958_17913 1.161905e-01
R12675 n2_14958_17913 n2_14958_17946 2.095238e-02
R12676 n2_14958_17946 n2_14958_17983 2.349206e-02
R12677 n2_14958_17983 n2_14958_18129 9.269841e-02
R12678 n2_14958_18129 n2_14958_18162 2.095238e-02
R12679 n2_14958_18162 n2_14958_18176 8.888889e-03
R12680 n2_14958_18176 n2_14958_18345 1.073016e-01
R12681 n2_14958_18345 n2_14958_18378 2.095238e-02
R12682 n2_14958_18378 n2_14958_18424 2.920635e-02
R12683 n2_14958_18424 n2_14958_18520 6.095238e-02
R12684 n2_14958_18520 n2_14958_18561 2.603175e-02
R12685 n2_14958_18561 n2_14958_18594 2.095238e-02
R12686 n2_14958_18594 n2_14958_18608 8.888889e-03
R12687 n2_14958_18608 n2_14958_18777 1.073016e-01
R12688 n2_14958_18777 n2_14958_18810 2.095238e-02
R12689 n2_14958_18810 n2_14958_18993 1.161905e-01
R12690 n2_14958_18993 n2_14958_19026 2.095238e-02
R12691 n2_14958_19026 n2_14958_19209 1.161905e-01
R12692 n2_14958_19209 n2_14958_19242 2.095238e-02
R12693 n2_14958_19242 n2_14958_19256 8.888889e-03
R12694 n2_14958_19256 n2_14958_19263 4.444444e-03
R12695 n2_14958_19263 n2_14958_19425 1.028571e-01
R12696 n2_14958_19425 n2_14958_19458 2.095238e-02
R12697 n2_14958_19458 n2_14958_19549 5.777778e-02
R12698 n2_14958_19549 n2_14958_19641 5.841270e-02
R12699 n2_14958_19641 n2_14958_19645 2.539683e-03
R12700 n2_14958_19645 n2_14958_19674 1.841270e-02
R12701 n2_14958_19674 n2_14958_19857 1.161905e-01
R12702 n2_14958_19857 n2_14958_19890 2.095238e-02
R12703 n2_14958_19890 n2_14958_20073 1.161905e-01
R12704 n2_14958_20073 n2_14958_20106 2.095238e-02
R12705 n2_14958_20106 n2_14958_20289 1.161905e-01
R12706 n2_14958_20289 n2_14958_20322 2.095238e-02
R12707 n2_14958_20322 n2_14958_20505 1.161905e-01
R12708 n2_14958_20505 n2_14958_20538 2.095238e-02
R12709 n2_14958_20538 n2_14958_20674 8.634921e-02
R12710 n2_14958_20674 n2_14958_20721 2.984127e-02
R12711 n2_14958_20721 n2_14958_20754 2.095238e-02
R12712 n2_14958_20754 n2_14958_20770 1.015873e-02
R12713 n2_14958_20770 n2_14958_20937 1.060317e-01
R12714 n2_14958_20937 n2_14958_20970 2.095238e-02
R12715 n2_15054_201 n2_15054_234 2.095238e-02
R12716 n2_15054_234 n2_15054_417 1.161905e-01
R12717 n2_15054_417 n2_15054_424 4.444444e-03
R12718 n2_15054_424 n2_15054_450 1.650794e-02
R12719 n2_15054_450 n2_15054_520 4.444444e-02
R12720 n2_15054_520 n2_15054_633 7.174603e-02
R12721 n2_15054_633 n2_15054_666 2.095238e-02
R12722 n2_15054_666 n2_15054_849 1.161905e-01
R12723 n2_15054_849 n2_15054_882 2.095238e-02
R12724 n2_15054_882 n2_15054_1065 1.161905e-01
R12725 n2_15054_1065 n2_15054_1098 2.095238e-02
R12726 n2_15054_1098 n2_15054_1281 1.161905e-01
R12727 n2_15054_1281 n2_15054_1314 2.095238e-02
R12728 n2_15054_1314 n2_15054_1497 1.161905e-01
R12729 n2_15054_1497 n2_15054_1530 2.095238e-02
R12730 n2_15054_1530 n2_15054_1549 1.206349e-02
R12731 n2_15054_1549 n2_15054_1645 6.095238e-02
R12732 n2_15054_1645 n2_15054_1713 4.317460e-02
R12733 n2_15054_1713 n2_15054_1746 2.095238e-02
R12734 n2_15054_1746 n2_15054_1783 2.349206e-02
R12735 n2_15054_1783 n2_15054_1929 9.269841e-02
R12736 n2_15054_1929 n2_15054_1962 2.095238e-02
R12737 n2_15054_1962 n2_15054_2145 1.161905e-01
R12738 n2_15054_2145 n2_15054_2178 2.095238e-02
R12739 n2_15054_2178 n2_15054_2361 1.161905e-01
R12740 n2_15054_2361 n2_15054_2394 2.095238e-02
R12741 n2_15054_2394 n2_15054_2431 2.349206e-02
R12742 n2_15054_2431 n2_15054_2577 9.269841e-02
R12743 n2_15054_2577 n2_15054_2610 2.095238e-02
R12744 n2_15054_2610 n2_15054_2674 4.063492e-02
R12745 n2_15054_2674 n2_15054_2770 6.095238e-02
R12746 n2_15054_2770 n2_15054_2793 1.460317e-02
R12747 n2_15054_2793 n2_15054_2826 2.095238e-02
R12748 n2_15054_2826 n2_15054_2863 2.349206e-02
R12749 n2_15054_2863 n2_15054_3009 9.269841e-02
R12750 n2_15054_3009 n2_15054_3042 2.095238e-02
R12751 n2_15054_3042 n2_15054_3225 1.161905e-01
R12752 n2_15054_3225 n2_15054_3258 2.095238e-02
R12753 n2_15054_3258 n2_15054_3295 2.349206e-02
R12754 n2_15054_3295 n2_15054_3441 9.269841e-02
R12755 n2_15054_3441 n2_15054_3474 2.095238e-02
R12756 n2_15054_3474 n2_15054_3511 2.349206e-02
R12757 n2_15054_3511 n2_15054_3657 9.269841e-02
R12758 n2_15054_3657 n2_15054_3690 2.095238e-02
R12759 n2_15054_3690 n2_15054_3799 6.920635e-02
R12760 n2_15054_3799 n2_15054_3873 4.698413e-02
R12761 n2_15054_3873 n2_15054_3895 1.396825e-02
R12762 n2_15054_3895 n2_15054_3906 6.984127e-03
R12763 n2_15054_3906 n2_15054_3943 2.349206e-02
R12764 n2_15054_3943 n2_15054_4089 9.269841e-02
R12765 n2_15054_4089 n2_15054_4122 2.095238e-02
R12766 n2_15054_4122 n2_15054_4159 2.349206e-02
R12767 n2_15054_4159 n2_15054_4305 9.269841e-02
R12768 n2_15054_4305 n2_15054_4338 2.095238e-02
R12769 n2_15054_4338 n2_15054_4375 2.349206e-02
R12770 n2_15054_4375 n2_15054_4521 9.269841e-02
R12771 n2_15054_4521 n2_15054_4554 2.095238e-02
R12772 n2_15054_4554 n2_15054_4591 2.349206e-02
R12773 n2_15054_4591 n2_15054_4737 9.269841e-02
R12774 n2_15054_4737 n2_15054_4770 2.095238e-02
R12775 n2_15054_4770 n2_15054_4807 2.349206e-02
R12776 n2_15054_4807 n2_15054_4924 7.428571e-02
R12777 n2_15054_4924 n2_15054_4953 1.841270e-02
R12778 n2_15054_4953 n2_15054_4986 2.095238e-02
R12779 n2_15054_4986 n2_15054_5020 2.158730e-02
R12780 n2_15054_5020 n2_15054_5169 9.460317e-02
R12781 n2_15054_5169 n2_15054_5202 2.095238e-02
R12782 n2_15054_5202 n2_15054_5239 2.349206e-02
R12783 n2_15054_5239 n2_15054_5385 9.269841e-02
R12784 n2_15054_5385 n2_15054_5418 2.095238e-02
R12785 n2_15054_5418 n2_15054_5455 2.349206e-02
R12786 n2_15054_5455 n2_15054_5601 9.269841e-02
R12787 n2_15054_5601 n2_15054_5634 2.095238e-02
R12788 n2_15054_5634 n2_15054_5671 2.349206e-02
R12789 n2_15054_5671 n2_15054_5817 9.269841e-02
R12790 n2_15054_5817 n2_15054_5850 2.095238e-02
R12791 n2_15054_5850 n2_15054_6033 1.161905e-01
R12792 n2_15054_6033 n2_15054_6049 1.015873e-02
R12793 n2_15054_6049 n2_15054_6066 1.079365e-02
R12794 n2_15054_6066 n2_15054_6145 5.015873e-02
R12795 n2_15054_6145 n2_15054_6249 6.603175e-02
R12796 n2_15054_6249 n2_15054_6282 2.095238e-02
R12797 n2_15054_6282 n2_15054_6319 2.349206e-02
R12798 n2_15054_6319 n2_15054_6465 9.269841e-02
R12799 n2_15054_6465 n2_15054_6498 2.095238e-02
R12800 n2_15054_6498 n2_15054_6535 2.349206e-02
R12801 n2_15054_6535 n2_15054_6681 9.269841e-02
R12802 n2_15054_6681 n2_15054_6714 2.095238e-02
R12803 n2_15054_6714 n2_15054_6897 1.161905e-01
R12804 n2_15054_6897 n2_15054_6930 2.095238e-02
R12805 n2_15054_6930 n2_15054_7113 1.161905e-01
R12806 n2_15054_7329 n2_15054_7362 2.095238e-02
R12807 n2_15054_7362 n2_15054_7545 1.161905e-01
R12808 n2_15054_7545 n2_15054_7578 2.095238e-02
R12809 n2_15054_7578 n2_15054_7761 1.161905e-01
R12810 n2_15054_7761 n2_15054_7794 2.095238e-02
R12811 n2_15054_7794 n2_15054_7831 2.349206e-02
R12812 n2_15054_7831 n2_15054_7977 9.269841e-02
R12813 n2_15054_7977 n2_15054_8010 2.095238e-02
R12814 n2_15054_8010 n2_15054_8193 1.161905e-01
R12815 n2_15054_8193 n2_15054_8226 2.095238e-02
R12816 n2_15054_8226 n2_15054_8299 4.634921e-02
R12817 n2_15054_8299 n2_15054_8395 6.095238e-02
R12818 n2_15054_8395 n2_15054_8409 8.888889e-03
R12819 n2_15054_8409 n2_15054_8442 2.095238e-02
R12820 n2_15054_8442 n2_15054_8625 1.161905e-01
R12821 n2_15054_8625 n2_15054_8658 2.095238e-02
R12822 n2_15054_8658 n2_15054_8841 1.161905e-01
R12823 n2_15054_8841 n2_15054_8874 2.095238e-02
R12824 n2_15054_8874 n2_15054_8911 2.349206e-02
R12825 n2_15054_8911 n2_15054_9057 9.269841e-02
R12826 n2_15054_9057 n2_15054_9090 2.095238e-02
R12827 n2_15054_9090 n2_15054_9273 1.161905e-01
R12828 n2_15054_9273 n2_15054_9306 2.095238e-02
R12829 n2_15054_9705 n2_15054_9738 2.095238e-02
R12830 n2_15054_9738 n2_15054_9921 1.161905e-01
R12831 n2_15054_9921 n2_15054_9954 2.095238e-02
R12832 n2_15054_9954 n2_15054_9991 2.349206e-02
R12833 n2_15054_9991 n2_15054_10137 9.269841e-02
R12834 n2_15054_10137 n2_15054_10170 2.095238e-02
R12835 n2_15054_10170 n2_15054_10353 1.161905e-01
R12836 n2_15054_10353 n2_15054_10386 2.095238e-02
R12837 n2_15054_10386 n2_15054_10549 1.034921e-01
R12838 n2_15054_10549 n2_15054_10569 1.269841e-02
R12839 n2_15054_10569 n2_15054_10602 2.095238e-02
R12840 n2_15054_10602 n2_15054_10645 2.730159e-02
R12841 n2_15054_10645 n2_15054_10785 8.888889e-02
R12842 n2_15054_10785 n2_15054_10818 2.095238e-02
R12843 n2_15054_10818 n2_15054_11001 1.161905e-01
R12844 n2_15054_11001 n2_15054_11034 2.095238e-02
R12845 n2_15054_11034 n2_15054_11048 8.888889e-03
R12846 n2_15054_11048 n2_15054_11217 1.073016e-01
R12847 n2_15054_11217 n2_15054_11250 2.095238e-02
R12848 n2_15054_11250 n2_15054_11433 1.161905e-01
R12849 n2_15054_11433 n2_15054_11466 2.095238e-02
R12850 n2_15054_11865 n2_15054_11898 2.095238e-02
R12851 n2_15054_11898 n2_15054_12081 1.161905e-01
R12852 n2_15054_12081 n2_15054_12114 2.095238e-02
R12853 n2_15054_12114 n2_15054_12128 8.888889e-03
R12854 n2_15054_12128 n2_15054_12135 4.444444e-03
R12855 n2_15054_12135 n2_15054_12297 1.028571e-01
R12856 n2_15054_12297 n2_15054_12330 2.095238e-02
R12857 n2_15054_12330 n2_15054_12513 1.161905e-01
R12858 n2_15054_12513 n2_15054_12546 2.095238e-02
R12859 n2_15054_12546 n2_15054_12729 1.161905e-01
R12860 n2_15054_12729 n2_15054_12762 2.095238e-02
R12861 n2_15054_12762 n2_15054_12776 8.888889e-03
R12862 n2_15054_12776 n2_15054_12799 1.460317e-02
R12863 n2_15054_12799 n2_15054_12895 6.095238e-02
R12864 n2_15054_12895 n2_15054_12945 3.174603e-02
R12865 n2_15054_12945 n2_15054_12978 2.095238e-02
R12866 n2_15054_12978 n2_15054_12992 8.888889e-03
R12867 n2_15054_12992 n2_15054_13161 1.073016e-01
R12868 n2_15054_13161 n2_15054_13194 2.095238e-02
R12869 n2_15054_13194 n2_15054_13377 1.161905e-01
R12870 n2_15054_13377 n2_15054_13410 2.095238e-02
R12871 n2_15054_13410 n2_15054_13423 8.253968e-03
R12872 n2_15054_13423 n2_15054_13593 1.079365e-01
R12873 n2_15054_13593 n2_15054_13626 2.095238e-02
R12874 n2_15054_13626 n2_15054_13809 1.161905e-01
R12875 n2_15054_13809 n2_15054_13842 2.095238e-02
R12876 n2_15054_14241 n2_15054_14274 2.095238e-02
R12877 n2_15054_14274 n2_15054_14457 1.161905e-01
R12878 n2_15054_14457 n2_15054_14490 2.095238e-02
R12879 n2_15054_14490 n2_15054_14511 1.333333e-02
R12880 n2_15054_14511 n2_15054_14673 1.028571e-01
R12881 n2_15054_14673 n2_15054_14706 2.095238e-02
R12882 n2_15054_14706 n2_15054_14889 1.161905e-01
R12883 n2_15054_14889 n2_15054_14922 2.095238e-02
R12884 n2_15054_14922 n2_15054_14943 1.333333e-02
R12885 n2_15054_14943 n2_15054_15049 6.730159e-02
R12886 n2_15054_15049 n2_15054_15105 3.555556e-02
R12887 n2_15054_15105 n2_15054_15138 2.095238e-02
R12888 n2_15054_15138 n2_15054_15145 4.444444e-03
R12889 n2_15054_15145 n2_15054_15159 8.888889e-03
R12890 n2_15054_15159 n2_15054_15321 1.028571e-01
R12891 n2_15054_15321 n2_15054_15354 2.095238e-02
R12892 n2_15054_15354 n2_15054_15368 8.888889e-03
R12893 n2_15054_15368 n2_15054_15537 1.073016e-01
R12894 n2_15054_15537 n2_15054_15570 2.095238e-02
R12895 n2_15054_15570 n2_15054_15584 8.888889e-03
R12896 n2_15054_15584 n2_15054_15753 1.073016e-01
R12897 n2_15054_15753 n2_15054_15786 2.095238e-02
R12898 n2_15054_15786 n2_15054_15800 8.888889e-03
R12899 n2_15054_15800 n2_15054_15969 1.073016e-01
R12900 n2_15054_15969 n2_15054_16002 2.095238e-02
R12901 n2_15054_16002 n2_15054_16174 1.092063e-01
R12902 n2_15054_16174 n2_15054_16185 6.984127e-03
R12903 n2_15054_16185 n2_15054_16218 2.095238e-02
R12904 n2_15054_16218 n2_15054_16270 3.301587e-02
R12905 n2_15054_16270 n2_15054_16401 8.317460e-02
R12906 n2_15054_16401 n2_15054_16434 2.095238e-02
R12907 n2_15054_16434 n2_15054_16448 8.888889e-03
R12908 n2_15054_16448 n2_15054_16617 1.073016e-01
R12909 n2_15054_16617 n2_15054_16650 2.095238e-02
R12910 n2_15054_16650 n2_15054_16687 2.349206e-02
R12911 n2_15054_16687 n2_15054_16833 9.269841e-02
R12912 n2_15054_16833 n2_15054_16866 2.095238e-02
R12913 n2_15054_16866 n2_15054_17049 1.161905e-01
R12914 n2_15054_17049 n2_15054_17082 2.095238e-02
R12915 n2_15054_17082 n2_15054_17096 8.888889e-03
R12916 n2_15054_17096 n2_15054_17265 1.073016e-01
R12917 n2_15054_17265 n2_15054_17298 2.095238e-02
R12918 n2_15054_17298 n2_15054_17299 6.349206e-04
R12919 n2_15054_17299 n2_15054_17395 6.095238e-02
R12920 n2_15054_17395 n2_15054_17481 5.460317e-02
R12921 n2_15054_17481 n2_15054_17514 2.095238e-02
R12922 n2_15054_17514 n2_15054_17528 8.888889e-03
R12923 n2_15054_17528 n2_15054_17697 1.073016e-01
R12924 n2_15054_17697 n2_15054_17730 2.095238e-02
R12925 n2_15054_17730 n2_15054_17913 1.161905e-01
R12926 n2_15054_17913 n2_15054_17946 2.095238e-02
R12927 n2_15054_17946 n2_15054_17983 2.349206e-02
R12928 n2_15054_17983 n2_15054_18129 9.269841e-02
R12929 n2_15054_18129 n2_15054_18162 2.095238e-02
R12930 n2_15054_18162 n2_15054_18176 8.888889e-03
R12931 n2_15054_18176 n2_15054_18345 1.073016e-01
R12932 n2_15054_18345 n2_15054_18378 2.095238e-02
R12933 n2_15054_18378 n2_15054_18424 2.920635e-02
R12934 n2_15054_18424 n2_15054_18520 6.095238e-02
R12935 n2_15054_18520 n2_15054_18561 2.603175e-02
R12936 n2_15054_18561 n2_15054_18594 2.095238e-02
R12937 n2_15054_18594 n2_15054_18608 8.888889e-03
R12938 n2_15054_18608 n2_15054_18777 1.073016e-01
R12939 n2_15054_18777 n2_15054_18810 2.095238e-02
R12940 n2_15054_18810 n2_15054_18993 1.161905e-01
R12941 n2_15054_18993 n2_15054_19026 2.095238e-02
R12942 n2_15054_19026 n2_15054_19209 1.161905e-01
R12943 n2_15054_19209 n2_15054_19242 2.095238e-02
R12944 n2_15054_19242 n2_15054_19256 8.888889e-03
R12945 n2_15054_19256 n2_15054_19263 4.444444e-03
R12946 n2_15054_19263 n2_15054_19425 1.028571e-01
R12947 n2_15054_19425 n2_15054_19458 2.095238e-02
R12948 n2_15054_19458 n2_15054_19549 5.777778e-02
R12949 n2_15054_19549 n2_15054_19641 5.841270e-02
R12950 n2_15054_19641 n2_15054_19645 2.539683e-03
R12951 n2_15054_19645 n2_15054_19674 1.841270e-02
R12952 n2_15054_19674 n2_15054_19857 1.161905e-01
R12953 n2_15054_19857 n2_15054_19890 2.095238e-02
R12954 n2_15054_19890 n2_15054_20073 1.161905e-01
R12955 n2_15054_20073 n2_15054_20106 2.095238e-02
R12956 n2_15054_20106 n2_15054_20289 1.161905e-01
R12957 n2_15054_20289 n2_15054_20322 2.095238e-02
R12958 n2_15054_20322 n2_15054_20505 1.161905e-01
R12959 n2_15054_20505 n2_15054_20538 2.095238e-02
R12960 n2_15054_20538 n2_15054_20674 8.634921e-02
R12961 n2_15054_20674 n2_15054_20721 2.984127e-02
R12962 n2_15054_20721 n2_15054_20754 2.095238e-02
R12963 n2_15054_20754 n2_15054_20770 1.015873e-02
R12964 n2_15054_20770 n2_15054_20937 1.060317e-01
R12965 n2_15054_20937 n2_15054_20970 2.095238e-02
R12966 n2_15146_201 n2_15146_234 2.095238e-02
R12967 n2_15146_234 n2_15146_417 1.161905e-01
R12968 n2_15146_417 n2_15146_424 4.444444e-03
R12969 n2_15146_424 n2_15146_450 1.650794e-02
R12970 n2_15146_520 n2_15146_633 7.174603e-02
R12971 n2_15146_633 n2_15146_666 2.095238e-02
R12972 n2_15146_666 n2_15146_849 1.161905e-01
R12973 n2_15146_849 n2_15146_882 2.095238e-02
R12974 n2_15146_882 n2_15146_1065 1.161905e-01
R12975 n2_15146_1065 n2_15146_1098 2.095238e-02
R12976 n2_15146_1098 n2_15146_1281 1.161905e-01
R12977 n2_15146_1281 n2_15146_1314 2.095238e-02
R12978 n2_15146_1314 n2_15146_1497 1.161905e-01
R12979 n2_15146_1497 n2_15146_1530 2.095238e-02
R12980 n2_15146_1530 n2_15146_1549 1.206349e-02
R12981 n2_15146_1645 n2_15146_1713 4.317460e-02
R12982 n2_15146_1713 n2_15146_1746 2.095238e-02
R12983 n2_15146_1746 n2_15146_1783 2.349206e-02
R12984 n2_15146_1783 n2_15146_1929 9.269841e-02
R12985 n2_15146_1929 n2_15146_1962 2.095238e-02
R12986 n2_15146_1962 n2_15146_2145 1.161905e-01
R12987 n2_15146_2145 n2_15146_2178 2.095238e-02
R12988 n2_15146_2178 n2_15146_2361 1.161905e-01
R12989 n2_15146_2361 n2_15146_2394 2.095238e-02
R12990 n2_15146_2394 n2_15146_2431 2.349206e-02
R12991 n2_15146_2431 n2_15146_2577 9.269841e-02
R12992 n2_15146_2577 n2_15146_2610 2.095238e-02
R12993 n2_15146_2610 n2_15146_2674 4.063492e-02
R12994 n2_15146_2770 n2_15146_2793 1.460317e-02
R12995 n2_15146_2793 n2_15146_2826 2.095238e-02
R12996 n2_15146_2826 n2_15146_2863 2.349206e-02
R12997 n2_15146_2863 n2_15146_3009 9.269841e-02
R12998 n2_15146_3009 n2_15146_3042 2.095238e-02
R12999 n2_15146_3042 n2_15146_3225 1.161905e-01
R13000 n2_15146_3225 n2_15146_3258 2.095238e-02
R13001 n2_15146_3258 n2_15146_3295 2.349206e-02
R13002 n2_15146_3295 n2_15146_3441 9.269841e-02
R13003 n2_15146_3441 n2_15146_3474 2.095238e-02
R13004 n2_15146_3474 n2_15146_3511 2.349206e-02
R13005 n2_15146_3511 n2_15146_3657 9.269841e-02
R13006 n2_15146_3657 n2_15146_3690 2.095238e-02
R13007 n2_15146_3690 n2_15146_3799 6.920635e-02
R13008 n2_15146_3873 n2_15146_3895 1.396825e-02
R13009 n2_15146_3895 n2_15146_3906 6.984127e-03
R13010 n2_15146_3906 n2_15146_3943 2.349206e-02
R13011 n2_15146_3943 n2_15146_4089 9.269841e-02
R13012 n2_15146_4089 n2_15146_4122 2.095238e-02
R13013 n2_15146_4122 n2_15146_4159 2.349206e-02
R13014 n2_15146_4159 n2_15146_4305 9.269841e-02
R13015 n2_15146_4305 n2_15146_4338 2.095238e-02
R13016 n2_15146_4338 n2_15146_4375 2.349206e-02
R13017 n2_15146_4375 n2_15146_4521 9.269841e-02
R13018 n2_15146_4521 n2_15146_4554 2.095238e-02
R13019 n2_15146_4554 n2_15146_4591 2.349206e-02
R13020 n2_15146_4591 n2_15146_4737 9.269841e-02
R13021 n2_15146_4737 n2_15146_4770 2.095238e-02
R13022 n2_15146_4770 n2_15146_4807 2.349206e-02
R13023 n2_15146_4807 n2_15146_4924 7.428571e-02
R13024 n2_15146_4924 n2_15146_4953 1.841270e-02
R13025 n2_15146_5020 n2_15146_5169 9.460317e-02
R13026 n2_15146_5169 n2_15146_5202 2.095238e-02
R13027 n2_15146_5202 n2_15146_5239 2.349206e-02
R13028 n2_15146_5239 n2_15146_5385 9.269841e-02
R13029 n2_15146_5385 n2_15146_5418 2.095238e-02
R13030 n2_15146_5418 n2_15146_5455 2.349206e-02
R13031 n2_15146_5455 n2_15146_5601 9.269841e-02
R13032 n2_15146_5601 n2_15146_5634 2.095238e-02
R13033 n2_15146_5634 n2_15146_5671 2.349206e-02
R13034 n2_15146_5671 n2_15146_5817 9.269841e-02
R13035 n2_15146_5817 n2_15146_5850 2.095238e-02
R13036 n2_15146_5850 n2_15146_6033 1.161905e-01
R13037 n2_15146_6033 n2_15146_6049 1.015873e-02
R13038 n2_15146_6049 n2_15146_6066 1.079365e-02
R13039 n2_15146_15138 n2_15146_15145 4.444444e-03
R13040 n2_15146_15145 n2_15146_15159 8.888889e-03
R13041 n2_15146_15159 n2_15146_15321 1.028571e-01
R13042 n2_15146_15321 n2_15146_15354 2.095238e-02
R13043 n2_15146_15354 n2_15146_15368 8.888889e-03
R13044 n2_15146_15368 n2_15146_15537 1.073016e-01
R13045 n2_15146_15537 n2_15146_15570 2.095238e-02
R13046 n2_15146_15570 n2_15146_15584 8.888889e-03
R13047 n2_15146_15584 n2_15146_15753 1.073016e-01
R13048 n2_15146_15753 n2_15146_15786 2.095238e-02
R13049 n2_15146_15786 n2_15146_15800 8.888889e-03
R13050 n2_15146_15800 n2_15146_15969 1.073016e-01
R13051 n2_15146_15969 n2_15146_16002 2.095238e-02
R13052 n2_15146_16002 n2_15146_16174 1.092063e-01
R13053 n2_15146_16174 n2_15146_16185 6.984127e-03
R13054 n2_15146_16270 n2_15146_16401 8.317460e-02
R13055 n2_15146_16401 n2_15146_16434 2.095238e-02
R13056 n2_15146_16434 n2_15146_16448 8.888889e-03
R13057 n2_15146_16448 n2_15146_16617 1.073016e-01
R13058 n2_15146_16617 n2_15146_16650 2.095238e-02
R13059 n2_15146_16650 n2_15146_16687 2.349206e-02
R13060 n2_15146_16687 n2_15146_16833 9.269841e-02
R13061 n2_15146_16833 n2_15146_16866 2.095238e-02
R13062 n2_15146_16866 n2_15146_17049 1.161905e-01
R13063 n2_15146_17049 n2_15146_17082 2.095238e-02
R13064 n2_15146_17082 n2_15146_17096 8.888889e-03
R13065 n2_15146_17096 n2_15146_17265 1.073016e-01
R13066 n2_15146_17265 n2_15146_17298 2.095238e-02
R13067 n2_15146_17298 n2_15146_17299 6.349206e-04
R13068 n2_15146_17395 n2_15146_17481 5.460317e-02
R13069 n2_15146_17481 n2_15146_17514 2.095238e-02
R13070 n2_15146_17514 n2_15146_17528 8.888889e-03
R13071 n2_15146_17528 n2_15146_17697 1.073016e-01
R13072 n2_15146_17697 n2_15146_17730 2.095238e-02
R13073 n2_15146_17730 n2_15146_17913 1.161905e-01
R13074 n2_15146_17913 n2_15146_17946 2.095238e-02
R13075 n2_15146_17946 n2_15146_17983 2.349206e-02
R13076 n2_15146_17983 n2_15146_18129 9.269841e-02
R13077 n2_15146_18129 n2_15146_18162 2.095238e-02
R13078 n2_15146_18162 n2_15146_18176 8.888889e-03
R13079 n2_15146_18176 n2_15146_18345 1.073016e-01
R13080 n2_15146_18345 n2_15146_18378 2.095238e-02
R13081 n2_15146_18378 n2_15146_18424 2.920635e-02
R13082 n2_15146_18520 n2_15146_18561 2.603175e-02
R13083 n2_15146_18561 n2_15146_18594 2.095238e-02
R13084 n2_15146_18594 n2_15146_18608 8.888889e-03
R13085 n2_15146_18608 n2_15146_18777 1.073016e-01
R13086 n2_15146_18777 n2_15146_18810 2.095238e-02
R13087 n2_15146_18810 n2_15146_18993 1.161905e-01
R13088 n2_15146_18993 n2_15146_19026 2.095238e-02
R13089 n2_15146_19026 n2_15146_19209 1.161905e-01
R13090 n2_15146_19209 n2_15146_19242 2.095238e-02
R13091 n2_15146_19242 n2_15146_19256 8.888889e-03
R13092 n2_15146_19256 n2_15146_19263 4.444444e-03
R13093 n2_15146_19263 n2_15146_19425 1.028571e-01
R13094 n2_15146_19425 n2_15146_19458 2.095238e-02
R13095 n2_15146_19458 n2_15146_19549 5.777778e-02
R13096 n2_15146_19641 n2_15146_19645 2.539683e-03
R13097 n2_15146_19645 n2_15146_19674 1.841270e-02
R13098 n2_15146_19674 n2_15146_19857 1.161905e-01
R13099 n2_15146_19857 n2_15146_19890 2.095238e-02
R13100 n2_15146_19890 n2_15146_20073 1.161905e-01
R13101 n2_15146_20073 n2_15146_20106 2.095238e-02
R13102 n2_15146_20106 n2_15146_20289 1.161905e-01
R13103 n2_15146_20289 n2_15146_20322 2.095238e-02
R13104 n2_15146_20322 n2_15146_20505 1.161905e-01
R13105 n2_15146_20505 n2_15146_20538 2.095238e-02
R13106 n2_15146_20538 n2_15146_20674 8.634921e-02
R13107 n2_15146_20754 n2_15146_20770 1.015873e-02
R13108 n2_15146_20770 n2_15146_20937 1.060317e-01
R13109 n2_15146_20937 n2_15146_20970 2.095238e-02
R13110 n2_15991_5023 n2_15991_5169 9.269841e-02
R13111 n2_15991_5169 n2_15991_5202 2.095238e-02
R13112 n2_15991_5202 n2_15991_5239 2.349206e-02
R13113 n2_15991_5239 n2_15991_5385 9.269841e-02
R13114 n2_15991_5385 n2_15991_5418 2.095238e-02
R13115 n2_15991_5418 n2_15991_5455 2.349206e-02
R13116 n2_15991_5455 n2_15991_5601 9.269841e-02
R13117 n2_15991_5601 n2_15991_5634 2.095238e-02
R13118 n2_15991_5634 n2_15991_5817 1.161905e-01
R13119 n2_15991_5817 n2_15991_5850 2.095238e-02
R13120 n2_15991_5850 n2_15991_6033 1.161905e-01
R13121 n2_15991_6033 n2_15991_6049 1.015873e-02
R13122 n2_15991_6049 n2_15991_6066 1.079365e-02
R13123 n2_15991_6145 n2_15991_6249 6.603175e-02
R13124 n2_15991_6249 n2_15991_6282 2.095238e-02
R13125 n2_15991_6282 n2_15991_6319 2.349206e-02
R13126 n2_15991_6319 n2_15991_6465 9.269841e-02
R13127 n2_15991_6465 n2_15991_6498 2.095238e-02
R13128 n2_15991_6498 n2_15991_6681 1.161905e-01
R13129 n2_15991_6681 n2_15991_6714 2.095238e-02
R13130 n2_15991_6714 n2_15991_6897 1.161905e-01
R13131 n2_15991_6897 n2_15991_6930 2.095238e-02
R13132 n2_15991_6930 n2_15991_7113 1.161905e-01
R13133 n2_15991_7113 n2_15991_7146 2.095238e-02
R13134 n2_15991_7146 n2_15991_7329 1.161905e-01
R13135 n2_15991_7329 n2_15991_7362 2.095238e-02
R13136 n2_15991_7362 n2_15991_7545 1.161905e-01
R13137 n2_15991_7545 n2_15991_7578 2.095238e-02
R13138 n2_15991_7578 n2_15991_7761 1.161905e-01
R13139 n2_15991_7761 n2_15991_7794 2.095238e-02
R13140 n2_15991_7794 n2_15991_7831 2.349206e-02
R13141 n2_15991_7831 n2_15991_7977 9.269841e-02
R13142 n2_15991_7977 n2_15991_8010 2.095238e-02
R13143 n2_15991_8010 n2_15991_8193 1.161905e-01
R13144 n2_15991_8193 n2_15991_8226 2.095238e-02
R13145 n2_15991_8226 n2_15991_8299 4.634921e-02
R13146 n2_15991_8395 n2_15991_8409 8.888889e-03
R13147 n2_15991_8409 n2_15991_8442 2.095238e-02
R13148 n2_15991_8442 n2_15991_8625 1.161905e-01
R13149 n2_15991_8625 n2_15991_8658 2.095238e-02
R13150 n2_15991_8658 n2_15991_8841 1.161905e-01
R13151 n2_15991_8841 n2_15991_8874 2.095238e-02
R13152 n2_15991_8874 n2_15991_8911 2.349206e-02
R13153 n2_15991_8911 n2_15991_9057 9.269841e-02
R13154 n2_15991_9057 n2_15991_9090 2.095238e-02
R13155 n2_15991_9090 n2_15991_9273 1.161905e-01
R13156 n2_15991_9273 n2_15991_9306 2.095238e-02
R13157 n2_15991_9306 n2_15991_9489 1.161905e-01
R13158 n2_15991_9489 n2_15991_9522 2.095238e-02
R13159 n2_15991_9522 n2_15991_9705 1.161905e-01
R13160 n2_15991_9705 n2_15991_9738 2.095238e-02
R13161 n2_15991_9738 n2_15991_9921 1.161905e-01
R13162 n2_15991_9921 n2_15991_9954 2.095238e-02
R13163 n2_15991_9954 n2_15991_9991 2.349206e-02
R13164 n2_15991_9991 n2_15991_10137 9.269841e-02
R13165 n2_15991_10137 n2_15991_10170 2.095238e-02
R13166 n2_15991_10170 n2_15991_10353 1.161905e-01
R13167 n2_15991_10353 n2_15991_10386 2.095238e-02
R13168 n2_15991_10386 n2_15991_10549 1.034921e-01
R13169 n2_15991_10549 n2_15991_10569 1.269841e-02
R13170 n2_15991_10645 n2_15991_10785 8.888889e-02
R13171 n2_15991_10785 n2_15991_10818 2.095238e-02
R13172 n2_15991_10818 n2_15991_11001 1.161905e-01
R13173 n2_15991_11001 n2_15991_11034 2.095238e-02
R13174 n2_15991_11034 n2_15991_11048 8.888889e-03
R13175 n2_15991_11048 n2_15991_11217 1.073016e-01
R13176 n2_15991_11217 n2_15991_11250 2.095238e-02
R13177 n2_15991_11250 n2_15991_11433 1.161905e-01
R13178 n2_15991_11433 n2_15991_11466 2.095238e-02
R13179 n2_15991_11466 n2_15991_11649 1.161905e-01
R13180 n2_15991_11649 n2_15991_11682 2.095238e-02
R13181 n2_15991_11682 n2_15991_11865 1.161905e-01
R13182 n2_15991_11865 n2_15991_11898 2.095238e-02
R13183 n2_15991_11898 n2_15991_12081 1.161905e-01
R13184 n2_15991_12081 n2_15991_12114 2.095238e-02
R13185 n2_15991_12114 n2_15991_12128 8.888889e-03
R13186 n2_15991_12128 n2_15991_12135 4.444444e-03
R13187 n2_15991_12135 n2_15991_12297 1.028571e-01
R13188 n2_15991_12297 n2_15991_12330 2.095238e-02
R13189 n2_15991_12330 n2_15991_12513 1.161905e-01
R13190 n2_15991_12513 n2_15991_12546 2.095238e-02
R13191 n2_15991_12546 n2_15991_12729 1.161905e-01
R13192 n2_15991_12729 n2_15991_12762 2.095238e-02
R13193 n2_15991_12762 n2_15991_12776 8.888889e-03
R13194 n2_15991_12776 n2_15991_12799 1.460317e-02
R13195 n2_15991_12895 n2_15991_12945 3.174603e-02
R13196 n2_15991_12945 n2_15991_12978 2.095238e-02
R13197 n2_15991_12978 n2_15991_12992 8.888889e-03
R13198 n2_15991_12992 n2_15991_13161 1.073016e-01
R13199 n2_15991_13161 n2_15991_13194 2.095238e-02
R13200 n2_15991_13194 n2_15991_13377 1.161905e-01
R13201 n2_15991_13377 n2_15991_13410 2.095238e-02
R13202 n2_15991_13410 n2_15991_13423 8.253968e-03
R13203 n2_15991_13423 n2_15991_13593 1.079365e-01
R13204 n2_15991_13593 n2_15991_13626 2.095238e-02
R13205 n2_15991_13626 n2_15991_13647 1.333333e-02
R13206 n2_15991_13647 n2_15991_13809 1.028571e-01
R13207 n2_15991_13809 n2_15991_13842 2.095238e-02
R13208 n2_15991_13842 n2_15991_14025 1.161905e-01
R13209 n2_15991_14025 n2_15991_14058 2.095238e-02
R13210 n2_15991_14058 n2_15991_14241 1.161905e-01
R13211 n2_15991_14241 n2_15991_14274 2.095238e-02
R13212 n2_15991_14274 n2_15991_14457 1.161905e-01
R13213 n2_15991_14457 n2_15991_14490 2.095238e-02
R13214 n2_15991_14490 n2_15991_14511 1.333333e-02
R13215 n2_15991_14511 n2_15991_14673 1.028571e-01
R13216 n2_15991_14673 n2_15991_14706 2.095238e-02
R13217 n2_15991_14706 n2_15991_14889 1.161905e-01
R13218 n2_15991_14889 n2_15991_14922 2.095238e-02
R13219 n2_15991_14922 n2_15991_14943 1.333333e-02
R13220 n2_15991_14943 n2_15991_15049 6.730159e-02
R13221 n2_15991_15138 n2_15991_15145 4.444444e-03
R13222 n2_15991_15145 n2_15991_15159 8.888889e-03
R13223 n2_15991_15159 n2_15991_15321 1.028571e-01
R13224 n2_15991_15321 n2_15991_15354 2.095238e-02
R13225 n2_15991_15354 n2_15991_15537 1.161905e-01
R13226 n2_15991_15537 n2_15991_15570 2.095238e-02
R13227 n2_15991_15570 n2_15991_15584 8.888889e-03
R13228 n2_15991_15584 n2_15991_15753 1.073016e-01
R13229 n2_15991_15753 n2_15991_15786 2.095238e-02
R13230 n2_15991_15786 n2_15991_15969 1.161905e-01
R13231 n2_15991_15969 n2_15991_16002 2.095238e-02
R13232 n2_15991_16002 n2_15991_16185 1.161905e-01
R13233 n2_15991_6049 n2_16130_6049 8.825397e-02
R13234 n2_16130_6049 n2_16179_6049 3.111111e-02
R13235 n2_15991_6145 n2_16130_6145 8.825397e-02
R13236 n2_16130_6145 n2_16179_6145 3.111111e-02
R13237 n2_15991_8299 n2_16130_8299 8.825397e-02
R13238 n2_16130_8299 n2_16179_8299 3.111111e-02
R13239 n2_15991_8395 n2_16130_8395 8.825397e-02
R13240 n2_16130_8395 n2_16179_8395 3.111111e-02
R13241 n2_15991_10549 n2_16130_10549 8.825397e-02
R13242 n2_16130_10549 n2_16179_10549 3.111111e-02
R13243 n2_15991_10645 n2_16130_10645 8.825397e-02
R13244 n2_16130_10645 n2_16179_10645 3.111111e-02
R13245 n2_15991_12799 n2_16130_12799 8.825397e-02
R13246 n2_16130_12799 n2_16179_12799 3.111111e-02
R13247 n2_15991_12895 n2_16130_12895 8.825397e-02
R13248 n2_16130_12895 n2_16179_12895 3.111111e-02
R13249 n2_15991_15049 n2_16130_15049 8.825397e-02
R13250 n2_16130_15049 n2_16179_15049 3.111111e-02
R13251 n2_15991_15145 n2_16130_15145 8.825397e-02
R13252 n2_16130_15145 n2_16179_15145 3.111111e-02
R13253 n2_16179_5169 n2_16179_5202 2.095238e-02
R13254 n2_16179_5202 n2_16179_5239 2.349206e-02
R13255 n2_16179_5239 n2_16179_5385 9.269841e-02
R13256 n2_16179_5385 n2_16179_5418 2.095238e-02
R13257 n2_16179_5418 n2_16179_5455 2.349206e-02
R13258 n2_16179_5455 n2_16179_5601 9.269841e-02
R13259 n2_16179_5601 n2_16179_5634 2.095238e-02
R13260 n2_16179_5634 n2_16179_5817 1.161905e-01
R13261 n2_16179_5817 n2_16179_5850 2.095238e-02
R13262 n2_16179_5850 n2_16179_6033 1.161905e-01
R13263 n2_16179_6033 n2_16179_6049 1.015873e-02
R13264 n2_16179_6049 n2_16179_6066 1.079365e-02
R13265 n2_16179_6066 n2_16179_6145 5.015873e-02
R13266 n2_16179_6145 n2_16179_6249 6.603175e-02
R13267 n2_16179_6249 n2_16179_6282 2.095238e-02
R13268 n2_16179_6282 n2_16179_6319 2.349206e-02
R13269 n2_16179_6319 n2_16179_6465 9.269841e-02
R13270 n2_16179_6465 n2_16179_6498 2.095238e-02
R13271 n2_16179_6498 n2_16179_6681 1.161905e-01
R13272 n2_16179_6681 n2_16179_6714 2.095238e-02
R13273 n2_16179_6714 n2_16179_6897 1.161905e-01
R13274 n2_16179_6897 n2_16179_6930 2.095238e-02
R13275 n2_16179_6930 n2_16179_7113 1.161905e-01
R13276 n2_16179_7329 n2_16179_7362 2.095238e-02
R13277 n2_16179_7362 n2_16179_7545 1.161905e-01
R13278 n2_16179_7545 n2_16179_7578 2.095238e-02
R13279 n2_16179_7578 n2_16179_7761 1.161905e-01
R13280 n2_16179_7761 n2_16179_7794 2.095238e-02
R13281 n2_16179_7794 n2_16179_7831 2.349206e-02
R13282 n2_16179_7831 n2_16179_7977 9.269841e-02
R13283 n2_16179_7977 n2_16179_8010 2.095238e-02
R13284 n2_16179_8010 n2_16179_8193 1.161905e-01
R13285 n2_16179_8193 n2_16179_8226 2.095238e-02
R13286 n2_16179_8226 n2_16179_8299 4.634921e-02
R13287 n2_16179_8299 n2_16179_8395 6.095238e-02
R13288 n2_16179_8395 n2_16179_8409 8.888889e-03
R13289 n2_16179_8409 n2_16179_8442 2.095238e-02
R13290 n2_16179_8442 n2_16179_8625 1.161905e-01
R13291 n2_16179_8625 n2_16179_8658 2.095238e-02
R13292 n2_16179_8658 n2_16179_8841 1.161905e-01
R13293 n2_16179_8841 n2_16179_8874 2.095238e-02
R13294 n2_16179_8874 n2_16179_8911 2.349206e-02
R13295 n2_16179_8911 n2_16179_9057 9.269841e-02
R13296 n2_16179_9057 n2_16179_9090 2.095238e-02
R13297 n2_16179_9090 n2_16179_9273 1.161905e-01
R13298 n2_16179_9273 n2_16179_9306 2.095238e-02
R13299 n2_16179_9705 n2_16179_9738 2.095238e-02
R13300 n2_16179_9738 n2_16179_9921 1.161905e-01
R13301 n2_16179_9921 n2_16179_9954 2.095238e-02
R13302 n2_16179_9954 n2_16179_9991 2.349206e-02
R13303 n2_16179_9991 n2_16179_10137 9.269841e-02
R13304 n2_16179_10137 n2_16179_10170 2.095238e-02
R13305 n2_16179_10170 n2_16179_10353 1.161905e-01
R13306 n2_16179_10353 n2_16179_10386 2.095238e-02
R13307 n2_16179_10386 n2_16179_10549 1.034921e-01
R13308 n2_16179_10549 n2_16179_10569 1.269841e-02
R13309 n2_16179_10569 n2_16179_10602 2.095238e-02
R13310 n2_16179_10602 n2_16179_10645 2.730159e-02
R13311 n2_16179_10645 n2_16179_10785 8.888889e-02
R13312 n2_16179_10785 n2_16179_10818 2.095238e-02
R13313 n2_16179_10818 n2_16179_11001 1.161905e-01
R13314 n2_16179_11001 n2_16179_11034 2.095238e-02
R13315 n2_16179_11034 n2_16179_11048 8.888889e-03
R13316 n2_16179_11048 n2_16179_11217 1.073016e-01
R13317 n2_16179_11217 n2_16179_11250 2.095238e-02
R13318 n2_16179_11250 n2_16179_11433 1.161905e-01
R13319 n2_16179_11433 n2_16179_11466 2.095238e-02
R13320 n2_16179_11865 n2_16179_11898 2.095238e-02
R13321 n2_16179_11898 n2_16179_12081 1.161905e-01
R13322 n2_16179_12081 n2_16179_12114 2.095238e-02
R13323 n2_16179_12114 n2_16179_12128 8.888889e-03
R13324 n2_16179_12128 n2_16179_12135 4.444444e-03
R13325 n2_16179_12135 n2_16179_12297 1.028571e-01
R13326 n2_16179_12297 n2_16179_12330 2.095238e-02
R13327 n2_16179_12330 n2_16179_12513 1.161905e-01
R13328 n2_16179_12513 n2_16179_12546 2.095238e-02
R13329 n2_16179_12546 n2_16179_12729 1.161905e-01
R13330 n2_16179_12729 n2_16179_12762 2.095238e-02
R13331 n2_16179_12762 n2_16179_12776 8.888889e-03
R13332 n2_16179_12776 n2_16179_12799 1.460317e-02
R13333 n2_16179_12799 n2_16179_12895 6.095238e-02
R13334 n2_16179_12895 n2_16179_12945 3.174603e-02
R13335 n2_16179_12945 n2_16179_12978 2.095238e-02
R13336 n2_16179_12978 n2_16179_12992 8.888889e-03
R13337 n2_16179_12992 n2_16179_13161 1.073016e-01
R13338 n2_16179_13161 n2_16179_13194 2.095238e-02
R13339 n2_16179_13194 n2_16179_13377 1.161905e-01
R13340 n2_16179_13377 n2_16179_13410 2.095238e-02
R13341 n2_16179_13410 n2_16179_13423 8.253968e-03
R13342 n2_16179_13423 n2_16179_13593 1.079365e-01
R13343 n2_16179_13593 n2_16179_13626 2.095238e-02
R13344 n2_16179_13626 n2_16179_13647 1.333333e-02
R13345 n2_16179_13647 n2_16179_13809 1.028571e-01
R13346 n2_16179_13809 n2_16179_13842 2.095238e-02
R13347 n2_16179_14241 n2_16179_14274 2.095238e-02
R13348 n2_16179_14274 n2_16179_14457 1.161905e-01
R13349 n2_16179_14457 n2_16179_14490 2.095238e-02
R13350 n2_16179_14490 n2_16179_14511 1.333333e-02
R13351 n2_16179_14511 n2_16179_14673 1.028571e-01
R13352 n2_16179_14673 n2_16179_14706 2.095238e-02
R13353 n2_16179_14706 n2_16179_14889 1.161905e-01
R13354 n2_16179_14889 n2_16179_14922 2.095238e-02
R13355 n2_16179_14922 n2_16179_14943 1.333333e-02
R13356 n2_16179_14943 n2_16179_15049 6.730159e-02
R13357 n2_16179_15049 n2_16179_15105 3.555556e-02
R13358 n2_16179_15105 n2_16179_15138 2.095238e-02
R13359 n2_16179_15138 n2_16179_15145 4.444444e-03
R13360 n2_16179_15145 n2_16179_15159 8.888889e-03
R13361 n2_16179_15159 n2_16179_15321 1.028571e-01
R13362 n2_16179_15321 n2_16179_15354 2.095238e-02
R13363 n2_16179_15354 n2_16179_15537 1.161905e-01
R13364 n2_16179_15537 n2_16179_15570 2.095238e-02
R13365 n2_16179_15570 n2_16179_15584 8.888889e-03
R13366 n2_16179_15584 n2_16179_15753 1.073016e-01
R13367 n2_16179_15753 n2_16179_15786 2.095238e-02
R13368 n2_16179_15786 n2_16179_15969 1.161905e-01
R13369 n2_16179_15969 n2_16179_16002 2.095238e-02
R13370 n2_17116_201 n2_17116_234 2.095238e-02
R13371 n2_17116_234 n2_17116_417 1.161905e-01
R13372 n2_17116_417 n2_17116_424 4.444444e-03
R13373 n2_17116_424 n2_17116_450 1.650794e-02
R13374 n2_17116_520 n2_17116_633 7.174603e-02
R13375 n2_17116_633 n2_17116_666 2.095238e-02
R13376 n2_17116_666 n2_17116_849 1.161905e-01
R13377 n2_17116_849 n2_17116_882 2.095238e-02
R13378 n2_17116_882 n2_17116_1065 1.161905e-01
R13379 n2_17116_1065 n2_17116_1098 2.095238e-02
R13380 n2_17116_1098 n2_17116_1281 1.161905e-01
R13381 n2_17116_1281 n2_17116_1314 2.095238e-02
R13382 n2_17116_1314 n2_17116_1497 1.161905e-01
R13383 n2_17116_1497 n2_17116_1530 2.095238e-02
R13384 n2_17116_1530 n2_17116_1549 1.206349e-02
R13385 n2_17116_1645 n2_17116_1713 4.317460e-02
R13386 n2_17116_1713 n2_17116_1746 2.095238e-02
R13387 n2_17116_1746 n2_17116_1783 2.349206e-02
R13388 n2_17116_1783 n2_17116_1929 9.269841e-02
R13389 n2_17116_1929 n2_17116_1962 2.095238e-02
R13390 n2_17116_1962 n2_17116_2145 1.161905e-01
R13391 n2_17116_2145 n2_17116_2178 2.095238e-02
R13392 n2_17116_2178 n2_17116_2361 1.161905e-01
R13393 n2_17116_2361 n2_17116_2394 2.095238e-02
R13394 n2_17116_2394 n2_17116_2431 2.349206e-02
R13395 n2_17116_2431 n2_17116_2577 9.269841e-02
R13396 n2_17116_2577 n2_17116_2610 2.095238e-02
R13397 n2_17116_2610 n2_17116_2674 4.063492e-02
R13398 n2_17116_2770 n2_17116_2793 1.460317e-02
R13399 n2_17116_2793 n2_17116_2826 2.095238e-02
R13400 n2_17116_2826 n2_17116_2863 2.349206e-02
R13401 n2_17116_2863 n2_17116_3009 9.269841e-02
R13402 n2_17116_3009 n2_17116_3042 2.095238e-02
R13403 n2_17116_3042 n2_17116_3225 1.161905e-01
R13404 n2_17116_3225 n2_17116_3258 2.095238e-02
R13405 n2_17116_3258 n2_17116_3295 2.349206e-02
R13406 n2_17116_3295 n2_17116_3441 9.269841e-02
R13407 n2_17116_3441 n2_17116_3474 2.095238e-02
R13408 n2_17116_3474 n2_17116_3657 1.161905e-01
R13409 n2_17116_3657 n2_17116_3690 2.095238e-02
R13410 n2_17116_3690 n2_17116_3799 6.920635e-02
R13411 n2_17116_3873 n2_17116_3895 1.396825e-02
R13412 n2_17116_3895 n2_17116_3906 6.984127e-03
R13413 n2_17116_3906 n2_17116_4089 1.161905e-01
R13414 n2_17116_4089 n2_17116_4122 2.095238e-02
R13415 n2_17116_4122 n2_17116_4305 1.161905e-01
R13416 n2_17116_4305 n2_17116_4338 2.095238e-02
R13417 n2_17116_4338 n2_17116_4375 2.349206e-02
R13418 n2_17116_4375 n2_17116_4521 9.269841e-02
R13419 n2_17116_4521 n2_17116_4554 2.095238e-02
R13420 n2_17116_4554 n2_17116_4591 2.349206e-02
R13421 n2_17116_4591 n2_17116_4737 9.269841e-02
R13422 n2_17116_4737 n2_17116_4770 2.095238e-02
R13423 n2_17116_4770 n2_17116_4807 2.349206e-02
R13424 n2_17116_4807 n2_17116_4953 9.269841e-02
R13425 n2_17116_4953 n2_17116_4986 2.095238e-02
R13426 n2_17116_4986 n2_17116_5023 2.349206e-02
R13427 n2_17116_5023 n2_17116_5169 9.269841e-02
R13428 n2_17116_5169 n2_17116_5202 2.095238e-02
R13429 n2_17116_5202 n2_17116_5239 2.349206e-02
R13430 n2_17116_5239 n2_17116_5385 9.269841e-02
R13431 n2_17116_5385 n2_17116_5418 2.095238e-02
R13432 n2_17116_5418 n2_17116_5455 2.349206e-02
R13433 n2_17116_5455 n2_17116_5601 9.269841e-02
R13434 n2_17116_5601 n2_17116_5634 2.095238e-02
R13435 n2_17116_5634 n2_17116_5817 1.161905e-01
R13436 n2_17116_5817 n2_17116_5850 2.095238e-02
R13437 n2_17116_5850 n2_17116_6033 1.161905e-01
R13438 n2_17116_6033 n2_17116_6049 1.015873e-02
R13439 n2_17116_6049 n2_17116_6066 1.079365e-02
R13440 n2_17116_6145 n2_17116_6249 6.603175e-02
R13441 n2_17116_6249 n2_17116_6282 2.095238e-02
R13442 n2_17116_6282 n2_17116_6319 2.349206e-02
R13443 n2_17116_6319 n2_17116_6465 9.269841e-02
R13444 n2_17116_6465 n2_17116_6498 2.095238e-02
R13445 n2_17116_6498 n2_17116_6681 1.161905e-01
R13446 n2_17116_6681 n2_17116_6714 2.095238e-02
R13447 n2_17116_6714 n2_17116_6897 1.161905e-01
R13448 n2_17116_6897 n2_17116_6930 2.095238e-02
R13449 n2_17116_6930 n2_17116_7113 1.161905e-01
R13450 n2_17116_7113 n2_17116_7146 2.095238e-02
R13451 n2_17116_7146 n2_17116_7329 1.161905e-01
R13452 n2_17116_7329 n2_17116_7362 2.095238e-02
R13453 n2_17116_7362 n2_17116_7545 1.161905e-01
R13454 n2_17116_7545 n2_17116_7578 2.095238e-02
R13455 n2_17116_7578 n2_17116_7761 1.161905e-01
R13456 n2_17116_7761 n2_17116_7794 2.095238e-02
R13457 n2_17116_7794 n2_17116_7831 2.349206e-02
R13458 n2_17116_7831 n2_17116_7977 9.269841e-02
R13459 n2_17116_7977 n2_17116_8010 2.095238e-02
R13460 n2_17116_8010 n2_17116_8193 1.161905e-01
R13461 n2_17116_8193 n2_17116_8226 2.095238e-02
R13462 n2_17116_8226 n2_17116_8299 4.634921e-02
R13463 n2_17116_8395 n2_17116_8409 8.888889e-03
R13464 n2_17116_8409 n2_17116_8442 2.095238e-02
R13465 n2_17116_8442 n2_17116_8625 1.161905e-01
R13466 n2_17116_8625 n2_17116_8658 2.095238e-02
R13467 n2_17116_8658 n2_17116_8841 1.161905e-01
R13468 n2_17116_8841 n2_17116_8874 2.095238e-02
R13469 n2_17116_8874 n2_17116_8911 2.349206e-02
R13470 n2_17116_8911 n2_17116_9057 9.269841e-02
R13471 n2_17116_9057 n2_17116_9090 2.095238e-02
R13472 n2_17116_9090 n2_17116_9273 1.161905e-01
R13473 n2_17116_9273 n2_17116_9306 2.095238e-02
R13474 n2_17116_9306 n2_17116_9489 1.161905e-01
R13475 n2_17116_9489 n2_17116_9522 2.095238e-02
R13476 n2_17116_9522 n2_17116_9705 1.161905e-01
R13477 n2_17116_9705 n2_17116_9738 2.095238e-02
R13478 n2_17116_9738 n2_17116_9921 1.161905e-01
R13479 n2_17116_9921 n2_17116_9954 2.095238e-02
R13480 n2_17116_9954 n2_17116_9991 2.349206e-02
R13481 n2_17116_9991 n2_17116_10137 9.269841e-02
R13482 n2_17116_10137 n2_17116_10170 2.095238e-02
R13483 n2_17116_10170 n2_17116_10353 1.161905e-01
R13484 n2_17116_10353 n2_17116_10386 2.095238e-02
R13485 n2_17116_10386 n2_17116_10549 1.034921e-01
R13486 n2_17116_10549 n2_17116_10569 1.269841e-02
R13487 n2_17116_10645 n2_17116_10785 8.888889e-02
R13488 n2_17116_10785 n2_17116_10818 2.095238e-02
R13489 n2_17116_10818 n2_17116_11001 1.161905e-01
R13490 n2_17116_11001 n2_17116_11034 2.095238e-02
R13491 n2_17116_11034 n2_17116_11048 8.888889e-03
R13492 n2_17116_11048 n2_17116_11055 4.444444e-03
R13493 n2_17116_11055 n2_17116_11217 1.028571e-01
R13494 n2_17116_11217 n2_17116_11250 2.095238e-02
R13495 n2_17116_11250 n2_17116_11433 1.161905e-01
R13496 n2_17116_11433 n2_17116_11466 2.095238e-02
R13497 n2_17116_11466 n2_17116_11649 1.161905e-01
R13498 n2_17116_11649 n2_17116_11682 2.095238e-02
R13499 n2_17116_11682 n2_17116_11865 1.161905e-01
R13500 n2_17116_11865 n2_17116_11898 2.095238e-02
R13501 n2_17116_11898 n2_17116_12081 1.161905e-01
R13502 n2_17116_12081 n2_17116_12114 2.095238e-02
R13503 n2_17116_12114 n2_17116_12128 8.888889e-03
R13504 n2_17116_12128 n2_17116_12135 4.444444e-03
R13505 n2_17116_12135 n2_17116_12297 1.028571e-01
R13506 n2_17116_12297 n2_17116_12330 2.095238e-02
R13507 n2_17116_12330 n2_17116_12513 1.161905e-01
R13508 n2_17116_12513 n2_17116_12546 2.095238e-02
R13509 n2_17116_12546 n2_17116_12729 1.161905e-01
R13510 n2_17116_12729 n2_17116_12762 2.095238e-02
R13511 n2_17116_12762 n2_17116_12799 2.349206e-02
R13512 n2_17116_12895 n2_17116_12945 3.174603e-02
R13513 n2_17116_12945 n2_17116_12978 2.095238e-02
R13514 n2_17116_12978 n2_17116_13161 1.161905e-01
R13515 n2_17116_13161 n2_17116_13194 2.095238e-02
R13516 n2_17116_13194 n2_17116_13377 1.161905e-01
R13517 n2_17116_13377 n2_17116_13410 2.095238e-02
R13518 n2_17116_13410 n2_17116_13593 1.161905e-01
R13519 n2_17116_13593 n2_17116_13626 2.095238e-02
R13520 n2_17116_13626 n2_17116_13640 8.888889e-03
R13521 n2_17116_13640 n2_17116_13647 4.444444e-03
R13522 n2_17116_13647 n2_17116_13809 1.028571e-01
R13523 n2_17116_13809 n2_17116_13842 2.095238e-02
R13524 n2_17116_13842 n2_17116_14025 1.161905e-01
R13525 n2_17116_14025 n2_17116_14058 2.095238e-02
R13526 n2_17116_14058 n2_17116_14241 1.161905e-01
R13527 n2_17116_14241 n2_17116_14274 2.095238e-02
R13528 n2_17116_14274 n2_17116_14457 1.161905e-01
R13529 n2_17116_14457 n2_17116_14490 2.095238e-02
R13530 n2_17116_14490 n2_17116_14511 1.333333e-02
R13531 n2_17116_14511 n2_17116_14673 1.028571e-01
R13532 n2_17116_14673 n2_17116_14706 2.095238e-02
R13533 n2_17116_14706 n2_17116_14889 1.161905e-01
R13534 n2_17116_14889 n2_17116_14922 2.095238e-02
R13535 n2_17116_14922 n2_17116_14936 8.888889e-03
R13536 n2_17116_14936 n2_17116_14943 4.444444e-03
R13537 n2_17116_14943 n2_17116_15049 6.730159e-02
R13538 n2_17116_15138 n2_17116_15145 4.444444e-03
R13539 n2_17116_15145 n2_17116_15152 4.444444e-03
R13540 n2_17116_15152 n2_17116_15159 4.444444e-03
R13541 n2_17116_15159 n2_17116_15321 1.028571e-01
R13542 n2_17116_15321 n2_17116_15354 2.095238e-02
R13543 n2_17116_15354 n2_17116_15537 1.161905e-01
R13544 n2_17116_15537 n2_17116_15570 2.095238e-02
R13545 n2_17116_15570 n2_17116_15584 8.888889e-03
R13546 n2_17116_15584 n2_17116_15753 1.073016e-01
R13547 n2_17116_15753 n2_17116_15786 2.095238e-02
R13548 n2_17116_15786 n2_17116_15969 1.161905e-01
R13549 n2_17116_15969 n2_17116_16002 2.095238e-02
R13550 n2_17116_16002 n2_17116_16185 1.161905e-01
R13551 n2_17116_16185 n2_17116_16218 2.095238e-02
R13552 n2_17116_16218 n2_17116_16401 1.161905e-01
R13553 n2_17116_16401 n2_17116_16434 2.095238e-02
R13554 n2_17116_16434 n2_17116_16617 1.161905e-01
R13555 n2_17116_16617 n2_17116_16650 2.095238e-02
R13556 n2_17116_16650 n2_17116_16664 8.888889e-03
R13557 n2_17116_16664 n2_17116_16687 1.460317e-02
R13558 n2_17116_16687 n2_17116_16833 9.269841e-02
R13559 n2_17116_16833 n2_17116_16866 2.095238e-02
R13560 n2_17116_16866 n2_17116_17049 1.161905e-01
R13561 n2_17116_17049 n2_17116_17082 2.095238e-02
R13562 n2_17116_17082 n2_17116_17119 2.349206e-02
R13563 n2_17116_17119 n2_17116_17265 9.269841e-02
R13564 n2_17116_17265 n2_17116_17298 2.095238e-02
R13565 n2_17116_17298 n2_17116_17299 6.349206e-04
R13566 n2_17116_17395 n2_17116_17481 5.460317e-02
R13567 n2_17116_17481 n2_17116_17514 2.095238e-02
R13568 n2_17116_17514 n2_17116_17535 1.333333e-02
R13569 n2_17116_17535 n2_17116_17697 1.028571e-01
R13570 n2_17116_17697 n2_17116_17730 2.095238e-02
R13571 n2_17116_17730 n2_17116_17913 1.161905e-01
R13572 n2_17116_17913 n2_17116_17946 2.095238e-02
R13573 n2_17116_17946 n2_17116_18129 1.161905e-01
R13574 n2_17116_18129 n2_17116_18162 2.095238e-02
R13575 n2_17116_18162 n2_17116_18176 8.888889e-03
R13576 n2_17116_18176 n2_17116_18345 1.073016e-01
R13577 n2_17116_18345 n2_17116_18378 2.095238e-02
R13578 n2_17116_18378 n2_17116_18424 2.920635e-02
R13579 n2_17116_18520 n2_17116_18561 2.603175e-02
R13580 n2_17116_18561 n2_17116_18594 2.095238e-02
R13581 n2_17116_18594 n2_17116_18777 1.161905e-01
R13582 n2_17116_18777 n2_17116_18810 2.095238e-02
R13583 n2_17116_18810 n2_17116_18993 1.161905e-01
R13584 n2_17116_18993 n2_17116_19026 2.095238e-02
R13585 n2_17116_19026 n2_17116_19040 8.888889e-03
R13586 n2_17116_19040 n2_17116_19209 1.073016e-01
R13587 n2_17116_19209 n2_17116_19242 2.095238e-02
R13588 n2_17116_19242 n2_17116_19425 1.161905e-01
R13589 n2_17116_19425 n2_17116_19458 2.095238e-02
R13590 n2_17116_19458 n2_17116_19549 5.777778e-02
R13591 n2_17116_19641 n2_17116_19645 2.539683e-03
R13592 n2_17116_19645 n2_17116_19674 1.841270e-02
R13593 n2_17116_19674 n2_17116_19857 1.161905e-01
R13594 n2_17116_19857 n2_17116_19890 2.095238e-02
R13595 n2_17116_19890 n2_17116_20073 1.161905e-01
R13596 n2_17116_20073 n2_17116_20106 2.095238e-02
R13597 n2_17116_20106 n2_17116_20289 1.161905e-01
R13598 n2_17116_20289 n2_17116_20322 2.095238e-02
R13599 n2_17116_20322 n2_17116_20505 1.161905e-01
R13600 n2_17116_20505 n2_17116_20538 2.095238e-02
R13601 n2_17116_20538 n2_17116_20674 8.634921e-02
R13602 n2_17116_20754 n2_17116_20770 1.015873e-02
R13603 n2_17116_20770 n2_17116_20937 1.060317e-01
R13604 n2_17116_20937 n2_17116_20970 2.095238e-02
R13605 n2_17116_3895 n2_17208_3895 5.841270e-02
R13606 n2_17208_3895 n2_17255_3895 2.984127e-02
R13607 n2_17255_3895 n2_17304_3895 3.111111e-02
R13608 n2_17116_6049 n2_17255_6049 8.825397e-02
R13609 n2_17255_6049 n2_17304_6049 3.111111e-02
R13610 n2_17116_6145 n2_17255_6145 8.825397e-02
R13611 n2_17255_6145 n2_17304_6145 3.111111e-02
R13612 n2_17116_8299 n2_17255_8299 8.825397e-02
R13613 n2_17255_8299 n2_17304_8299 3.111111e-02
R13614 n2_17116_8395 n2_17255_8395 8.825397e-02
R13615 n2_17255_8395 n2_17304_8395 3.111111e-02
R13616 n2_17116_10549 n2_17255_10549 8.825397e-02
R13617 n2_17255_10549 n2_17304_10549 3.111111e-02
R13618 n2_17116_10645 n2_17255_10645 8.825397e-02
R13619 n2_17255_10645 n2_17304_10645 3.111111e-02
R13620 n2_17116_12799 n2_17255_12799 8.825397e-02
R13621 n2_17255_12799 n2_17304_12799 3.111111e-02
R13622 n2_17116_12895 n2_17255_12895 8.825397e-02
R13623 n2_17255_12895 n2_17304_12895 3.111111e-02
R13624 n2_17116_15049 n2_17255_15049 8.825397e-02
R13625 n2_17255_15049 n2_17304_15049 3.111111e-02
R13626 n2_17116_15145 n2_17255_15145 8.825397e-02
R13627 n2_17255_15145 n2_17304_15145 3.111111e-02
R13628 n2_17116_17299 n2_17208_17299 5.841270e-02
R13629 n2_17208_17299 n2_17255_17299 2.984127e-02
R13630 n2_17255_17299 n2_17304_17299 3.111111e-02
R13631 n2_17116_424 n2_17208_424 5.841270e-02
R13632 n2_17208_424 n2_17255_424 2.984127e-02
R13633 n2_17255_424 n2_17304_424 3.111111e-02
R13634 n2_17304_424 n2_17396_424 5.841270e-02
R13635 n2_17116_520 n2_17208_520 5.841270e-02
R13636 n2_17208_520 n2_17255_520 2.984127e-02
R13637 n2_17255_520 n2_17304_520 3.111111e-02
R13638 n2_17304_520 n2_17396_520 5.841270e-02
R13639 n2_17116_1549 n2_17208_1549 5.841270e-02
R13640 n2_17208_1549 n2_17255_1549 2.984127e-02
R13641 n2_17255_1549 n2_17304_1549 3.111111e-02
R13642 n2_17304_1549 n2_17396_1549 5.841270e-02
R13643 n2_17116_1645 n2_17208_1645 5.841270e-02
R13644 n2_17208_1645 n2_17255_1645 2.984127e-02
R13645 n2_17255_1645 n2_17304_1645 3.111111e-02
R13646 n2_17304_1645 n2_17396_1645 5.841270e-02
R13647 n2_17116_2674 n2_17208_2674 5.841270e-02
R13648 n2_17208_2674 n2_17255_2674 2.984127e-02
R13649 n2_17255_2674 n2_17304_2674 3.111111e-02
R13650 n2_17304_2674 n2_17396_2674 5.841270e-02
R13651 n2_17116_2770 n2_17208_2770 5.841270e-02
R13652 n2_17208_2770 n2_17255_2770 2.984127e-02
R13653 n2_17255_2770 n2_17304_2770 3.111111e-02
R13654 n2_17304_2770 n2_17396_2770 5.841270e-02
R13655 n2_17116_3799 n2_17208_3799 5.841270e-02
R13656 n2_17208_3799 n2_17255_3799 2.984127e-02
R13657 n2_17255_3799 n2_17304_3799 3.111111e-02
R13658 n2_17304_3799 n2_17396_3799 5.841270e-02
R13659 n2_17116_17395 n2_17208_17395 5.841270e-02
R13660 n2_17208_17395 n2_17255_17395 2.984127e-02
R13661 n2_17255_17395 n2_17304_17395 3.111111e-02
R13662 n2_17304_17395 n2_17396_17395 5.841270e-02
R13663 n2_17116_18424 n2_17208_18424 5.841270e-02
R13664 n2_17208_18424 n2_17255_18424 2.984127e-02
R13665 n2_17255_18424 n2_17304_18424 3.111111e-02
R13666 n2_17304_18424 n2_17396_18424 5.841270e-02
R13667 n2_17116_18520 n2_17208_18520 5.841270e-02
R13668 n2_17208_18520 n2_17255_18520 2.984127e-02
R13669 n2_17255_18520 n2_17304_18520 3.111111e-02
R13670 n2_17304_18520 n2_17396_18520 5.841270e-02
R13671 n2_17116_19549 n2_17208_19549 5.841270e-02
R13672 n2_17208_19549 n2_17255_19549 2.984127e-02
R13673 n2_17255_19549 n2_17304_19549 3.111111e-02
R13674 n2_17304_19549 n2_17396_19549 5.841270e-02
R13675 n2_17116_19645 n2_17208_19645 5.841270e-02
R13676 n2_17208_19645 n2_17255_19645 2.984127e-02
R13677 n2_17255_19645 n2_17304_19645 3.111111e-02
R13678 n2_17304_19645 n2_17396_19645 5.841270e-02
R13679 n2_17116_20674 n2_17208_20674 5.841270e-02
R13680 n2_17208_20674 n2_17255_20674 2.984127e-02
R13681 n2_17255_20674 n2_17304_20674 3.111111e-02
R13682 n2_17304_20674 n2_17396_20674 5.841270e-02
R13683 n2_17116_20770 n2_17208_20770 5.841270e-02
R13684 n2_17208_20770 n2_17255_20770 2.984127e-02
R13685 n2_17255_20770 n2_17304_20770 3.111111e-02
R13686 n2_17304_20770 n2_17396_20770 5.841270e-02
R13687 n2_17208_201 n2_17208_234 2.095238e-02
R13688 n2_17208_234 n2_17208_417 1.161905e-01
R13689 n2_17208_417 n2_17208_424 4.444444e-03
R13690 n2_17208_424 n2_17208_450 1.650794e-02
R13691 n2_17208_450 n2_17208_520 4.444444e-02
R13692 n2_17208_520 n2_17208_633 7.174603e-02
R13693 n2_17208_633 n2_17208_666 2.095238e-02
R13694 n2_17208_666 n2_17208_849 1.161905e-01
R13695 n2_17208_849 n2_17208_882 2.095238e-02
R13696 n2_17208_882 n2_17208_1065 1.161905e-01
R13697 n2_17208_1065 n2_17208_1098 2.095238e-02
R13698 n2_17208_1098 n2_17208_1281 1.161905e-01
R13699 n2_17208_1281 n2_17208_1314 2.095238e-02
R13700 n2_17208_1314 n2_17208_1497 1.161905e-01
R13701 n2_17208_1497 n2_17208_1530 2.095238e-02
R13702 n2_17208_1530 n2_17208_1549 1.206349e-02
R13703 n2_17208_1549 n2_17208_1645 6.095238e-02
R13704 n2_17208_1645 n2_17208_1713 4.317460e-02
R13705 n2_17208_1713 n2_17208_1746 2.095238e-02
R13706 n2_17208_1746 n2_17208_1783 2.349206e-02
R13707 n2_17208_1783 n2_17208_1929 9.269841e-02
R13708 n2_17208_1929 n2_17208_1962 2.095238e-02
R13709 n2_17208_1962 n2_17208_2145 1.161905e-01
R13710 n2_17208_2145 n2_17208_2178 2.095238e-02
R13711 n2_17208_2178 n2_17208_2361 1.161905e-01
R13712 n2_17208_2361 n2_17208_2394 2.095238e-02
R13713 n2_17208_2394 n2_17208_2431 2.349206e-02
R13714 n2_17208_2431 n2_17208_2577 9.269841e-02
R13715 n2_17208_2577 n2_17208_2610 2.095238e-02
R13716 n2_17208_2610 n2_17208_2674 4.063492e-02
R13717 n2_17208_2674 n2_17208_2770 6.095238e-02
R13718 n2_17208_2770 n2_17208_2793 1.460317e-02
R13719 n2_17208_2793 n2_17208_2826 2.095238e-02
R13720 n2_17208_2826 n2_17208_2863 2.349206e-02
R13721 n2_17208_2863 n2_17208_3009 9.269841e-02
R13722 n2_17208_3009 n2_17208_3042 2.095238e-02
R13723 n2_17208_3042 n2_17208_3225 1.161905e-01
R13724 n2_17208_3225 n2_17208_3258 2.095238e-02
R13725 n2_17208_3258 n2_17208_3295 2.349206e-02
R13726 n2_17208_3295 n2_17208_3441 9.269841e-02
R13727 n2_17208_3441 n2_17208_3474 2.095238e-02
R13728 n2_17208_3474 n2_17208_3657 1.161905e-01
R13729 n2_17208_3657 n2_17208_3690 2.095238e-02
R13730 n2_17208_3690 n2_17208_3799 6.920635e-02
R13731 n2_17208_3799 n2_17208_3873 4.698413e-02
R13732 n2_17208_3873 n2_17208_3895 1.396825e-02
R13733 n2_17208_3895 n2_17208_3906 6.984127e-03
R13734 n2_17208_17265 n2_17208_17298 2.095238e-02
R13735 n2_17208_17298 n2_17208_17299 6.349206e-04
R13736 n2_17208_17299 n2_17208_17395 6.095238e-02
R13737 n2_17208_17395 n2_17208_17481 5.460317e-02
R13738 n2_17208_17481 n2_17208_17514 2.095238e-02
R13739 n2_17208_17514 n2_17208_17535 1.333333e-02
R13740 n2_17208_17535 n2_17208_17697 1.028571e-01
R13741 n2_17208_17697 n2_17208_17730 2.095238e-02
R13742 n2_17208_17730 n2_17208_17913 1.161905e-01
R13743 n2_17208_17913 n2_17208_17946 2.095238e-02
R13744 n2_17208_17946 n2_17208_18129 1.161905e-01
R13745 n2_17208_18129 n2_17208_18162 2.095238e-02
R13746 n2_17208_18162 n2_17208_18176 8.888889e-03
R13747 n2_17208_18176 n2_17208_18345 1.073016e-01
R13748 n2_17208_18345 n2_17208_18378 2.095238e-02
R13749 n2_17208_18378 n2_17208_18424 2.920635e-02
R13750 n2_17208_18424 n2_17208_18520 6.095238e-02
R13751 n2_17208_18520 n2_17208_18561 2.603175e-02
R13752 n2_17208_18561 n2_17208_18594 2.095238e-02
R13753 n2_17208_18594 n2_17208_18777 1.161905e-01
R13754 n2_17208_18777 n2_17208_18810 2.095238e-02
R13755 n2_17208_18810 n2_17208_18993 1.161905e-01
R13756 n2_17208_18993 n2_17208_19026 2.095238e-02
R13757 n2_17208_19026 n2_17208_19040 8.888889e-03
R13758 n2_17208_19040 n2_17208_19209 1.073016e-01
R13759 n2_17208_19209 n2_17208_19242 2.095238e-02
R13760 n2_17208_19242 n2_17208_19425 1.161905e-01
R13761 n2_17208_19425 n2_17208_19458 2.095238e-02
R13762 n2_17208_19458 n2_17208_19549 5.777778e-02
R13763 n2_17208_19549 n2_17208_19641 5.841270e-02
R13764 n2_17208_19641 n2_17208_19645 2.539683e-03
R13765 n2_17208_19645 n2_17208_19674 1.841270e-02
R13766 n2_17208_19674 n2_17208_19857 1.161905e-01
R13767 n2_17208_19857 n2_17208_19890 2.095238e-02
R13768 n2_17208_19890 n2_17208_20073 1.161905e-01
R13769 n2_17208_20073 n2_17208_20106 2.095238e-02
R13770 n2_17208_20106 n2_17208_20289 1.161905e-01
R13771 n2_17208_20289 n2_17208_20322 2.095238e-02
R13772 n2_17208_20322 n2_17208_20505 1.161905e-01
R13773 n2_17208_20505 n2_17208_20538 2.095238e-02
R13774 n2_17208_20538 n2_17208_20674 8.634921e-02
R13775 n2_17208_20674 n2_17208_20721 2.984127e-02
R13776 n2_17208_20721 n2_17208_20754 2.095238e-02
R13777 n2_17208_20754 n2_17208_20770 1.015873e-02
R13778 n2_17208_20770 n2_17208_20937 1.060317e-01
R13779 n2_17208_20937 n2_17208_20970 2.095238e-02
R13780 n2_17304_201 n2_17304_234 2.095238e-02
R13781 n2_17304_234 n2_17304_417 1.161905e-01
R13782 n2_17304_417 n2_17304_424 4.444444e-03
R13783 n2_17304_424 n2_17304_450 1.650794e-02
R13784 n2_17304_450 n2_17304_520 4.444444e-02
R13785 n2_17304_520 n2_17304_633 7.174603e-02
R13786 n2_17304_633 n2_17304_666 2.095238e-02
R13787 n2_17304_666 n2_17304_849 1.161905e-01
R13788 n2_17304_849 n2_17304_882 2.095238e-02
R13789 n2_17304_882 n2_17304_1065 1.161905e-01
R13790 n2_17304_1065 n2_17304_1098 2.095238e-02
R13791 n2_17304_1098 n2_17304_1281 1.161905e-01
R13792 n2_17304_1281 n2_17304_1314 2.095238e-02
R13793 n2_17304_1314 n2_17304_1497 1.161905e-01
R13794 n2_17304_1497 n2_17304_1530 2.095238e-02
R13795 n2_17304_1530 n2_17304_1549 1.206349e-02
R13796 n2_17304_1549 n2_17304_1645 6.095238e-02
R13797 n2_17304_1645 n2_17304_1713 4.317460e-02
R13798 n2_17304_1713 n2_17304_1746 2.095238e-02
R13799 n2_17304_1746 n2_17304_1783 2.349206e-02
R13800 n2_17304_1783 n2_17304_1929 9.269841e-02
R13801 n2_17304_1929 n2_17304_1962 2.095238e-02
R13802 n2_17304_1962 n2_17304_2145 1.161905e-01
R13803 n2_17304_2145 n2_17304_2178 2.095238e-02
R13804 n2_17304_2178 n2_17304_2361 1.161905e-01
R13805 n2_17304_2361 n2_17304_2394 2.095238e-02
R13806 n2_17304_2394 n2_17304_2431 2.349206e-02
R13807 n2_17304_2431 n2_17304_2577 9.269841e-02
R13808 n2_17304_2577 n2_17304_2610 2.095238e-02
R13809 n2_17304_2610 n2_17304_2674 4.063492e-02
R13810 n2_17304_2674 n2_17304_2770 6.095238e-02
R13811 n2_17304_2770 n2_17304_2793 1.460317e-02
R13812 n2_17304_2793 n2_17304_2826 2.095238e-02
R13813 n2_17304_2826 n2_17304_2863 2.349206e-02
R13814 n2_17304_2863 n2_17304_3009 9.269841e-02
R13815 n2_17304_3009 n2_17304_3042 2.095238e-02
R13816 n2_17304_3042 n2_17304_3225 1.161905e-01
R13817 n2_17304_3225 n2_17304_3258 2.095238e-02
R13818 n2_17304_3258 n2_17304_3295 2.349206e-02
R13819 n2_17304_3295 n2_17304_3441 9.269841e-02
R13820 n2_17304_3441 n2_17304_3474 2.095238e-02
R13821 n2_17304_3474 n2_17304_3657 1.161905e-01
R13822 n2_17304_3657 n2_17304_3690 2.095238e-02
R13823 n2_17304_3690 n2_17304_3799 6.920635e-02
R13824 n2_17304_3799 n2_17304_3873 4.698413e-02
R13825 n2_17304_3873 n2_17304_3895 1.396825e-02
R13826 n2_17304_3895 n2_17304_3906 6.984127e-03
R13827 n2_17304_3906 n2_17304_4089 1.161905e-01
R13828 n2_17304_4089 n2_17304_4122 2.095238e-02
R13829 n2_17304_4122 n2_17304_4305 1.161905e-01
R13830 n2_17304_4305 n2_17304_4338 2.095238e-02
R13831 n2_17304_4338 n2_17304_4375 2.349206e-02
R13832 n2_17304_4375 n2_17304_4521 9.269841e-02
R13833 n2_17304_4521 n2_17304_4554 2.095238e-02
R13834 n2_17304_4554 n2_17304_4591 2.349206e-02
R13835 n2_17304_4591 n2_17304_4737 9.269841e-02
R13836 n2_17304_4737 n2_17304_4770 2.095238e-02
R13837 n2_17304_4770 n2_17304_4807 2.349206e-02
R13838 n2_17304_5169 n2_17304_5202 2.095238e-02
R13839 n2_17304_5202 n2_17304_5239 2.349206e-02
R13840 n2_17304_5239 n2_17304_5385 9.269841e-02
R13841 n2_17304_5385 n2_17304_5418 2.095238e-02
R13842 n2_17304_5418 n2_17304_5455 2.349206e-02
R13843 n2_17304_5455 n2_17304_5601 9.269841e-02
R13844 n2_17304_5601 n2_17304_5634 2.095238e-02
R13845 n2_17304_5634 n2_17304_5817 1.161905e-01
R13846 n2_17304_5817 n2_17304_5850 2.095238e-02
R13847 n2_17304_5850 n2_17304_6033 1.161905e-01
R13848 n2_17304_6033 n2_17304_6049 1.015873e-02
R13849 n2_17304_6049 n2_17304_6066 1.079365e-02
R13850 n2_17304_6066 n2_17304_6145 5.015873e-02
R13851 n2_17304_6145 n2_17304_6249 6.603175e-02
R13852 n2_17304_6249 n2_17304_6282 2.095238e-02
R13853 n2_17304_6282 n2_17304_6319 2.349206e-02
R13854 n2_17304_6319 n2_17304_6465 9.269841e-02
R13855 n2_17304_6465 n2_17304_6498 2.095238e-02
R13856 n2_17304_6498 n2_17304_6681 1.161905e-01
R13857 n2_17304_6681 n2_17304_6714 2.095238e-02
R13858 n2_17304_6714 n2_17304_6897 1.161905e-01
R13859 n2_17304_6897 n2_17304_6930 2.095238e-02
R13860 n2_17304_6930 n2_17304_7113 1.161905e-01
R13861 n2_17304_7329 n2_17304_7362 2.095238e-02
R13862 n2_17304_7362 n2_17304_7545 1.161905e-01
R13863 n2_17304_7545 n2_17304_7578 2.095238e-02
R13864 n2_17304_7578 n2_17304_7761 1.161905e-01
R13865 n2_17304_7761 n2_17304_7794 2.095238e-02
R13866 n2_17304_7794 n2_17304_7831 2.349206e-02
R13867 n2_17304_7831 n2_17304_7977 9.269841e-02
R13868 n2_17304_7977 n2_17304_8010 2.095238e-02
R13869 n2_17304_8010 n2_17304_8193 1.161905e-01
R13870 n2_17304_8193 n2_17304_8226 2.095238e-02
R13871 n2_17304_8226 n2_17304_8299 4.634921e-02
R13872 n2_17304_8299 n2_17304_8395 6.095238e-02
R13873 n2_17304_8395 n2_17304_8409 8.888889e-03
R13874 n2_17304_8409 n2_17304_8442 2.095238e-02
R13875 n2_17304_8442 n2_17304_8625 1.161905e-01
R13876 n2_17304_8625 n2_17304_8658 2.095238e-02
R13877 n2_17304_8658 n2_17304_8841 1.161905e-01
R13878 n2_17304_8841 n2_17304_8874 2.095238e-02
R13879 n2_17304_8874 n2_17304_8911 2.349206e-02
R13880 n2_17304_8911 n2_17304_9057 9.269841e-02
R13881 n2_17304_9057 n2_17304_9090 2.095238e-02
R13882 n2_17304_9090 n2_17304_9273 1.161905e-01
R13883 n2_17304_9273 n2_17304_9306 2.095238e-02
R13884 n2_17304_9705 n2_17304_9738 2.095238e-02
R13885 n2_17304_9738 n2_17304_9921 1.161905e-01
R13886 n2_17304_9921 n2_17304_9954 2.095238e-02
R13887 n2_17304_9954 n2_17304_9991 2.349206e-02
R13888 n2_17304_9991 n2_17304_10137 9.269841e-02
R13889 n2_17304_10137 n2_17304_10170 2.095238e-02
R13890 n2_17304_10170 n2_17304_10353 1.161905e-01
R13891 n2_17304_10353 n2_17304_10386 2.095238e-02
R13892 n2_17304_10386 n2_17304_10549 1.034921e-01
R13893 n2_17304_10549 n2_17304_10569 1.269841e-02
R13894 n2_17304_10569 n2_17304_10602 2.095238e-02
R13895 n2_17304_10602 n2_17304_10645 2.730159e-02
R13896 n2_17304_10645 n2_17304_10785 8.888889e-02
R13897 n2_17304_10785 n2_17304_10818 2.095238e-02
R13898 n2_17304_10818 n2_17304_11001 1.161905e-01
R13899 n2_17304_11001 n2_17304_11034 2.095238e-02
R13900 n2_17304_11034 n2_17304_11048 8.888889e-03
R13901 n2_17304_11048 n2_17304_11055 4.444444e-03
R13902 n2_17304_11055 n2_17304_11217 1.028571e-01
R13903 n2_17304_11217 n2_17304_11250 2.095238e-02
R13904 n2_17304_11250 n2_17304_11433 1.161905e-01
R13905 n2_17304_11433 n2_17304_11466 2.095238e-02
R13906 n2_17304_11865 n2_17304_11898 2.095238e-02
R13907 n2_17304_11898 n2_17304_12081 1.161905e-01
R13908 n2_17304_12081 n2_17304_12114 2.095238e-02
R13909 n2_17304_12114 n2_17304_12128 8.888889e-03
R13910 n2_17304_12128 n2_17304_12135 4.444444e-03
R13911 n2_17304_12135 n2_17304_12297 1.028571e-01
R13912 n2_17304_12297 n2_17304_12330 2.095238e-02
R13913 n2_17304_12330 n2_17304_12513 1.161905e-01
R13914 n2_17304_12513 n2_17304_12546 2.095238e-02
R13915 n2_17304_12546 n2_17304_12729 1.161905e-01
R13916 n2_17304_12729 n2_17304_12762 2.095238e-02
R13917 n2_17304_12762 n2_17304_12799 2.349206e-02
R13918 n2_17304_12799 n2_17304_12895 6.095238e-02
R13919 n2_17304_12895 n2_17304_12945 3.174603e-02
R13920 n2_17304_12945 n2_17304_12978 2.095238e-02
R13921 n2_17304_12978 n2_17304_13161 1.161905e-01
R13922 n2_17304_13161 n2_17304_13194 2.095238e-02
R13923 n2_17304_13194 n2_17304_13377 1.161905e-01
R13924 n2_17304_13377 n2_17304_13410 2.095238e-02
R13925 n2_17304_13410 n2_17304_13423 8.253968e-03
R13926 n2_17304_13423 n2_17304_13593 1.079365e-01
R13927 n2_17304_13593 n2_17304_13626 2.095238e-02
R13928 n2_17304_13626 n2_17304_13640 8.888889e-03
R13929 n2_17304_13640 n2_17304_13647 4.444444e-03
R13930 n2_17304_13647 n2_17304_13809 1.028571e-01
R13931 n2_17304_13809 n2_17304_13842 2.095238e-02
R13932 n2_17304_14241 n2_17304_14274 2.095238e-02
R13933 n2_17304_14274 n2_17304_14457 1.161905e-01
R13934 n2_17304_14457 n2_17304_14490 2.095238e-02
R13935 n2_17304_14490 n2_17304_14511 1.333333e-02
R13936 n2_17304_14511 n2_17304_14673 1.028571e-01
R13937 n2_17304_14673 n2_17304_14706 2.095238e-02
R13938 n2_17304_14706 n2_17304_14889 1.161905e-01
R13939 n2_17304_14889 n2_17304_14922 2.095238e-02
R13940 n2_17304_14922 n2_17304_14936 8.888889e-03
R13941 n2_17304_14936 n2_17304_14943 4.444444e-03
R13942 n2_17304_14943 n2_17304_15049 6.730159e-02
R13943 n2_17304_15049 n2_17304_15105 3.555556e-02
R13944 n2_17304_15105 n2_17304_15138 2.095238e-02
R13945 n2_17304_15138 n2_17304_15145 4.444444e-03
R13946 n2_17304_15145 n2_17304_15152 4.444444e-03
R13947 n2_17304_15152 n2_17304_15159 4.444444e-03
R13948 n2_17304_15159 n2_17304_15321 1.028571e-01
R13949 n2_17304_15321 n2_17304_15354 2.095238e-02
R13950 n2_17304_15354 n2_17304_15537 1.161905e-01
R13951 n2_17304_15537 n2_17304_15570 2.095238e-02
R13952 n2_17304_15570 n2_17304_15584 8.888889e-03
R13953 n2_17304_15584 n2_17304_15753 1.073016e-01
R13954 n2_17304_15753 n2_17304_15786 2.095238e-02
R13955 n2_17304_15786 n2_17304_15969 1.161905e-01
R13956 n2_17304_15969 n2_17304_16002 2.095238e-02
R13957 n2_17304_16401 n2_17304_16434 2.095238e-02
R13958 n2_17304_16434 n2_17304_16617 1.161905e-01
R13959 n2_17304_16617 n2_17304_16650 2.095238e-02
R13960 n2_17304_16650 n2_17304_16664 8.888889e-03
R13961 n2_17304_16664 n2_17304_16687 1.460317e-02
R13962 n2_17304_16687 n2_17304_16833 9.269841e-02
R13963 n2_17304_16833 n2_17304_16866 2.095238e-02
R13964 n2_17304_16866 n2_17304_17049 1.161905e-01
R13965 n2_17304_17049 n2_17304_17082 2.095238e-02
R13966 n2_17304_17082 n2_17304_17119 2.349206e-02
R13967 n2_17304_17119 n2_17304_17265 9.269841e-02
R13968 n2_17304_17265 n2_17304_17298 2.095238e-02
R13969 n2_17304_17298 n2_17304_17299 6.349206e-04
R13970 n2_17304_17299 n2_17304_17395 6.095238e-02
R13971 n2_17304_17395 n2_17304_17481 5.460317e-02
R13972 n2_17304_17481 n2_17304_17514 2.095238e-02
R13973 n2_17304_17514 n2_17304_17535 1.333333e-02
R13974 n2_17304_17535 n2_17304_17697 1.028571e-01
R13975 n2_17304_17697 n2_17304_17730 2.095238e-02
R13976 n2_17304_17730 n2_17304_17913 1.161905e-01
R13977 n2_17304_17913 n2_17304_17946 2.095238e-02
R13978 n2_17304_17946 n2_17304_18129 1.161905e-01
R13979 n2_17304_18129 n2_17304_18162 2.095238e-02
R13980 n2_17304_18162 n2_17304_18176 8.888889e-03
R13981 n2_17304_18176 n2_17304_18345 1.073016e-01
R13982 n2_17304_18345 n2_17304_18378 2.095238e-02
R13983 n2_17304_18378 n2_17304_18424 2.920635e-02
R13984 n2_17304_18424 n2_17304_18520 6.095238e-02
R13985 n2_17304_18520 n2_17304_18561 2.603175e-02
R13986 n2_17304_18561 n2_17304_18594 2.095238e-02
R13987 n2_17304_18594 n2_17304_18777 1.161905e-01
R13988 n2_17304_18777 n2_17304_18810 2.095238e-02
R13989 n2_17304_18810 n2_17304_18993 1.161905e-01
R13990 n2_17304_18993 n2_17304_19026 2.095238e-02
R13991 n2_17304_19026 n2_17304_19040 8.888889e-03
R13992 n2_17304_19040 n2_17304_19209 1.073016e-01
R13993 n2_17304_19209 n2_17304_19242 2.095238e-02
R13994 n2_17304_19242 n2_17304_19425 1.161905e-01
R13995 n2_17304_19425 n2_17304_19458 2.095238e-02
R13996 n2_17304_19458 n2_17304_19549 5.777778e-02
R13997 n2_17304_19549 n2_17304_19641 5.841270e-02
R13998 n2_17304_19641 n2_17304_19645 2.539683e-03
R13999 n2_17304_19645 n2_17304_19674 1.841270e-02
R14000 n2_17304_19674 n2_17304_19857 1.161905e-01
R14001 n2_17304_19857 n2_17304_19890 2.095238e-02
R14002 n2_17304_19890 n2_17304_20073 1.161905e-01
R14003 n2_17304_20073 n2_17304_20106 2.095238e-02
R14004 n2_17304_20106 n2_17304_20289 1.161905e-01
R14005 n2_17304_20289 n2_17304_20322 2.095238e-02
R14006 n2_17304_20322 n2_17304_20505 1.161905e-01
R14007 n2_17304_20505 n2_17304_20538 2.095238e-02
R14008 n2_17304_20538 n2_17304_20674 8.634921e-02
R14009 n2_17304_20674 n2_17304_20721 2.984127e-02
R14010 n2_17304_20721 n2_17304_20754 2.095238e-02
R14011 n2_17304_20754 n2_17304_20770 1.015873e-02
R14012 n2_17304_20770 n2_17304_20937 1.060317e-01
R14013 n2_17304_20937 n2_17304_20970 2.095238e-02
R14014 n2_17396_201 n2_17396_234 2.095238e-02
R14015 n2_17396_234 n2_17396_417 1.161905e-01
R14016 n2_17396_417 n2_17396_424 4.444444e-03
R14017 n2_17396_424 n2_17396_450 1.650794e-02
R14018 n2_17396_520 n2_17396_633 7.174603e-02
R14019 n2_17396_633 n2_17396_666 2.095238e-02
R14020 n2_17396_666 n2_17396_849 1.161905e-01
R14021 n2_17396_849 n2_17396_882 2.095238e-02
R14022 n2_17396_882 n2_17396_1065 1.161905e-01
R14023 n2_17396_1065 n2_17396_1098 2.095238e-02
R14024 n2_17396_1098 n2_17396_1281 1.161905e-01
R14025 n2_17396_1281 n2_17396_1314 2.095238e-02
R14026 n2_17396_1314 n2_17396_1497 1.161905e-01
R14027 n2_17396_1497 n2_17396_1530 2.095238e-02
R14028 n2_17396_1530 n2_17396_1549 1.206349e-02
R14029 n2_17396_1645 n2_17396_1713 4.317460e-02
R14030 n2_17396_1713 n2_17396_1746 2.095238e-02
R14031 n2_17396_1746 n2_17396_1783 2.349206e-02
R14032 n2_17396_1783 n2_17396_1929 9.269841e-02
R14033 n2_17396_1929 n2_17396_1962 2.095238e-02
R14034 n2_17396_1962 n2_17396_2145 1.161905e-01
R14035 n2_17396_2145 n2_17396_2178 2.095238e-02
R14036 n2_17396_2178 n2_17396_2361 1.161905e-01
R14037 n2_17396_2361 n2_17396_2394 2.095238e-02
R14038 n2_17396_2394 n2_17396_2431 2.349206e-02
R14039 n2_17396_2431 n2_17396_2577 9.269841e-02
R14040 n2_17396_2577 n2_17396_2610 2.095238e-02
R14041 n2_17396_2610 n2_17396_2674 4.063492e-02
R14042 n2_17396_2770 n2_17396_2793 1.460317e-02
R14043 n2_17396_2793 n2_17396_2826 2.095238e-02
R14044 n2_17396_2826 n2_17396_2863 2.349206e-02
R14045 n2_17396_2863 n2_17396_3009 9.269841e-02
R14046 n2_17396_3009 n2_17396_3042 2.095238e-02
R14047 n2_17396_3042 n2_17396_3225 1.161905e-01
R14048 n2_17396_3225 n2_17396_3258 2.095238e-02
R14049 n2_17396_3258 n2_17396_3295 2.349206e-02
R14050 n2_17396_3295 n2_17396_3441 9.269841e-02
R14051 n2_17396_3441 n2_17396_3474 2.095238e-02
R14052 n2_17396_3474 n2_17396_3657 1.161905e-01
R14053 n2_17396_3657 n2_17396_3690 2.095238e-02
R14054 n2_17396_3690 n2_17396_3799 6.920635e-02
R14055 n2_17396_17395 n2_17396_17481 5.460317e-02
R14056 n2_17396_17481 n2_17396_17514 2.095238e-02
R14057 n2_17396_17514 n2_17396_17535 1.333333e-02
R14058 n2_17396_17535 n2_17396_17697 1.028571e-01
R14059 n2_17396_17697 n2_17396_17730 2.095238e-02
R14060 n2_17396_17730 n2_17396_17913 1.161905e-01
R14061 n2_17396_17913 n2_17396_17946 2.095238e-02
R14062 n2_17396_17946 n2_17396_18129 1.161905e-01
R14063 n2_17396_18129 n2_17396_18162 2.095238e-02
R14064 n2_17396_18162 n2_17396_18176 8.888889e-03
R14065 n2_17396_18176 n2_17396_18345 1.073016e-01
R14066 n2_17396_18345 n2_17396_18378 2.095238e-02
R14067 n2_17396_18378 n2_17396_18424 2.920635e-02
R14068 n2_17396_18520 n2_17396_18561 2.603175e-02
R14069 n2_17396_18561 n2_17396_18594 2.095238e-02
R14070 n2_17396_18594 n2_17396_18777 1.161905e-01
R14071 n2_17396_18777 n2_17396_18810 2.095238e-02
R14072 n2_17396_18810 n2_17396_18993 1.161905e-01
R14073 n2_17396_18993 n2_17396_19026 2.095238e-02
R14074 n2_17396_19026 n2_17396_19040 8.888889e-03
R14075 n2_17396_19040 n2_17396_19209 1.073016e-01
R14076 n2_17396_19209 n2_17396_19242 2.095238e-02
R14077 n2_17396_19242 n2_17396_19425 1.161905e-01
R14078 n2_17396_19425 n2_17396_19458 2.095238e-02
R14079 n2_17396_19458 n2_17396_19549 5.777778e-02
R14080 n2_17396_19641 n2_17396_19645 2.539683e-03
R14081 n2_17396_19645 n2_17396_19674 1.841270e-02
R14082 n2_17396_19674 n2_17396_19857 1.161905e-01
R14083 n2_17396_19857 n2_17396_19890 2.095238e-02
R14084 n2_17396_19890 n2_17396_20073 1.161905e-01
R14085 n2_17396_20073 n2_17396_20106 2.095238e-02
R14086 n2_17396_20106 n2_17396_20289 1.161905e-01
R14087 n2_17396_20289 n2_17396_20322 2.095238e-02
R14088 n2_17396_20322 n2_17396_20505 1.161905e-01
R14089 n2_17396_20505 n2_17396_20538 2.095238e-02
R14090 n2_17396_20538 n2_17396_20674 8.634921e-02
R14091 n2_17396_20754 n2_17396_20770 1.015873e-02
R14092 n2_17396_20770 n2_17396_20937 1.060317e-01
R14093 n2_17396_20937 n2_17396_20970 2.095238e-02
R14094 n2_18241_2793 n2_18241_2826 2.095238e-02
R14095 n2_18241_2826 n2_18241_3009 1.161905e-01
R14096 n2_18241_3009 n2_18241_3042 2.095238e-02
R14097 n2_18241_3042 n2_18241_3225 1.161905e-01
R14098 n2_18241_3225 n2_18241_3258 2.095238e-02
R14099 n2_18241_3258 n2_18241_3295 2.349206e-02
R14100 n2_18241_3295 n2_18241_3441 9.269841e-02
R14101 n2_18241_3441 n2_18241_3474 2.095238e-02
R14102 n2_18241_3474 n2_18241_3657 1.161905e-01
R14103 n2_18241_3657 n2_18241_3690 2.095238e-02
R14104 n2_18241_3690 n2_18241_3799 6.920635e-02
R14105 n2_18241_3873 n2_18241_3895 1.396825e-02
R14106 n2_18241_3895 n2_18241_3906 6.984127e-03
R14107 n2_18241_3906 n2_18241_4089 1.161905e-01
R14108 n2_18241_4089 n2_18241_4122 2.095238e-02
R14109 n2_18241_4122 n2_18241_4305 1.161905e-01
R14110 n2_18241_4305 n2_18241_4338 2.095238e-02
R14111 n2_18241_4338 n2_18241_4375 2.349206e-02
R14112 n2_18241_4375 n2_18241_4521 9.269841e-02
R14113 n2_18241_4521 n2_18241_4554 2.095238e-02
R14114 n2_18241_4554 n2_18241_4591 2.349206e-02
R14115 n2_18241_4591 n2_18241_4737 9.269841e-02
R14116 n2_18241_4737 n2_18241_4770 2.095238e-02
R14117 n2_18241_4770 n2_18241_4807 2.349206e-02
R14118 n2_18241_4807 n2_18241_4953 9.269841e-02
R14119 n2_18241_4953 n2_18241_4986 2.095238e-02
R14120 n2_18241_4986 n2_18241_5023 2.349206e-02
R14121 n2_18241_5023 n2_18241_5169 9.269841e-02
R14122 n2_18241_5169 n2_18241_5202 2.095238e-02
R14123 n2_18241_5202 n2_18241_5239 2.349206e-02
R14124 n2_18241_5239 n2_18241_5385 9.269841e-02
R14125 n2_18241_5385 n2_18241_5418 2.095238e-02
R14126 n2_18241_5418 n2_18241_5455 2.349206e-02
R14127 n2_18241_5455 n2_18241_5601 9.269841e-02
R14128 n2_18241_5601 n2_18241_5634 2.095238e-02
R14129 n2_18241_5634 n2_18241_5817 1.161905e-01
R14130 n2_18241_5817 n2_18241_5850 2.095238e-02
R14131 n2_18241_5850 n2_18241_6033 1.161905e-01
R14132 n2_18241_6033 n2_18241_6049 1.015873e-02
R14133 n2_18241_6049 n2_18241_6066 1.079365e-02
R14134 n2_18241_6145 n2_18241_6249 6.603175e-02
R14135 n2_18241_6249 n2_18241_6282 2.095238e-02
R14136 n2_18241_6282 n2_18241_6319 2.349206e-02
R14137 n2_18241_6319 n2_18241_6465 9.269841e-02
R14138 n2_18241_6465 n2_18241_6498 2.095238e-02
R14139 n2_18241_6498 n2_18241_6681 1.161905e-01
R14140 n2_18241_6681 n2_18241_6714 2.095238e-02
R14141 n2_18241_6714 n2_18241_6897 1.161905e-01
R14142 n2_18241_6897 n2_18241_6930 2.095238e-02
R14143 n2_18241_6930 n2_18241_7113 1.161905e-01
R14144 n2_18241_7113 n2_18241_7146 2.095238e-02
R14145 n2_18241_7146 n2_18241_7329 1.161905e-01
R14146 n2_18241_7329 n2_18241_7362 2.095238e-02
R14147 n2_18241_7362 n2_18241_7545 1.161905e-01
R14148 n2_18241_7545 n2_18241_7578 2.095238e-02
R14149 n2_18241_7578 n2_18241_7761 1.161905e-01
R14150 n2_18241_7761 n2_18241_7794 2.095238e-02
R14151 n2_18241_7794 n2_18241_7831 2.349206e-02
R14152 n2_18241_7831 n2_18241_7977 9.269841e-02
R14153 n2_18241_7977 n2_18241_8010 2.095238e-02
R14154 n2_18241_8010 n2_18241_8193 1.161905e-01
R14155 n2_18241_8193 n2_18241_8226 2.095238e-02
R14156 n2_18241_8226 n2_18241_8299 4.634921e-02
R14157 n2_18241_8395 n2_18241_8409 8.888889e-03
R14158 n2_18241_8409 n2_18241_8442 2.095238e-02
R14159 n2_18241_8442 n2_18241_8625 1.161905e-01
R14160 n2_18241_8625 n2_18241_8658 2.095238e-02
R14161 n2_18241_8658 n2_18241_8841 1.161905e-01
R14162 n2_18241_8841 n2_18241_8874 2.095238e-02
R14163 n2_18241_8874 n2_18241_8911 2.349206e-02
R14164 n2_18241_8911 n2_18241_9057 9.269841e-02
R14165 n2_18241_9057 n2_18241_9090 2.095238e-02
R14166 n2_18241_9090 n2_18241_9273 1.161905e-01
R14167 n2_18241_9273 n2_18241_9306 2.095238e-02
R14168 n2_18241_9306 n2_18241_9489 1.161905e-01
R14169 n2_18241_9489 n2_18241_9522 2.095238e-02
R14170 n2_18241_9522 n2_18241_9705 1.161905e-01
R14171 n2_18241_9705 n2_18241_9738 2.095238e-02
R14172 n2_18241_9738 n2_18241_9921 1.161905e-01
R14173 n2_18241_9921 n2_18241_9954 2.095238e-02
R14174 n2_18241_9954 n2_18241_9991 2.349206e-02
R14175 n2_18241_9991 n2_18241_10137 9.269841e-02
R14176 n2_18241_10137 n2_18241_10170 2.095238e-02
R14177 n2_18241_10170 n2_18241_10353 1.161905e-01
R14178 n2_18241_10353 n2_18241_10386 2.095238e-02
R14179 n2_18241_10386 n2_18241_10549 1.034921e-01
R14180 n2_18241_10549 n2_18241_10569 1.269841e-02
R14181 n2_18241_10645 n2_18241_10785 8.888889e-02
R14182 n2_18241_10785 n2_18241_10818 2.095238e-02
R14183 n2_18241_10818 n2_18241_11001 1.161905e-01
R14184 n2_18241_11001 n2_18241_11034 2.095238e-02
R14185 n2_18241_11034 n2_18241_11055 1.333333e-02
R14186 n2_18241_11055 n2_18241_11217 1.028571e-01
R14187 n2_18241_11217 n2_18241_11250 2.095238e-02
R14188 n2_18241_11250 n2_18241_11433 1.161905e-01
R14189 n2_18241_11433 n2_18241_11466 2.095238e-02
R14190 n2_18241_11466 n2_18241_11649 1.161905e-01
R14191 n2_18241_11649 n2_18241_11682 2.095238e-02
R14192 n2_18241_11682 n2_18241_11865 1.161905e-01
R14193 n2_18241_11865 n2_18241_11898 2.095238e-02
R14194 n2_18241_11898 n2_18241_12081 1.161905e-01
R14195 n2_18241_12081 n2_18241_12114 2.095238e-02
R14196 n2_18241_12114 n2_18241_12128 8.888889e-03
R14197 n2_18241_12128 n2_18241_12297 1.073016e-01
R14198 n2_18241_12297 n2_18241_12330 2.095238e-02
R14199 n2_18241_12330 n2_18241_12513 1.161905e-01
R14200 n2_18241_12513 n2_18241_12546 2.095238e-02
R14201 n2_18241_12546 n2_18241_12729 1.161905e-01
R14202 n2_18241_12729 n2_18241_12762 2.095238e-02
R14203 n2_18241_12762 n2_18241_12799 2.349206e-02
R14204 n2_18241_12895 n2_18241_12945 3.174603e-02
R14205 n2_18241_12945 n2_18241_12978 2.095238e-02
R14206 n2_18241_12978 n2_18241_13161 1.161905e-01
R14207 n2_18241_13161 n2_18241_13194 2.095238e-02
R14208 n2_18241_13194 n2_18241_13377 1.161905e-01
R14209 n2_18241_13377 n2_18241_13410 2.095238e-02
R14210 n2_18241_13410 n2_18241_13593 1.161905e-01
R14211 n2_18241_13593 n2_18241_13626 2.095238e-02
R14212 n2_18241_13626 n2_18241_13640 8.888889e-03
R14213 n2_18241_13640 n2_18241_13647 4.444444e-03
R14214 n2_18241_13647 n2_18241_13809 1.028571e-01
R14215 n2_18241_13809 n2_18241_13842 2.095238e-02
R14216 n2_18241_13842 n2_18241_14025 1.161905e-01
R14217 n2_18241_14025 n2_18241_14058 2.095238e-02
R14218 n2_18241_14058 n2_18241_14241 1.161905e-01
R14219 n2_18241_14241 n2_18241_14274 2.095238e-02
R14220 n2_18241_14274 n2_18241_14457 1.161905e-01
R14221 n2_18241_14457 n2_18241_14490 2.095238e-02
R14222 n2_18241_14490 n2_18241_14504 8.888889e-03
R14223 n2_18241_14504 n2_18241_14511 4.444444e-03
R14224 n2_18241_14511 n2_18241_14673 1.028571e-01
R14225 n2_18241_14673 n2_18241_14706 2.095238e-02
R14226 n2_18241_14706 n2_18241_14889 1.161905e-01
R14227 n2_18241_14889 n2_18241_14922 2.095238e-02
R14228 n2_18241_14922 n2_18241_14936 8.888889e-03
R14229 n2_18241_14936 n2_18241_15049 7.174603e-02
R14230 n2_18241_15138 n2_18241_15145 4.444444e-03
R14231 n2_18241_15145 n2_18241_15152 4.444444e-03
R14232 n2_18241_15152 n2_18241_15321 1.073016e-01
R14233 n2_18241_15321 n2_18241_15354 2.095238e-02
R14234 n2_18241_15354 n2_18241_15537 1.161905e-01
R14235 n2_18241_15537 n2_18241_15570 2.095238e-02
R14236 n2_18241_15570 n2_18241_15584 8.888889e-03
R14237 n2_18241_15584 n2_18241_15753 1.073016e-01
R14238 n2_18241_15753 n2_18241_15786 2.095238e-02
R14239 n2_18241_15786 n2_18241_15969 1.161905e-01
R14240 n2_18241_15969 n2_18241_16002 2.095238e-02
R14241 n2_18241_16002 n2_18241_16185 1.161905e-01
R14242 n2_18241_16185 n2_18241_16218 2.095238e-02
R14243 n2_18241_16218 n2_18241_16401 1.161905e-01
R14244 n2_18241_16401 n2_18241_16434 2.095238e-02
R14245 n2_18241_16434 n2_18241_16617 1.161905e-01
R14246 n2_18241_16617 n2_18241_16650 2.095238e-02
R14247 n2_18241_16650 n2_18241_16664 8.888889e-03
R14248 n2_18241_16664 n2_18241_16671 4.444444e-03
R14249 n2_18241_16671 n2_18241_16833 1.028571e-01
R14250 n2_18241_16833 n2_18241_16866 2.095238e-02
R14251 n2_18241_16866 n2_18241_17049 1.161905e-01
R14252 n2_18241_17049 n2_18241_17082 2.095238e-02
R14253 n2_18241_17082 n2_18241_17119 2.349206e-02
R14254 n2_18241_17119 n2_18241_17265 9.269841e-02
R14255 n2_18241_17265 n2_18241_17298 2.095238e-02
R14256 n2_18241_17298 n2_18241_17299 6.349206e-04
R14257 n2_18241_17395 n2_18241_17481 5.460317e-02
R14258 n2_18241_17481 n2_18241_17514 2.095238e-02
R14259 n2_18241_17514 n2_18241_17697 1.161905e-01
R14260 n2_18241_17697 n2_18241_17730 2.095238e-02
R14261 n2_18241_17730 n2_18241_17744 8.888889e-03
R14262 n2_18241_17744 n2_18241_17913 1.073016e-01
R14263 n2_18241_17913 n2_18241_17946 2.095238e-02
R14264 n2_18241_17946 n2_18241_18129 1.161905e-01
R14265 n2_18241_18129 n2_18241_18162 2.095238e-02
R14266 n2_18241_18162 n2_18241_18345 1.161905e-01
R14267 n2_18241_18345 n2_18241_18378 2.095238e-02
R14268 n2_18241_3799 n2_18380_3799 8.825397e-02
R14269 n2_18380_3799 n2_18429_3799 3.111111e-02
R14270 n2_18241_3895 n2_18380_3895 8.825397e-02
R14271 n2_18380_3895 n2_18429_3895 3.111111e-02
R14272 n2_18241_6049 n2_18380_6049 8.825397e-02
R14273 n2_18380_6049 n2_18429_6049 3.111111e-02
R14274 n2_18241_6145 n2_18380_6145 8.825397e-02
R14275 n2_18380_6145 n2_18429_6145 3.111111e-02
R14276 n2_18241_8299 n2_18380_8299 8.825397e-02
R14277 n2_18380_8299 n2_18429_8299 3.111111e-02
R14278 n2_18241_8395 n2_18380_8395 8.825397e-02
R14279 n2_18380_8395 n2_18429_8395 3.111111e-02
R14280 n2_18241_10549 n2_18380_10549 8.825397e-02
R14281 n2_18380_10549 n2_18429_10549 3.111111e-02
R14282 n2_18241_10645 n2_18380_10645 8.825397e-02
R14283 n2_18380_10645 n2_18429_10645 3.111111e-02
R14284 n2_18241_12799 n2_18380_12799 8.825397e-02
R14285 n2_18380_12799 n2_18429_12799 3.111111e-02
R14286 n2_18241_12895 n2_18380_12895 8.825397e-02
R14287 n2_18380_12895 n2_18429_12895 3.111111e-02
R14288 n2_18241_15049 n2_18380_15049 8.825397e-02
R14289 n2_18380_15049 n2_18429_15049 3.111111e-02
R14290 n2_18241_15145 n2_18380_15145 8.825397e-02
R14291 n2_18380_15145 n2_18429_15145 3.111111e-02
R14292 n2_18241_17299 n2_18380_17299 8.825397e-02
R14293 n2_18380_17299 n2_18429_17299 3.111111e-02
R14294 n2_18241_17395 n2_18380_17395 8.825397e-02
R14295 n2_18380_17395 n2_18429_17395 3.111111e-02
R14296 n2_18429_2826 n2_18429_3009 1.161905e-01
R14297 n2_18429_3009 n2_18429_3042 2.095238e-02
R14298 n2_18429_3042 n2_18429_3225 1.161905e-01
R14299 n2_18429_3225 n2_18429_3258 2.095238e-02
R14300 n2_18429_3258 n2_18429_3295 2.349206e-02
R14301 n2_18429_3295 n2_18429_3441 9.269841e-02
R14302 n2_18429_3441 n2_18429_3474 2.095238e-02
R14303 n2_18429_3474 n2_18429_3657 1.161905e-01
R14304 n2_18429_3657 n2_18429_3690 2.095238e-02
R14305 n2_18429_3690 n2_18429_3799 6.920635e-02
R14306 n2_18429_3799 n2_18429_3873 4.698413e-02
R14307 n2_18429_3873 n2_18429_3895 1.396825e-02
R14308 n2_18429_3895 n2_18429_3906 6.984127e-03
R14309 n2_18429_3906 n2_18429_4089 1.161905e-01
R14310 n2_18429_4089 n2_18429_4122 2.095238e-02
R14311 n2_18429_4122 n2_18429_4305 1.161905e-01
R14312 n2_18429_4305 n2_18429_4338 2.095238e-02
R14313 n2_18429_4338 n2_18429_4375 2.349206e-02
R14314 n2_18429_4375 n2_18429_4521 9.269841e-02
R14315 n2_18429_4521 n2_18429_4554 2.095238e-02
R14316 n2_18429_4554 n2_18429_4591 2.349206e-02
R14317 n2_18429_4591 n2_18429_4737 9.269841e-02
R14318 n2_18429_4737 n2_18429_4770 2.095238e-02
R14319 n2_18429_4770 n2_18429_4807 2.349206e-02
R14320 n2_18429_5169 n2_18429_5202 2.095238e-02
R14321 n2_18429_5202 n2_18429_5239 2.349206e-02
R14322 n2_18429_5239 n2_18429_5385 9.269841e-02
R14323 n2_18429_5385 n2_18429_5418 2.095238e-02
R14324 n2_18429_5418 n2_18429_5455 2.349206e-02
R14325 n2_18429_5455 n2_18429_5601 9.269841e-02
R14326 n2_18429_5601 n2_18429_5634 2.095238e-02
R14327 n2_18429_5634 n2_18429_5817 1.161905e-01
R14328 n2_18429_5817 n2_18429_5850 2.095238e-02
R14329 n2_18429_5850 n2_18429_6033 1.161905e-01
R14330 n2_18429_6033 n2_18429_6049 1.015873e-02
R14331 n2_18429_6049 n2_18429_6066 1.079365e-02
R14332 n2_18429_6066 n2_18429_6145 5.015873e-02
R14333 n2_18429_6145 n2_18429_6249 6.603175e-02
R14334 n2_18429_6249 n2_18429_6282 2.095238e-02
R14335 n2_18429_6282 n2_18429_6319 2.349206e-02
R14336 n2_18429_6319 n2_18429_6465 9.269841e-02
R14337 n2_18429_6465 n2_18429_6498 2.095238e-02
R14338 n2_18429_6498 n2_18429_6681 1.161905e-01
R14339 n2_18429_6681 n2_18429_6714 2.095238e-02
R14340 n2_18429_6714 n2_18429_6897 1.161905e-01
R14341 n2_18429_6897 n2_18429_6930 2.095238e-02
R14342 n2_18429_6930 n2_18429_7113 1.161905e-01
R14343 n2_18429_7329 n2_18429_7362 2.095238e-02
R14344 n2_18429_7362 n2_18429_7545 1.161905e-01
R14345 n2_18429_7545 n2_18429_7578 2.095238e-02
R14346 n2_18429_7578 n2_18429_7761 1.161905e-01
R14347 n2_18429_7761 n2_18429_7794 2.095238e-02
R14348 n2_18429_7794 n2_18429_7831 2.349206e-02
R14349 n2_18429_7831 n2_18429_7977 9.269841e-02
R14350 n2_18429_7977 n2_18429_8010 2.095238e-02
R14351 n2_18429_8010 n2_18429_8193 1.161905e-01
R14352 n2_18429_8193 n2_18429_8226 2.095238e-02
R14353 n2_18429_8226 n2_18429_8299 4.634921e-02
R14354 n2_18429_8299 n2_18429_8395 6.095238e-02
R14355 n2_18429_8395 n2_18429_8409 8.888889e-03
R14356 n2_18429_8409 n2_18429_8442 2.095238e-02
R14357 n2_18429_8442 n2_18429_8625 1.161905e-01
R14358 n2_18429_8625 n2_18429_8658 2.095238e-02
R14359 n2_18429_8658 n2_18429_8841 1.161905e-01
R14360 n2_18429_8841 n2_18429_8874 2.095238e-02
R14361 n2_18429_8874 n2_18429_8911 2.349206e-02
R14362 n2_18429_8911 n2_18429_9057 9.269841e-02
R14363 n2_18429_9057 n2_18429_9090 2.095238e-02
R14364 n2_18429_9090 n2_18429_9273 1.161905e-01
R14365 n2_18429_9273 n2_18429_9306 2.095238e-02
R14366 n2_18429_9705 n2_18429_9738 2.095238e-02
R14367 n2_18429_9738 n2_18429_9921 1.161905e-01
R14368 n2_18429_9921 n2_18429_9954 2.095238e-02
R14369 n2_18429_9954 n2_18429_9991 2.349206e-02
R14370 n2_18429_9991 n2_18429_10137 9.269841e-02
R14371 n2_18429_10137 n2_18429_10170 2.095238e-02
R14372 n2_18429_10170 n2_18429_10353 1.161905e-01
R14373 n2_18429_10353 n2_18429_10386 2.095238e-02
R14374 n2_18429_10386 n2_18429_10549 1.034921e-01
R14375 n2_18429_10549 n2_18429_10569 1.269841e-02
R14376 n2_18429_10569 n2_18429_10602 2.095238e-02
R14377 n2_18429_10602 n2_18429_10645 2.730159e-02
R14378 n2_18429_10645 n2_18429_10785 8.888889e-02
R14379 n2_18429_10785 n2_18429_10818 2.095238e-02
R14380 n2_18429_10818 n2_18429_11001 1.161905e-01
R14381 n2_18429_11001 n2_18429_11034 2.095238e-02
R14382 n2_18429_11034 n2_18429_11055 1.333333e-02
R14383 n2_18429_11055 n2_18429_11217 1.028571e-01
R14384 n2_18429_11217 n2_18429_11250 2.095238e-02
R14385 n2_18429_11250 n2_18429_11433 1.161905e-01
R14386 n2_18429_11433 n2_18429_11466 2.095238e-02
R14387 n2_18429_11865 n2_18429_11898 2.095238e-02
R14388 n2_18429_11898 n2_18429_12081 1.161905e-01
R14389 n2_18429_12081 n2_18429_12114 2.095238e-02
R14390 n2_18429_12114 n2_18429_12128 8.888889e-03
R14391 n2_18429_12128 n2_18429_12297 1.073016e-01
R14392 n2_18429_12297 n2_18429_12330 2.095238e-02
R14393 n2_18429_12330 n2_18429_12513 1.161905e-01
R14394 n2_18429_12513 n2_18429_12546 2.095238e-02
R14395 n2_18429_12546 n2_18429_12729 1.161905e-01
R14396 n2_18429_12729 n2_18429_12762 2.095238e-02
R14397 n2_18429_12762 n2_18429_12799 2.349206e-02
R14398 n2_18429_12799 n2_18429_12895 6.095238e-02
R14399 n2_18429_12895 n2_18429_12945 3.174603e-02
R14400 n2_18429_12945 n2_18429_12978 2.095238e-02
R14401 n2_18429_12978 n2_18429_13161 1.161905e-01
R14402 n2_18429_13161 n2_18429_13194 2.095238e-02
R14403 n2_18429_13194 n2_18429_13377 1.161905e-01
R14404 n2_18429_13377 n2_18429_13410 2.095238e-02
R14405 n2_18429_13410 n2_18429_13423 8.253968e-03
R14406 n2_18429_13423 n2_18429_13593 1.079365e-01
R14407 n2_18429_13593 n2_18429_13626 2.095238e-02
R14408 n2_18429_13626 n2_18429_13640 8.888889e-03
R14409 n2_18429_13640 n2_18429_13647 4.444444e-03
R14410 n2_18429_13647 n2_18429_13809 1.028571e-01
R14411 n2_18429_13809 n2_18429_13842 2.095238e-02
R14412 n2_18429_14241 n2_18429_14274 2.095238e-02
R14413 n2_18429_14274 n2_18429_14457 1.161905e-01
R14414 n2_18429_14457 n2_18429_14490 2.095238e-02
R14415 n2_18429_14490 n2_18429_14504 8.888889e-03
R14416 n2_18429_14504 n2_18429_14511 4.444444e-03
R14417 n2_18429_14511 n2_18429_14673 1.028571e-01
R14418 n2_18429_14673 n2_18429_14706 2.095238e-02
R14419 n2_18429_14706 n2_18429_14889 1.161905e-01
R14420 n2_18429_14889 n2_18429_14922 2.095238e-02
R14421 n2_18429_14922 n2_18429_14936 8.888889e-03
R14422 n2_18429_14936 n2_18429_15049 7.174603e-02
R14423 n2_18429_15049 n2_18429_15105 3.555556e-02
R14424 n2_18429_15105 n2_18429_15138 2.095238e-02
R14425 n2_18429_15138 n2_18429_15145 4.444444e-03
R14426 n2_18429_15145 n2_18429_15152 4.444444e-03
R14427 n2_18429_15152 n2_18429_15321 1.073016e-01
R14428 n2_18429_15321 n2_18429_15354 2.095238e-02
R14429 n2_18429_15354 n2_18429_15537 1.161905e-01
R14430 n2_18429_15537 n2_18429_15570 2.095238e-02
R14431 n2_18429_15570 n2_18429_15584 8.888889e-03
R14432 n2_18429_15584 n2_18429_15753 1.073016e-01
R14433 n2_18429_15753 n2_18429_15786 2.095238e-02
R14434 n2_18429_15786 n2_18429_15969 1.161905e-01
R14435 n2_18429_15969 n2_18429_16002 2.095238e-02
R14436 n2_18429_16401 n2_18429_16434 2.095238e-02
R14437 n2_18429_16434 n2_18429_16617 1.161905e-01
R14438 n2_18429_16617 n2_18429_16650 2.095238e-02
R14439 n2_18429_16650 n2_18429_16664 8.888889e-03
R14440 n2_18429_16664 n2_18429_16671 4.444444e-03
R14441 n2_18429_16671 n2_18429_16833 1.028571e-01
R14442 n2_18429_16833 n2_18429_16866 2.095238e-02
R14443 n2_18429_16866 n2_18429_17049 1.161905e-01
R14444 n2_18429_17049 n2_18429_17082 2.095238e-02
R14445 n2_18429_17082 n2_18429_17119 2.349206e-02
R14446 n2_18429_17119 n2_18429_17265 9.269841e-02
R14447 n2_18429_17265 n2_18429_17298 2.095238e-02
R14448 n2_18429_17298 n2_18429_17299 6.349206e-04
R14449 n2_18429_17299 n2_18429_17395 6.095238e-02
R14450 n2_18429_17395 n2_18429_17481 5.460317e-02
R14451 n2_18429_17481 n2_18429_17514 2.095238e-02
R14452 n2_18429_17514 n2_18429_17697 1.161905e-01
R14453 n2_18429_17697 n2_18429_17730 2.095238e-02
R14454 n2_18429_17730 n2_18429_17744 8.888889e-03
R14455 n2_18429_17744 n2_18429_17913 1.073016e-01
R14456 n2_18429_17913 n2_18429_17946 2.095238e-02
R14457 n2_18429_17946 n2_18429_18129 1.161905e-01
R14458 n2_18429_18129 n2_18429_18162 2.095238e-02
R14459 n2_18429_18162 n2_18429_18345 1.161905e-01
R14460 n2_19366_201 n2_19366_234 2.095238e-02
R14461 n2_19366_234 n2_19366_417 1.161905e-01
R14462 n2_19366_417 n2_19366_424 4.444444e-03
R14463 n2_19366_424 n2_19366_450 1.650794e-02
R14464 n2_19366_520 n2_19366_633 7.174603e-02
R14465 n2_19366_633 n2_19366_666 2.095238e-02
R14466 n2_19366_666 n2_19366_849 1.161905e-01
R14467 n2_19366_849 n2_19366_882 2.095238e-02
R14468 n2_19366_882 n2_19366_1065 1.161905e-01
R14469 n2_19366_1065 n2_19366_1098 2.095238e-02
R14470 n2_19366_1098 n2_19366_1281 1.161905e-01
R14471 n2_19366_1281 n2_19366_1314 2.095238e-02
R14472 n2_19366_1314 n2_19366_1497 1.161905e-01
R14473 n2_19366_1497 n2_19366_1530 2.095238e-02
R14474 n2_19366_1530 n2_19366_1713 1.161905e-01
R14475 n2_19366_1713 n2_19366_1746 2.095238e-02
R14476 n2_19366_1746 n2_19366_1929 1.161905e-01
R14477 n2_19366_1929 n2_19366_1962 2.095238e-02
R14478 n2_19366_1962 n2_19366_1976 8.888889e-03
R14479 n2_19366_1976 n2_19366_1999 1.460317e-02
R14480 n2_19366_1999 n2_19366_2145 9.269841e-02
R14481 n2_19366_2145 n2_19366_2178 2.095238e-02
R14482 n2_19366_2178 n2_19366_2361 1.161905e-01
R14483 n2_19366_2361 n2_19366_2394 2.095238e-02
R14484 n2_19366_2394 n2_19366_2577 1.161905e-01
R14485 n2_19366_2577 n2_19366_2610 2.095238e-02
R14486 n2_19366_2610 n2_19366_2793 1.161905e-01
R14487 n2_19366_2793 n2_19366_2826 2.095238e-02
R14488 n2_19366_2826 n2_19366_3009 1.161905e-01
R14489 n2_19366_3009 n2_19366_3042 2.095238e-02
R14490 n2_19366_3042 n2_19366_3225 1.161905e-01
R14491 n2_19366_3225 n2_19366_3258 2.095238e-02
R14492 n2_19366_3258 n2_19366_3295 2.349206e-02
R14493 n2_19366_3295 n2_19366_3441 9.269841e-02
R14494 n2_19366_3441 n2_19366_3474 2.095238e-02
R14495 n2_19366_3474 n2_19366_3657 1.161905e-01
R14496 n2_19366_3657 n2_19366_3690 2.095238e-02
R14497 n2_19366_3690 n2_19366_3799 6.920635e-02
R14498 n2_19366_3873 n2_19366_3895 1.396825e-02
R14499 n2_19366_3895 n2_19366_3906 6.984127e-03
R14500 n2_19366_3906 n2_19366_4089 1.161905e-01
R14501 n2_19366_4089 n2_19366_4122 2.095238e-02
R14502 n2_19366_4122 n2_19366_4305 1.161905e-01
R14503 n2_19366_4305 n2_19366_4338 2.095238e-02
R14504 n2_19366_4338 n2_19366_4375 2.349206e-02
R14505 n2_19366_4375 n2_19366_4521 9.269841e-02
R14506 n2_19366_4521 n2_19366_4554 2.095238e-02
R14507 n2_19366_4554 n2_19366_4737 1.161905e-01
R14508 n2_19366_4737 n2_19366_4770 2.095238e-02
R14509 n2_19366_4770 n2_19366_4953 1.161905e-01
R14510 n2_19366_4953 n2_19366_4986 2.095238e-02
R14511 n2_19366_4986 n2_19366_5169 1.161905e-01
R14512 n2_19366_5169 n2_19366_5202 2.095238e-02
R14513 n2_19366_5202 n2_19366_5239 2.349206e-02
R14514 n2_19366_5239 n2_19366_5385 9.269841e-02
R14515 n2_19366_5385 n2_19366_5418 2.095238e-02
R14516 n2_19366_5418 n2_19366_5455 2.349206e-02
R14517 n2_19366_5455 n2_19366_5601 9.269841e-02
R14518 n2_19366_5601 n2_19366_5634 2.095238e-02
R14519 n2_19366_5634 n2_19366_5671 2.349206e-02
R14520 n2_19366_5671 n2_19366_5817 9.269841e-02
R14521 n2_19366_5817 n2_19366_5850 2.095238e-02
R14522 n2_19366_5850 n2_19366_6033 1.161905e-01
R14523 n2_19366_6033 n2_19366_6049 1.015873e-02
R14524 n2_19366_6049 n2_19366_6066 1.079365e-02
R14525 n2_19366_6145 n2_19366_6249 6.603175e-02
R14526 n2_19366_6249 n2_19366_6282 2.095238e-02
R14527 n2_19366_6282 n2_19366_6319 2.349206e-02
R14528 n2_19366_6319 n2_19366_6465 9.269841e-02
R14529 n2_19366_6465 n2_19366_6498 2.095238e-02
R14530 n2_19366_6498 n2_19366_6681 1.161905e-01
R14531 n2_19366_6681 n2_19366_6714 2.095238e-02
R14532 n2_19366_6714 n2_19366_6897 1.161905e-01
R14533 n2_19366_6897 n2_19366_6930 2.095238e-02
R14534 n2_19366_6930 n2_19366_7113 1.161905e-01
R14535 n2_19366_7113 n2_19366_7146 2.095238e-02
R14536 n2_19366_7146 n2_19366_7329 1.161905e-01
R14537 n2_19366_7329 n2_19366_7362 2.095238e-02
R14538 n2_19366_7362 n2_19366_7545 1.161905e-01
R14539 n2_19366_7545 n2_19366_7578 2.095238e-02
R14540 n2_19366_7578 n2_19366_7761 1.161905e-01
R14541 n2_19366_7761 n2_19366_7794 2.095238e-02
R14542 n2_19366_7794 n2_19366_7831 2.349206e-02
R14543 n2_19366_7831 n2_19366_7977 9.269841e-02
R14544 n2_19366_7977 n2_19366_8010 2.095238e-02
R14545 n2_19366_8010 n2_19366_8193 1.161905e-01
R14546 n2_19366_8193 n2_19366_8226 2.095238e-02
R14547 n2_19366_8226 n2_19366_8299 4.634921e-02
R14548 n2_19366_8395 n2_19366_8409 8.888889e-03
R14549 n2_19366_8409 n2_19366_8442 2.095238e-02
R14550 n2_19366_8442 n2_19366_8625 1.161905e-01
R14551 n2_19366_8625 n2_19366_8658 2.095238e-02
R14552 n2_19366_8658 n2_19366_8841 1.161905e-01
R14553 n2_19366_8841 n2_19366_8874 2.095238e-02
R14554 n2_19366_8874 n2_19366_8911 2.349206e-02
R14555 n2_19366_8911 n2_19366_9057 9.269841e-02
R14556 n2_19366_9057 n2_19366_9090 2.095238e-02
R14557 n2_19366_9090 n2_19366_9273 1.161905e-01
R14558 n2_19366_9273 n2_19366_9306 2.095238e-02
R14559 n2_19366_9306 n2_19366_9489 1.161905e-01
R14560 n2_19366_9489 n2_19366_9522 2.095238e-02
R14561 n2_19366_9522 n2_19366_9705 1.161905e-01
R14562 n2_19366_9705 n2_19366_9738 2.095238e-02
R14563 n2_19366_9738 n2_19366_9921 1.161905e-01
R14564 n2_19366_9921 n2_19366_9954 2.095238e-02
R14565 n2_19366_9954 n2_19366_9991 2.349206e-02
R14566 n2_19366_9991 n2_19366_10137 9.269841e-02
R14567 n2_19366_10137 n2_19366_10170 2.095238e-02
R14568 n2_19366_10170 n2_19366_10353 1.161905e-01
R14569 n2_19366_10353 n2_19366_10386 2.095238e-02
R14570 n2_19366_10386 n2_19366_10549 1.034921e-01
R14571 n2_19366_10549 n2_19366_10569 1.269841e-02
R14572 n2_19366_10645 n2_19366_10785 8.888889e-02
R14573 n2_19366_10785 n2_19366_10818 2.095238e-02
R14574 n2_19366_10818 n2_19366_11001 1.161905e-01
R14575 n2_19366_11001 n2_19366_11034 2.095238e-02
R14576 n2_19366_11034 n2_19366_11055 1.333333e-02
R14577 n2_19366_11055 n2_19366_11217 1.028571e-01
R14578 n2_19366_11217 n2_19366_11250 2.095238e-02
R14579 n2_19366_11250 n2_19366_11433 1.161905e-01
R14580 n2_19366_11433 n2_19366_11466 2.095238e-02
R14581 n2_19366_11466 n2_19366_11649 1.161905e-01
R14582 n2_19366_11649 n2_19366_11682 2.095238e-02
R14583 n2_19366_11682 n2_19366_11865 1.161905e-01
R14584 n2_19366_11865 n2_19366_11898 2.095238e-02
R14585 n2_19366_11898 n2_19366_12081 1.161905e-01
R14586 n2_19366_12081 n2_19366_12114 2.095238e-02
R14587 n2_19366_12114 n2_19366_12128 8.888889e-03
R14588 n2_19366_12128 n2_19366_12297 1.073016e-01
R14589 n2_19366_12297 n2_19366_12330 2.095238e-02
R14590 n2_19366_12330 n2_19366_12513 1.161905e-01
R14591 n2_19366_12513 n2_19366_12546 2.095238e-02
R14592 n2_19366_12546 n2_19366_12729 1.161905e-01
R14593 n2_19366_12729 n2_19366_12762 2.095238e-02
R14594 n2_19366_12762 n2_19366_12799 2.349206e-02
R14595 n2_19366_12895 n2_19366_12945 3.174603e-02
R14596 n2_19366_12945 n2_19366_12978 2.095238e-02
R14597 n2_19366_12978 n2_19366_13161 1.161905e-01
R14598 n2_19366_13161 n2_19366_13194 2.095238e-02
R14599 n2_19366_13194 n2_19366_13377 1.161905e-01
R14600 n2_19366_13377 n2_19366_13410 2.095238e-02
R14601 n2_19366_13410 n2_19366_13593 1.161905e-01
R14602 n2_19366_13593 n2_19366_13626 2.095238e-02
R14603 n2_19366_13626 n2_19366_13647 1.333333e-02
R14604 n2_19366_13647 n2_19366_13809 1.028571e-01
R14605 n2_19366_13809 n2_19366_13842 2.095238e-02
R14606 n2_19366_13842 n2_19366_14025 1.161905e-01
R14607 n2_19366_14025 n2_19366_14058 2.095238e-02
R14608 n2_19366_14058 n2_19366_14241 1.161905e-01
R14609 n2_19366_14241 n2_19366_14274 2.095238e-02
R14610 n2_19366_14274 n2_19366_14457 1.161905e-01
R14611 n2_19366_14457 n2_19366_14490 2.095238e-02
R14612 n2_19366_14490 n2_19366_14504 8.888889e-03
R14613 n2_19366_14504 n2_19366_14511 4.444444e-03
R14614 n2_19366_14511 n2_19366_14673 1.028571e-01
R14615 n2_19366_14673 n2_19366_14706 2.095238e-02
R14616 n2_19366_14706 n2_19366_14889 1.161905e-01
R14617 n2_19366_14889 n2_19366_14922 2.095238e-02
R14618 n2_19366_14922 n2_19366_14936 8.888889e-03
R14619 n2_19366_14936 n2_19366_15049 7.174603e-02
R14620 n2_19366_15138 n2_19366_15145 4.444444e-03
R14621 n2_19366_15145 n2_19366_15152 4.444444e-03
R14622 n2_19366_15152 n2_19366_15321 1.073016e-01
R14623 n2_19366_15321 n2_19366_15354 2.095238e-02
R14624 n2_19366_15354 n2_19366_15537 1.161905e-01
R14625 n2_19366_15537 n2_19366_15570 2.095238e-02
R14626 n2_19366_15570 n2_19366_15584 8.888889e-03
R14627 n2_19366_15584 n2_19366_15753 1.073016e-01
R14628 n2_19366_15753 n2_19366_15786 2.095238e-02
R14629 n2_19366_15786 n2_19366_15969 1.161905e-01
R14630 n2_19366_15969 n2_19366_16002 2.095238e-02
R14631 n2_19366_16002 n2_19366_16185 1.161905e-01
R14632 n2_19366_16185 n2_19366_16218 2.095238e-02
R14633 n2_19366_16218 n2_19366_16401 1.161905e-01
R14634 n2_19366_16401 n2_19366_16434 2.095238e-02
R14635 n2_19366_16434 n2_19366_16617 1.161905e-01
R14636 n2_19366_16617 n2_19366_16650 2.095238e-02
R14637 n2_19366_16650 n2_19366_16664 8.888889e-03
R14638 n2_19366_16664 n2_19366_16671 4.444444e-03
R14639 n2_19366_16671 n2_19366_16687 1.015873e-02
R14640 n2_19366_16687 n2_19366_16833 9.269841e-02
R14641 n2_19366_16833 n2_19366_16866 2.095238e-02
R14642 n2_19366_16866 n2_19366_17049 1.161905e-01
R14643 n2_19366_17049 n2_19366_17082 2.095238e-02
R14644 n2_19366_17082 n2_19366_17119 2.349206e-02
R14645 n2_19366_17119 n2_19366_17265 9.269841e-02
R14646 n2_19366_17265 n2_19366_17298 2.095238e-02
R14647 n2_19366_17298 n2_19366_17299 6.349206e-04
R14648 n2_19366_17395 n2_19366_17481 5.460317e-02
R14649 n2_19366_17481 n2_19366_17514 2.095238e-02
R14650 n2_19366_17514 n2_19366_17697 1.161905e-01
R14651 n2_19366_17697 n2_19366_17730 2.095238e-02
R14652 n2_19366_17730 n2_19366_17744 8.888889e-03
R14653 n2_19366_17744 n2_19366_17913 1.073016e-01
R14654 n2_19366_17913 n2_19366_17946 2.095238e-02
R14655 n2_19366_17946 n2_19366_18129 1.161905e-01
R14656 n2_19366_18129 n2_19366_18162 2.095238e-02
R14657 n2_19366_18162 n2_19366_18345 1.161905e-01
R14658 n2_19366_18345 n2_19366_18378 2.095238e-02
R14659 n2_19366_18378 n2_19366_18561 1.161905e-01
R14660 n2_19366_18561 n2_19366_18594 2.095238e-02
R14661 n2_19366_18594 n2_19366_18777 1.161905e-01
R14662 n2_19366_18777 n2_19366_18810 2.095238e-02
R14663 n2_19366_18810 n2_19366_18932 7.746032e-02
R14664 n2_19366_18932 n2_19366_18993 3.873016e-02
R14665 n2_19366_18993 n2_19366_19026 2.095238e-02
R14666 n2_19366_19026 n2_19366_19040 8.888889e-03
R14667 n2_19366_19040 n2_19366_19209 1.073016e-01
R14668 n2_19366_19209 n2_19366_19242 2.095238e-02
R14669 n2_19366_19242 n2_19366_19425 1.161905e-01
R14670 n2_19366_19425 n2_19366_19458 2.095238e-02
R14671 n2_19366_19458 n2_19366_19641 1.161905e-01
R14672 n2_19366_19641 n2_19366_19674 2.095238e-02
R14673 n2_19366_19674 n2_19366_19857 1.161905e-01
R14674 n2_19366_19857 n2_19366_19890 2.095238e-02
R14675 n2_19366_19890 n2_19366_20073 1.161905e-01
R14676 n2_19366_20073 n2_19366_20106 2.095238e-02
R14677 n2_19366_20106 n2_19366_20289 1.161905e-01
R14678 n2_19366_20289 n2_19366_20322 2.095238e-02
R14679 n2_19366_20322 n2_19366_20505 1.161905e-01
R14680 n2_19366_20505 n2_19366_20538 2.095238e-02
R14681 n2_19366_20538 n2_19366_20674 8.634921e-02
R14682 n2_19366_20754 n2_19366_20770 1.015873e-02
R14683 n2_19366_20770 n2_19366_20937 1.060317e-01
R14684 n2_19366_20937 n2_19366_20970 2.095238e-02
R14685 n2_19366_3799 n2_19505_3799 8.825397e-02
R14686 n2_19505_3799 n2_19554_3799 3.111111e-02
R14687 n2_19366_3895 n2_19505_3895 8.825397e-02
R14688 n2_19505_3895 n2_19554_3895 3.111111e-02
R14689 n2_19366_6049 n2_19505_6049 8.825397e-02
R14690 n2_19505_6049 n2_19554_6049 3.111111e-02
R14691 n2_19366_6145 n2_19505_6145 8.825397e-02
R14692 n2_19505_6145 n2_19554_6145 3.111111e-02
R14693 n2_19366_8299 n2_19505_8299 8.825397e-02
R14694 n2_19505_8299 n2_19554_8299 3.111111e-02
R14695 n2_19366_8395 n2_19505_8395 8.825397e-02
R14696 n2_19505_8395 n2_19554_8395 3.111111e-02
R14697 n2_19366_10549 n2_19505_10549 8.825397e-02
R14698 n2_19505_10549 n2_19554_10549 3.111111e-02
R14699 n2_19366_10645 n2_19505_10645 8.825397e-02
R14700 n2_19505_10645 n2_19554_10645 3.111111e-02
R14701 n2_19366_12799 n2_19505_12799 8.825397e-02
R14702 n2_19505_12799 n2_19554_12799 3.111111e-02
R14703 n2_19366_12895 n2_19505_12895 8.825397e-02
R14704 n2_19505_12895 n2_19554_12895 3.111111e-02
R14705 n2_19366_15049 n2_19505_15049 8.825397e-02
R14706 n2_19505_15049 n2_19554_15049 3.111111e-02
R14707 n2_19366_15145 n2_19505_15145 8.825397e-02
R14708 n2_19505_15145 n2_19554_15145 3.111111e-02
R14709 n2_19366_17299 n2_19505_17299 8.825397e-02
R14710 n2_19505_17299 n2_19554_17299 3.111111e-02
R14711 n2_19366_17395 n2_19505_17395 8.825397e-02
R14712 n2_19505_17395 n2_19554_17395 3.111111e-02
R14713 n2_19366_424 n2_19458_424 5.841270e-02
R14714 n2_19458_424 n2_19505_424 2.984127e-02
R14715 n2_19505_424 n2_19554_424 3.111111e-02
R14716 n2_19554_424 n2_19646_424 5.841270e-02
R14717 n2_19366_520 n2_19458_520 5.841270e-02
R14718 n2_19458_520 n2_19505_520 2.984127e-02
R14719 n2_19505_520 n2_19554_520 3.111111e-02
R14720 n2_19554_520 n2_19646_520 5.841270e-02
R14721 n2_19366_20674 n2_19458_20674 5.841270e-02
R14722 n2_19458_20674 n2_19505_20674 2.984127e-02
R14723 n2_19505_20674 n2_19554_20674 3.111111e-02
R14724 n2_19554_20674 n2_19646_20674 5.841270e-02
R14725 n2_19366_20770 n2_19458_20770 5.841270e-02
R14726 n2_19458_20770 n2_19505_20770 2.984127e-02
R14727 n2_19505_20770 n2_19554_20770 3.111111e-02
R14728 n2_19554_20770 n2_19646_20770 5.841270e-02
R14729 n2_19458_201 n2_19458_234 2.095238e-02
R14730 n2_19458_234 n2_19458_417 1.161905e-01
R14731 n2_19458_417 n2_19458_424 4.444444e-03
R14732 n2_19458_424 n2_19458_450 1.650794e-02
R14733 n2_19458_450 n2_19458_520 4.444444e-02
R14734 n2_19458_520 n2_19458_633 7.174603e-02
R14735 n2_19458_633 n2_19458_666 2.095238e-02
R14736 n2_19458_666 n2_19458_849 1.161905e-01
R14737 n2_19458_849 n2_19458_882 2.095238e-02
R14738 n2_19458_882 n2_19458_1065 1.161905e-01
R14739 n2_19458_1065 n2_19458_1098 2.095238e-02
R14740 n2_19458_1098 n2_19458_1281 1.161905e-01
R14741 n2_19458_1281 n2_19458_1314 2.095238e-02
R14742 n2_19458_1314 n2_19458_1497 1.161905e-01
R14743 n2_19458_19857 n2_19458_19890 2.095238e-02
R14744 n2_19458_19890 n2_19458_20073 1.161905e-01
R14745 n2_19458_20073 n2_19458_20106 2.095238e-02
R14746 n2_19458_20106 n2_19458_20289 1.161905e-01
R14747 n2_19458_20289 n2_19458_20322 2.095238e-02
R14748 n2_19458_20322 n2_19458_20505 1.161905e-01
R14749 n2_19458_20505 n2_19458_20538 2.095238e-02
R14750 n2_19458_20538 n2_19458_20674 8.634921e-02
R14751 n2_19458_20674 n2_19458_20721 2.984127e-02
R14752 n2_19458_20721 n2_19458_20754 2.095238e-02
R14753 n2_19458_20754 n2_19458_20770 1.015873e-02
R14754 n2_19458_20770 n2_19458_20937 1.060317e-01
R14755 n2_19458_20937 n2_19458_20970 2.095238e-02
R14756 n2_19554_201 n2_19554_234 2.095238e-02
R14757 n2_19554_234 n2_19554_417 1.161905e-01
R14758 n2_19554_417 n2_19554_424 4.444444e-03
R14759 n2_19554_424 n2_19554_450 1.650794e-02
R14760 n2_19554_450 n2_19554_520 4.444444e-02
R14761 n2_19554_520 n2_19554_633 7.174603e-02
R14762 n2_19554_633 n2_19554_666 2.095238e-02
R14763 n2_19554_666 n2_19554_849 1.161905e-01
R14764 n2_19554_849 n2_19554_882 2.095238e-02
R14765 n2_19554_882 n2_19554_1065 1.161905e-01
R14766 n2_19554_1065 n2_19554_1098 2.095238e-02
R14767 n2_19554_1098 n2_19554_1281 1.161905e-01
R14768 n2_19554_1281 n2_19554_1314 2.095238e-02
R14769 n2_19554_1314 n2_19554_1497 1.161905e-01
R14770 n2_19554_1713 n2_19554_1746 2.095238e-02
R14771 n2_19554_1746 n2_19554_1929 1.161905e-01
R14772 n2_19554_1929 n2_19554_1962 2.095238e-02
R14773 n2_19554_1962 n2_19554_1976 8.888889e-03
R14774 n2_19554_1976 n2_19554_1999 1.460317e-02
R14775 n2_19554_1999 n2_19554_2145 9.269841e-02
R14776 n2_19554_2145 n2_19554_2178 2.095238e-02
R14777 n2_19554_2178 n2_19554_2361 1.161905e-01
R14778 n2_19554_2361 n2_19554_2394 2.095238e-02
R14779 n2_19554_2394 n2_19554_2577 1.161905e-01
R14780 n2_19554_2577 n2_19554_2610 2.095238e-02
R14781 n2_19554_2826 n2_19554_3009 1.161905e-01
R14782 n2_19554_3009 n2_19554_3042 2.095238e-02
R14783 n2_19554_3042 n2_19554_3225 1.161905e-01
R14784 n2_19554_3225 n2_19554_3258 2.095238e-02
R14785 n2_19554_3258 n2_19554_3295 2.349206e-02
R14786 n2_19554_3295 n2_19554_3441 9.269841e-02
R14787 n2_19554_3441 n2_19554_3474 2.095238e-02
R14788 n2_19554_3474 n2_19554_3657 1.161905e-01
R14789 n2_19554_3657 n2_19554_3690 2.095238e-02
R14790 n2_19554_3690 n2_19554_3799 6.920635e-02
R14791 n2_19554_3799 n2_19554_3873 4.698413e-02
R14792 n2_19554_3873 n2_19554_3895 1.396825e-02
R14793 n2_19554_3895 n2_19554_3906 6.984127e-03
R14794 n2_19554_3906 n2_19554_4089 1.161905e-01
R14795 n2_19554_4089 n2_19554_4122 2.095238e-02
R14796 n2_19554_4122 n2_19554_4305 1.161905e-01
R14797 n2_19554_4305 n2_19554_4338 2.095238e-02
R14798 n2_19554_4338 n2_19554_4375 2.349206e-02
R14799 n2_19554_4375 n2_19554_4521 9.269841e-02
R14800 n2_19554_4521 n2_19554_4554 2.095238e-02
R14801 n2_19554_4554 n2_19554_4737 1.161905e-01
R14802 n2_19554_4737 n2_19554_4770 2.095238e-02
R14803 n2_19554_5169 n2_19554_5202 2.095238e-02
R14804 n2_19554_5202 n2_19554_5239 2.349206e-02
R14805 n2_19554_5239 n2_19554_5385 9.269841e-02
R14806 n2_19554_5385 n2_19554_5418 2.095238e-02
R14807 n2_19554_5418 n2_19554_5455 2.349206e-02
R14808 n2_19554_5455 n2_19554_5601 9.269841e-02
R14809 n2_19554_5601 n2_19554_5634 2.095238e-02
R14810 n2_19554_5634 n2_19554_5671 2.349206e-02
R14811 n2_19554_5671 n2_19554_5817 9.269841e-02
R14812 n2_19554_5817 n2_19554_5850 2.095238e-02
R14813 n2_19554_5850 n2_19554_6033 1.161905e-01
R14814 n2_19554_6033 n2_19554_6049 1.015873e-02
R14815 n2_19554_6049 n2_19554_6066 1.079365e-02
R14816 n2_19554_6066 n2_19554_6145 5.015873e-02
R14817 n2_19554_6145 n2_19554_6249 6.603175e-02
R14818 n2_19554_6249 n2_19554_6282 2.095238e-02
R14819 n2_19554_6282 n2_19554_6319 2.349206e-02
R14820 n2_19554_6319 n2_19554_6465 9.269841e-02
R14821 n2_19554_6465 n2_19554_6498 2.095238e-02
R14822 n2_19554_6498 n2_19554_6681 1.161905e-01
R14823 n2_19554_6681 n2_19554_6714 2.095238e-02
R14824 n2_19554_6714 n2_19554_6897 1.161905e-01
R14825 n2_19554_6897 n2_19554_6930 2.095238e-02
R14826 n2_19554_6930 n2_19554_7113 1.161905e-01
R14827 n2_19554_7329 n2_19554_7362 2.095238e-02
R14828 n2_19554_7362 n2_19554_7545 1.161905e-01
R14829 n2_19554_7545 n2_19554_7578 2.095238e-02
R14830 n2_19554_7578 n2_19554_7761 1.161905e-01
R14831 n2_19554_7761 n2_19554_7794 2.095238e-02
R14832 n2_19554_7794 n2_19554_7831 2.349206e-02
R14833 n2_19554_7831 n2_19554_7977 9.269841e-02
R14834 n2_19554_7977 n2_19554_8010 2.095238e-02
R14835 n2_19554_8010 n2_19554_8193 1.161905e-01
R14836 n2_19554_8193 n2_19554_8226 2.095238e-02
R14837 n2_19554_8226 n2_19554_8299 4.634921e-02
R14838 n2_19554_8299 n2_19554_8395 6.095238e-02
R14839 n2_19554_8395 n2_19554_8409 8.888889e-03
R14840 n2_19554_8409 n2_19554_8442 2.095238e-02
R14841 n2_19554_8442 n2_19554_8625 1.161905e-01
R14842 n2_19554_8625 n2_19554_8658 2.095238e-02
R14843 n2_19554_8658 n2_19554_8841 1.161905e-01
R14844 n2_19554_8841 n2_19554_8874 2.095238e-02
R14845 n2_19554_8874 n2_19554_8911 2.349206e-02
R14846 n2_19554_8911 n2_19554_9057 9.269841e-02
R14847 n2_19554_9057 n2_19554_9090 2.095238e-02
R14848 n2_19554_9090 n2_19554_9273 1.161905e-01
R14849 n2_19554_9273 n2_19554_9306 2.095238e-02
R14850 n2_19554_9705 n2_19554_9738 2.095238e-02
R14851 n2_19554_9738 n2_19554_9921 1.161905e-01
R14852 n2_19554_9921 n2_19554_9954 2.095238e-02
R14853 n2_19554_9954 n2_19554_9991 2.349206e-02
R14854 n2_19554_9991 n2_19554_10137 9.269841e-02
R14855 n2_19554_10137 n2_19554_10170 2.095238e-02
R14856 n2_19554_10170 n2_19554_10353 1.161905e-01
R14857 n2_19554_10353 n2_19554_10386 2.095238e-02
R14858 n2_19554_10386 n2_19554_10549 1.034921e-01
R14859 n2_19554_10549 n2_19554_10569 1.269841e-02
R14860 n2_19554_10569 n2_19554_10602 2.095238e-02
R14861 n2_19554_10602 n2_19554_10645 2.730159e-02
R14862 n2_19554_10645 n2_19554_10785 8.888889e-02
R14863 n2_19554_10785 n2_19554_10818 2.095238e-02
R14864 n2_19554_10818 n2_19554_11001 1.161905e-01
R14865 n2_19554_11001 n2_19554_11034 2.095238e-02
R14866 n2_19554_11034 n2_19554_11055 1.333333e-02
R14867 n2_19554_11055 n2_19554_11217 1.028571e-01
R14868 n2_19554_11217 n2_19554_11250 2.095238e-02
R14869 n2_19554_11250 n2_19554_11433 1.161905e-01
R14870 n2_19554_11433 n2_19554_11466 2.095238e-02
R14871 n2_19554_11865 n2_19554_11898 2.095238e-02
R14872 n2_19554_11898 n2_19554_12081 1.161905e-01
R14873 n2_19554_12081 n2_19554_12114 2.095238e-02
R14874 n2_19554_12114 n2_19554_12128 8.888889e-03
R14875 n2_19554_12128 n2_19554_12297 1.073016e-01
R14876 n2_19554_12297 n2_19554_12330 2.095238e-02
R14877 n2_19554_12330 n2_19554_12513 1.161905e-01
R14878 n2_19554_12513 n2_19554_12546 2.095238e-02
R14879 n2_19554_12546 n2_19554_12729 1.161905e-01
R14880 n2_19554_12729 n2_19554_12762 2.095238e-02
R14881 n2_19554_12762 n2_19554_12799 2.349206e-02
R14882 n2_19554_12799 n2_19554_12895 6.095238e-02
R14883 n2_19554_12895 n2_19554_12945 3.174603e-02
R14884 n2_19554_12945 n2_19554_12978 2.095238e-02
R14885 n2_19554_12978 n2_19554_13161 1.161905e-01
R14886 n2_19554_13161 n2_19554_13194 2.095238e-02
R14887 n2_19554_13194 n2_19554_13377 1.161905e-01
R14888 n2_19554_13377 n2_19554_13410 2.095238e-02
R14889 n2_19554_13410 n2_19554_13593 1.161905e-01
R14890 n2_19554_13593 n2_19554_13626 2.095238e-02
R14891 n2_19554_13626 n2_19554_13647 1.333333e-02
R14892 n2_19554_13647 n2_19554_13809 1.028571e-01
R14893 n2_19554_13809 n2_19554_13842 2.095238e-02
R14894 n2_19554_14241 n2_19554_14274 2.095238e-02
R14895 n2_19554_14274 n2_19554_14457 1.161905e-01
R14896 n2_19554_14457 n2_19554_14490 2.095238e-02
R14897 n2_19554_14490 n2_19554_14504 8.888889e-03
R14898 n2_19554_14504 n2_19554_14511 4.444444e-03
R14899 n2_19554_14511 n2_19554_14673 1.028571e-01
R14900 n2_19554_14673 n2_19554_14706 2.095238e-02
R14901 n2_19554_14706 n2_19554_14889 1.161905e-01
R14902 n2_19554_14889 n2_19554_14922 2.095238e-02
R14903 n2_19554_14922 n2_19554_14936 8.888889e-03
R14904 n2_19554_14936 n2_19554_15049 7.174603e-02
R14905 n2_19554_15049 n2_19554_15105 3.555556e-02
R14906 n2_19554_15105 n2_19554_15138 2.095238e-02
R14907 n2_19554_15138 n2_19554_15145 4.444444e-03
R14908 n2_19554_15145 n2_19554_15152 4.444444e-03
R14909 n2_19554_15152 n2_19554_15321 1.073016e-01
R14910 n2_19554_15321 n2_19554_15354 2.095238e-02
R14911 n2_19554_15354 n2_19554_15537 1.161905e-01
R14912 n2_19554_15537 n2_19554_15570 2.095238e-02
R14913 n2_19554_15570 n2_19554_15584 8.888889e-03
R14914 n2_19554_15584 n2_19554_15753 1.073016e-01
R14915 n2_19554_15753 n2_19554_15786 2.095238e-02
R14916 n2_19554_15786 n2_19554_15969 1.161905e-01
R14917 n2_19554_15969 n2_19554_16002 2.095238e-02
R14918 n2_19554_16401 n2_19554_16434 2.095238e-02
R14919 n2_19554_16434 n2_19554_16617 1.161905e-01
R14920 n2_19554_16617 n2_19554_16650 2.095238e-02
R14921 n2_19554_16650 n2_19554_16664 8.888889e-03
R14922 n2_19554_16664 n2_19554_16671 4.444444e-03
R14923 n2_19554_16671 n2_19554_16687 1.015873e-02
R14924 n2_19554_16687 n2_19554_16833 9.269841e-02
R14925 n2_19554_16833 n2_19554_16866 2.095238e-02
R14926 n2_19554_16866 n2_19554_17049 1.161905e-01
R14927 n2_19554_17049 n2_19554_17082 2.095238e-02
R14928 n2_19554_17082 n2_19554_17119 2.349206e-02
R14929 n2_19554_17119 n2_19554_17265 9.269841e-02
R14930 n2_19554_17265 n2_19554_17298 2.095238e-02
R14931 n2_19554_17298 n2_19554_17299 6.349206e-04
R14932 n2_19554_17299 n2_19554_17395 6.095238e-02
R14933 n2_19554_17395 n2_19554_17481 5.460317e-02
R14934 n2_19554_17481 n2_19554_17514 2.095238e-02
R14935 n2_19554_17514 n2_19554_17697 1.161905e-01
R14936 n2_19554_17697 n2_19554_17730 2.095238e-02
R14937 n2_19554_17730 n2_19554_17744 8.888889e-03
R14938 n2_19554_17744 n2_19554_17913 1.073016e-01
R14939 n2_19554_17913 n2_19554_17946 2.095238e-02
R14940 n2_19554_17946 n2_19554_18129 1.161905e-01
R14941 n2_19554_18129 n2_19554_18162 2.095238e-02
R14942 n2_19554_18162 n2_19554_18345 1.161905e-01
R14943 n2_19554_18594 n2_19554_18777 1.161905e-01
R14944 n2_19554_18777 n2_19554_18810 2.095238e-02
R14945 n2_19554_18810 n2_19554_18932 7.746032e-02
R14946 n2_19554_18932 n2_19554_18993 3.873016e-02
R14947 n2_19554_18993 n2_19554_19026 2.095238e-02
R14948 n2_19554_19026 n2_19554_19040 8.888889e-03
R14949 n2_19554_19040 n2_19554_19209 1.073016e-01
R14950 n2_19554_19209 n2_19554_19242 2.095238e-02
R14951 n2_19554_19242 n2_19554_19425 1.161905e-01
R14952 n2_19554_19425 n2_19554_19458 2.095238e-02
R14953 n2_19554_19857 n2_19554_19890 2.095238e-02
R14954 n2_19554_19890 n2_19554_20073 1.161905e-01
R14955 n2_19554_20073 n2_19554_20106 2.095238e-02
R14956 n2_19554_20106 n2_19554_20289 1.161905e-01
R14957 n2_19554_20289 n2_19554_20322 2.095238e-02
R14958 n2_19554_20322 n2_19554_20505 1.161905e-01
R14959 n2_19554_20505 n2_19554_20538 2.095238e-02
R14960 n2_19554_20538 n2_19554_20674 8.634921e-02
R14961 n2_19554_20674 n2_19554_20721 2.984127e-02
R14962 n2_19554_20721 n2_19554_20754 2.095238e-02
R14963 n2_19554_20754 n2_19554_20770 1.015873e-02
R14964 n2_19554_20770 n2_19554_20937 1.060317e-01
R14965 n2_19554_20937 n2_19554_20970 2.095238e-02
R14966 n2_19646_201 n2_19646_234 2.095238e-02
R14967 n2_19646_234 n2_19646_417 1.161905e-01
R14968 n2_19646_417 n2_19646_424 4.444444e-03
R14969 n2_19646_424 n2_19646_450 1.650794e-02
R14970 n2_19646_520 n2_19646_633 7.174603e-02
R14971 n2_19646_633 n2_19646_666 2.095238e-02
R14972 n2_19646_666 n2_19646_849 1.161905e-01
R14973 n2_19646_849 n2_19646_882 2.095238e-02
R14974 n2_19646_882 n2_19646_1065 1.161905e-01
R14975 n2_19646_1065 n2_19646_1098 2.095238e-02
R14976 n2_19646_1098 n2_19646_1281 1.161905e-01
R14977 n2_19646_1281 n2_19646_1314 2.095238e-02
R14978 n2_19646_1314 n2_19646_1497 1.161905e-01
R14979 n2_19646_1497 n2_19646_1530 2.095238e-02
R14980 n2_19646_19641 n2_19646_19674 2.095238e-02
R14981 n2_19646_19674 n2_19646_19857 1.161905e-01
R14982 n2_19646_19857 n2_19646_19890 2.095238e-02
R14983 n2_19646_19890 n2_19646_20073 1.161905e-01
R14984 n2_19646_20073 n2_19646_20106 2.095238e-02
R14985 n2_19646_20106 n2_19646_20289 1.161905e-01
R14986 n2_19646_20289 n2_19646_20322 2.095238e-02
R14987 n2_19646_20322 n2_19646_20505 1.161905e-01
R14988 n2_19646_20505 n2_19646_20538 2.095238e-02
R14989 n2_19646_20538 n2_19646_20674 8.634921e-02
R14990 n2_19646_20754 n2_19646_20770 1.015873e-02
R14991 n2_19646_20770 n2_19646_20937 1.060317e-01
R14992 n2_19646_20937 n2_19646_20970 2.095238e-02
R14993 n2_20491_633 n2_20491_666 2.095238e-02
R14994 n2_20491_666 n2_20491_849 1.161905e-01
R14995 n2_20491_849 n2_20491_882 2.095238e-02
R14996 n2_20491_882 n2_20491_1065 1.161905e-01
R14997 n2_20491_1065 n2_20491_1098 2.095238e-02
R14998 n2_20491_1098 n2_20491_1281 1.161905e-01
R14999 n2_20491_1281 n2_20491_1314 2.095238e-02
R15000 n2_20491_1314 n2_20491_1497 1.161905e-01
R15001 n2_20491_1497 n2_20491_1530 2.095238e-02
R15002 n2_20491_1530 n2_20491_1549 1.206349e-02
R15003 n2_20491_1645 n2_20491_1713 4.317460e-02
R15004 n2_20491_1713 n2_20491_1746 2.095238e-02
R15005 n2_20491_1746 n2_20491_1929 1.161905e-01
R15006 n2_20491_1929 n2_20491_1962 2.095238e-02
R15007 n2_20491_1962 n2_20491_1976 8.888889e-03
R15008 n2_20491_1976 n2_20491_2145 1.073016e-01
R15009 n2_20491_2145 n2_20491_2178 2.095238e-02
R15010 n2_20491_2178 n2_20491_2361 1.161905e-01
R15011 n2_20491_2361 n2_20491_2394 2.095238e-02
R15012 n2_20491_2394 n2_20491_2577 1.161905e-01
R15013 n2_20491_2577 n2_20491_2610 2.095238e-02
R15014 n2_20491_2610 n2_20491_2793 1.161905e-01
R15015 n2_20491_2793 n2_20491_2826 2.095238e-02
R15016 n2_20491_2826 n2_20491_3009 1.161905e-01
R15017 n2_20491_3009 n2_20491_3042 2.095238e-02
R15018 n2_20491_3042 n2_20491_3225 1.161905e-01
R15019 n2_20491_3225 n2_20491_3258 2.095238e-02
R15020 n2_20491_3258 n2_20491_3441 1.161905e-01
R15021 n2_20491_3441 n2_20491_3474 2.095238e-02
R15022 n2_20491_3474 n2_20491_3657 1.161905e-01
R15023 n2_20491_3657 n2_20491_3690 2.095238e-02
R15024 n2_20491_3690 n2_20491_3799 6.920635e-02
R15025 n2_20491_3873 n2_20491_3895 1.396825e-02
R15026 n2_20491_3895 n2_20491_3906 6.984127e-03
R15027 n2_20491_3906 n2_20491_4089 1.161905e-01
R15028 n2_20491_4089 n2_20491_4122 2.095238e-02
R15029 n2_20491_4122 n2_20491_4305 1.161905e-01
R15030 n2_20491_4305 n2_20491_4338 2.095238e-02
R15031 n2_20491_4338 n2_20491_4521 1.161905e-01
R15032 n2_20491_4521 n2_20491_4554 2.095238e-02
R15033 n2_20491_4554 n2_20491_4737 1.161905e-01
R15034 n2_20491_4737 n2_20491_4770 2.095238e-02
R15035 n2_20491_4770 n2_20491_4953 1.161905e-01
R15036 n2_20491_4953 n2_20491_4986 2.095238e-02
R15037 n2_20491_4986 n2_20491_5169 1.161905e-01
R15038 n2_20491_5169 n2_20491_5202 2.095238e-02
R15039 n2_20491_5202 n2_20491_5385 1.161905e-01
R15040 n2_20491_5385 n2_20491_5418 2.095238e-02
R15041 n2_20491_5418 n2_20491_5601 1.161905e-01
R15042 n2_20491_5601 n2_20491_5634 2.095238e-02
R15043 n2_20491_5634 n2_20491_5671 2.349206e-02
R15044 n2_20491_5671 n2_20491_5817 9.269841e-02
R15045 n2_20491_5817 n2_20491_5850 2.095238e-02
R15046 n2_20491_5850 n2_20491_6033 1.161905e-01
R15047 n2_20491_6033 n2_20491_6049 1.015873e-02
R15048 n2_20491_6049 n2_20491_6066 1.079365e-02
R15049 n2_20491_6145 n2_20491_6249 6.603175e-02
R15050 n2_20491_6249 n2_20491_6282 2.095238e-02
R15051 n2_20491_6282 n2_20491_6319 2.349206e-02
R15052 n2_20491_6319 n2_20491_6465 9.269841e-02
R15053 n2_20491_6465 n2_20491_6498 2.095238e-02
R15054 n2_20491_6498 n2_20491_6681 1.161905e-01
R15055 n2_20491_6681 n2_20491_6714 2.095238e-02
R15056 n2_20491_6714 n2_20491_6897 1.161905e-01
R15057 n2_20491_6897 n2_20491_6930 2.095238e-02
R15058 n2_20491_6930 n2_20491_7113 1.161905e-01
R15059 n2_20491_7113 n2_20491_7146 2.095238e-02
R15060 n2_20491_7146 n2_20491_7329 1.161905e-01
R15061 n2_20491_7329 n2_20491_7362 2.095238e-02
R15062 n2_20491_7362 n2_20491_7545 1.161905e-01
R15063 n2_20491_7545 n2_20491_7578 2.095238e-02
R15064 n2_20491_7578 n2_20491_7761 1.161905e-01
R15065 n2_20491_7761 n2_20491_7794 2.095238e-02
R15066 n2_20491_7794 n2_20491_7977 1.161905e-01
R15067 n2_20491_7977 n2_20491_8010 2.095238e-02
R15068 n2_20491_8010 n2_20491_8193 1.161905e-01
R15069 n2_20491_8193 n2_20491_8226 2.095238e-02
R15070 n2_20491_8226 n2_20491_8299 4.634921e-02
R15071 n2_20491_8395 n2_20491_8409 8.888889e-03
R15072 n2_20491_8409 n2_20491_8442 2.095238e-02
R15073 n2_20491_8442 n2_20491_8625 1.161905e-01
R15074 n2_20491_8625 n2_20491_8658 2.095238e-02
R15075 n2_20491_8658 n2_20491_8841 1.161905e-01
R15076 n2_20491_8841 n2_20491_8874 2.095238e-02
R15077 n2_20491_8874 n2_20491_9057 1.161905e-01
R15078 n2_20491_9057 n2_20491_9090 2.095238e-02
R15079 n2_20491_9090 n2_20491_9213 7.809524e-02
R15080 n2_20491_9213 n2_20491_10549 8.482540e-01
R15081 n2_20491_10645 n2_20491_11956 8.323810e-01
R15082 n2_20491_11956 n2_20491_12081 7.936508e-02
R15083 n2_20491_12081 n2_20491_12114 2.095238e-02
R15084 n2_20491_12114 n2_20491_12297 1.161905e-01
R15085 n2_20491_12297 n2_20491_12330 2.095238e-02
R15086 n2_20491_12330 n2_20491_12513 1.161905e-01
R15087 n2_20491_12513 n2_20491_12546 2.095238e-02
R15088 n2_20491_12546 n2_20491_12729 1.161905e-01
R15089 n2_20491_12729 n2_20491_12762 2.095238e-02
R15090 n2_20491_12762 n2_20491_12799 2.349206e-02
R15091 n2_20491_12895 n2_20491_12945 3.174603e-02
R15092 n2_20491_12945 n2_20491_12978 2.095238e-02
R15093 n2_20491_12978 n2_20491_13161 1.161905e-01
R15094 n2_20491_13161 n2_20491_13194 2.095238e-02
R15095 n2_20491_13194 n2_20491_13377 1.161905e-01
R15096 n2_20491_13377 n2_20491_13410 2.095238e-02
R15097 n2_20491_13410 n2_20491_13593 1.161905e-01
R15098 n2_20491_13593 n2_20491_13626 2.095238e-02
R15099 n2_20491_13626 n2_20491_13809 1.161905e-01
R15100 n2_20491_13809 n2_20491_13842 2.095238e-02
R15101 n2_20491_13842 n2_20491_14025 1.161905e-01
R15102 n2_20491_14025 n2_20491_14058 2.095238e-02
R15103 n2_20491_14058 n2_20491_14241 1.161905e-01
R15104 n2_20491_14241 n2_20491_14274 2.095238e-02
R15105 n2_20491_14274 n2_20491_14457 1.161905e-01
R15106 n2_20491_14457 n2_20491_14490 2.095238e-02
R15107 n2_20491_14490 n2_20491_14673 1.161905e-01
R15108 n2_20491_14673 n2_20491_14706 2.095238e-02
R15109 n2_20491_14706 n2_20491_14889 1.161905e-01
R15110 n2_20491_14889 n2_20491_14922 2.095238e-02
R15111 n2_20491_14922 n2_20491_14936 8.888889e-03
R15112 n2_20491_14936 n2_20491_15049 7.174603e-02
R15113 n2_20491_15138 n2_20491_15145 4.444444e-03
R15114 n2_20491_15145 n2_20491_15152 4.444444e-03
R15115 n2_20491_15152 n2_20491_15321 1.073016e-01
R15116 n2_20491_15321 n2_20491_15354 2.095238e-02
R15117 n2_20491_15354 n2_20491_15537 1.161905e-01
R15118 n2_20491_15537 n2_20491_15570 2.095238e-02
R15119 n2_20491_15570 n2_20491_15753 1.161905e-01
R15120 n2_20491_15753 n2_20491_15786 2.095238e-02
R15121 n2_20491_15786 n2_20491_15969 1.161905e-01
R15122 n2_20491_15969 n2_20491_16002 2.095238e-02
R15123 n2_20491_16002 n2_20491_16185 1.161905e-01
R15124 n2_20491_16185 n2_20491_16218 2.095238e-02
R15125 n2_20491_16218 n2_20491_16401 1.161905e-01
R15126 n2_20491_16401 n2_20491_16434 2.095238e-02
R15127 n2_20491_16434 n2_20491_16617 1.161905e-01
R15128 n2_20491_16617 n2_20491_16650 2.095238e-02
R15129 n2_20491_16650 n2_20491_16687 2.349206e-02
R15130 n2_20491_16687 n2_20491_16833 9.269841e-02
R15131 n2_20491_16833 n2_20491_16866 2.095238e-02
R15132 n2_20491_16866 n2_20491_17049 1.161905e-01
R15133 n2_20491_17049 n2_20491_17082 2.095238e-02
R15134 n2_20491_17082 n2_20491_17265 1.161905e-01
R15135 n2_20491_17265 n2_20491_17298 2.095238e-02
R15136 n2_20491_17298 n2_20491_17299 6.349206e-04
R15137 n2_20491_17395 n2_20491_17481 5.460317e-02
R15138 n2_20491_17481 n2_20491_17514 2.095238e-02
R15139 n2_20491_17514 n2_20491_17697 1.161905e-01
R15140 n2_20491_17697 n2_20491_17730 2.095238e-02
R15141 n2_20491_17730 n2_20491_17913 1.161905e-01
R15142 n2_20491_17913 n2_20491_17946 2.095238e-02
R15143 n2_20491_17946 n2_20491_18129 1.161905e-01
R15144 n2_20491_18129 n2_20491_18162 2.095238e-02
R15145 n2_20491_18162 n2_20491_18345 1.161905e-01
R15146 n2_20491_18345 n2_20491_18378 2.095238e-02
R15147 n2_20491_18378 n2_20491_18561 1.161905e-01
R15148 n2_20491_18561 n2_20491_18594 2.095238e-02
R15149 n2_20491_18594 n2_20491_18777 1.161905e-01
R15150 n2_20491_18777 n2_20491_18810 2.095238e-02
R15151 n2_20491_18810 n2_20491_18993 1.161905e-01
R15152 n2_20491_18993 n2_20491_19026 2.095238e-02
R15153 n2_20491_19026 n2_20491_19040 8.888889e-03
R15154 n2_20491_19040 n2_20491_19209 1.073016e-01
R15155 n2_20491_19209 n2_20491_19242 2.095238e-02
R15156 n2_20491_19242 n2_20491_19425 1.161905e-01
R15157 n2_20491_19425 n2_20491_19458 2.095238e-02
R15158 n2_20491_19458 n2_20491_19549 5.777778e-02
R15159 n2_20491_19641 n2_20491_19645 2.539683e-03
R15160 n2_20491_19645 n2_20491_19674 1.841270e-02
R15161 n2_20491_19674 n2_20491_19857 1.161905e-01
R15162 n2_20491_19857 n2_20491_19890 2.095238e-02
R15163 n2_20491_19890 n2_20491_20073 1.161905e-01
R15164 n2_20491_20073 n2_20491_20106 2.095238e-02
R15165 n2_20491_20106 n2_20491_20289 1.161905e-01
R15166 n2_20491_20289 n2_20491_20322 2.095238e-02
R15167 n2_20491_20322 n2_20491_20505 1.161905e-01
R15168 n2_20491_20505 n2_20491_20538 2.095238e-02
R15169 n2_20491_1549 n2_20630_1549 8.825397e-02
R15170 n2_20630_1549 n2_20679_1549 3.111111e-02
R15171 n2_20491_1645 n2_20630_1645 8.825397e-02
R15172 n2_20630_1645 n2_20679_1645 3.111111e-02
R15173 n2_20491_3799 n2_20630_3799 8.825397e-02
R15174 n2_20630_3799 n2_20679_3799 3.111111e-02
R15175 n2_20491_3895 n2_20630_3895 8.825397e-02
R15176 n2_20630_3895 n2_20679_3895 3.111111e-02
R15177 n2_20491_6049 n2_20630_6049 8.825397e-02
R15178 n2_20630_6049 n2_20679_6049 3.111111e-02
R15179 n2_20491_6145 n2_20630_6145 8.825397e-02
R15180 n2_20630_6145 n2_20679_6145 3.111111e-02
R15181 n2_20491_8299 n2_20630_8299 8.825397e-02
R15182 n2_20630_8299 n2_20679_8299 3.111111e-02
R15183 n2_20491_8395 n2_20630_8395 8.825397e-02
R15184 n2_20630_8395 n2_20679_8395 3.111111e-02
R15185 n2_20491_10549 n2_20630_10549 8.825397e-02
R15186 n2_20630_10549 n2_20679_10549 3.111111e-02
R15187 n2_20491_10645 n2_20630_10645 8.825397e-02
R15188 n2_20630_10645 n2_20679_10645 3.111111e-02
R15189 n2_20491_12799 n2_20630_12799 8.825397e-02
R15190 n2_20630_12799 n2_20679_12799 3.111111e-02
R15191 n2_20491_12895 n2_20630_12895 8.825397e-02
R15192 n2_20630_12895 n2_20679_12895 3.111111e-02
R15193 n2_20491_15049 n2_20630_15049 8.825397e-02
R15194 n2_20630_15049 n2_20679_15049 3.111111e-02
R15195 n2_20491_15145 n2_20630_15145 8.825397e-02
R15196 n2_20630_15145 n2_20679_15145 3.111111e-02
R15197 n2_20491_17299 n2_20630_17299 8.825397e-02
R15198 n2_20630_17299 n2_20679_17299 3.111111e-02
R15199 n2_20491_17395 n2_20630_17395 8.825397e-02
R15200 n2_20630_17395 n2_20679_17395 3.111111e-02
R15201 n2_20491_19549 n2_20630_19549 8.825397e-02
R15202 n2_20630_19549 n2_20679_19549 3.111111e-02
R15203 n2_20491_19645 n2_20630_19645 8.825397e-02
R15204 n2_20630_19645 n2_20679_19645 3.111111e-02
R15205 n2_20679_633 n2_20679_666 2.095238e-02
R15206 n2_20679_666 n2_20679_849 1.161905e-01
R15207 n2_20679_849 n2_20679_882 2.095238e-02
R15208 n2_20679_882 n2_20679_1065 1.161905e-01
R15209 n2_20679_1065 n2_20679_1098 2.095238e-02
R15210 n2_20679_1098 n2_20679_1281 1.161905e-01
R15211 n2_20679_1281 n2_20679_1314 2.095238e-02
R15212 n2_20679_1314 n2_20679_1497 1.161905e-01
R15213 n2_20679_1497 n2_20679_1530 2.095238e-02
R15214 n2_20679_1530 n2_20679_1549 1.206349e-02
R15215 n2_20679_1549 n2_20679_1645 6.095238e-02
R15216 n2_20679_1645 n2_20679_1713 4.317460e-02
R15217 n2_20679_1713 n2_20679_1746 2.095238e-02
R15218 n2_20679_1746 n2_20679_1929 1.161905e-01
R15219 n2_20679_1929 n2_20679_1962 2.095238e-02
R15220 n2_20679_1962 n2_20679_1976 8.888889e-03
R15221 n2_20679_1976 n2_20679_2145 1.073016e-01
R15222 n2_20679_2145 n2_20679_2178 2.095238e-02
R15223 n2_20679_2178 n2_20679_2361 1.161905e-01
R15224 n2_20679_2361 n2_20679_2394 2.095238e-02
R15225 n2_20679_2394 n2_20679_2577 1.161905e-01
R15226 n2_20679_2577 n2_20679_2610 2.095238e-02
R15227 n2_20679_2826 n2_20679_3009 1.161905e-01
R15228 n2_20679_3009 n2_20679_3042 2.095238e-02
R15229 n2_20679_3042 n2_20679_3225 1.161905e-01
R15230 n2_20679_3225 n2_20679_3258 2.095238e-02
R15231 n2_20679_3258 n2_20679_3441 1.161905e-01
R15232 n2_20679_3441 n2_20679_3474 2.095238e-02
R15233 n2_20679_3474 n2_20679_3657 1.161905e-01
R15234 n2_20679_3657 n2_20679_3690 2.095238e-02
R15235 n2_20679_3690 n2_20679_3799 6.920635e-02
R15236 n2_20679_3799 n2_20679_3873 4.698413e-02
R15237 n2_20679_3873 n2_20679_3895 1.396825e-02
R15238 n2_20679_3895 n2_20679_3906 6.984127e-03
R15239 n2_20679_3906 n2_20679_4089 1.161905e-01
R15240 n2_20679_4089 n2_20679_4122 2.095238e-02
R15241 n2_20679_4122 n2_20679_4305 1.161905e-01
R15242 n2_20679_4305 n2_20679_4338 2.095238e-02
R15243 n2_20679_4338 n2_20679_4521 1.161905e-01
R15244 n2_20679_4521 n2_20679_4554 2.095238e-02
R15245 n2_20679_4554 n2_20679_4737 1.161905e-01
R15246 n2_20679_4737 n2_20679_4770 2.095238e-02
R15247 n2_20679_5169 n2_20679_5202 2.095238e-02
R15248 n2_20679_5202 n2_20679_5385 1.161905e-01
R15249 n2_20679_5385 n2_20679_5418 2.095238e-02
R15250 n2_20679_5418 n2_20679_5601 1.161905e-01
R15251 n2_20679_5601 n2_20679_5634 2.095238e-02
R15252 n2_20679_5634 n2_20679_5671 2.349206e-02
R15253 n2_20679_5671 n2_20679_5817 9.269841e-02
R15254 n2_20679_5817 n2_20679_5850 2.095238e-02
R15255 n2_20679_5850 n2_20679_6033 1.161905e-01
R15256 n2_20679_6033 n2_20679_6049 1.015873e-02
R15257 n2_20679_6049 n2_20679_6066 1.079365e-02
R15258 n2_20679_6066 n2_20679_6145 5.015873e-02
R15259 n2_20679_6145 n2_20679_6249 6.603175e-02
R15260 n2_20679_6249 n2_20679_6282 2.095238e-02
R15261 n2_20679_6282 n2_20679_6319 2.349206e-02
R15262 n2_20679_6319 n2_20679_6465 9.269841e-02
R15263 n2_20679_6465 n2_20679_6498 2.095238e-02
R15264 n2_20679_6498 n2_20679_6681 1.161905e-01
R15265 n2_20679_6681 n2_20679_6714 2.095238e-02
R15266 n2_20679_6714 n2_20679_6897 1.161905e-01
R15267 n2_20679_6897 n2_20679_6930 2.095238e-02
R15268 n2_20679_6930 n2_20679_7113 1.161905e-01
R15269 n2_20679_7329 n2_20679_7362 2.095238e-02
R15270 n2_20679_7362 n2_20679_7545 1.161905e-01
R15271 n2_20679_7545 n2_20679_7578 2.095238e-02
R15272 n2_20679_7578 n2_20679_7761 1.161905e-01
R15273 n2_20679_7761 n2_20679_7794 2.095238e-02
R15274 n2_20679_7794 n2_20679_7977 1.161905e-01
R15275 n2_20679_7977 n2_20679_8010 2.095238e-02
R15276 n2_20679_8010 n2_20679_8193 1.161905e-01
R15277 n2_20679_8193 n2_20679_8226 2.095238e-02
R15278 n2_20679_8226 n2_20679_8299 4.634921e-02
R15279 n2_20679_8299 n2_20679_8395 6.095238e-02
R15280 n2_20679_8395 n2_20679_8409 8.888889e-03
R15281 n2_20679_8409 n2_20679_8442 2.095238e-02
R15282 n2_20679_8442 n2_20679_8625 1.161905e-01
R15283 n2_20679_8625 n2_20679_8658 2.095238e-02
R15284 n2_20679_8658 n2_20679_8841 1.161905e-01
R15285 n2_20679_8841 n2_20679_8874 2.095238e-02
R15286 n2_20679_8874 n2_20679_9057 1.161905e-01
R15287 n2_20679_9057 n2_20679_9090 2.095238e-02
R15288 n2_20679_9090 n2_20679_9213 7.809524e-02
R15289 n2_20679_10549 n2_20679_10645 6.095238e-02
R15290 n2_20679_11956 n2_20679_12081 7.936508e-02
R15291 n2_20679_12081 n2_20679_12114 2.095238e-02
R15292 n2_20679_12114 n2_20679_12297 1.161905e-01
R15293 n2_20679_12297 n2_20679_12330 2.095238e-02
R15294 n2_20679_12330 n2_20679_12513 1.161905e-01
R15295 n2_20679_12513 n2_20679_12546 2.095238e-02
R15296 n2_20679_12546 n2_20679_12729 1.161905e-01
R15297 n2_20679_12729 n2_20679_12762 2.095238e-02
R15298 n2_20679_12762 n2_20679_12799 2.349206e-02
R15299 n2_20679_12799 n2_20679_12895 6.095238e-02
R15300 n2_20679_12895 n2_20679_12945 3.174603e-02
R15301 n2_20679_12945 n2_20679_12978 2.095238e-02
R15302 n2_20679_12978 n2_20679_13161 1.161905e-01
R15303 n2_20679_13161 n2_20679_13194 2.095238e-02
R15304 n2_20679_13194 n2_20679_13377 1.161905e-01
R15305 n2_20679_13377 n2_20679_13410 2.095238e-02
R15306 n2_20679_13410 n2_20679_13593 1.161905e-01
R15307 n2_20679_13593 n2_20679_13626 2.095238e-02
R15308 n2_20679_13626 n2_20679_13809 1.161905e-01
R15309 n2_20679_13809 n2_20679_13842 2.095238e-02
R15310 n2_20679_14241 n2_20679_14274 2.095238e-02
R15311 n2_20679_14274 n2_20679_14457 1.161905e-01
R15312 n2_20679_14457 n2_20679_14490 2.095238e-02
R15313 n2_20679_14490 n2_20679_14673 1.161905e-01
R15314 n2_20679_14673 n2_20679_14706 2.095238e-02
R15315 n2_20679_14706 n2_20679_14889 1.161905e-01
R15316 n2_20679_14889 n2_20679_14922 2.095238e-02
R15317 n2_20679_14922 n2_20679_14936 8.888889e-03
R15318 n2_20679_14936 n2_20679_15049 7.174603e-02
R15319 n2_20679_15049 n2_20679_15105 3.555556e-02
R15320 n2_20679_15105 n2_20679_15138 2.095238e-02
R15321 n2_20679_15138 n2_20679_15145 4.444444e-03
R15322 n2_20679_15145 n2_20679_15152 4.444444e-03
R15323 n2_20679_15152 n2_20679_15321 1.073016e-01
R15324 n2_20679_15321 n2_20679_15354 2.095238e-02
R15325 n2_20679_15354 n2_20679_15537 1.161905e-01
R15326 n2_20679_15537 n2_20679_15570 2.095238e-02
R15327 n2_20679_15570 n2_20679_15753 1.161905e-01
R15328 n2_20679_15753 n2_20679_15786 2.095238e-02
R15329 n2_20679_15786 n2_20679_15969 1.161905e-01
R15330 n2_20679_15969 n2_20679_16002 2.095238e-02
R15331 n2_20679_16401 n2_20679_16434 2.095238e-02
R15332 n2_20679_16434 n2_20679_16617 1.161905e-01
R15333 n2_20679_16617 n2_20679_16650 2.095238e-02
R15334 n2_20679_16650 n2_20679_16687 2.349206e-02
R15335 n2_20679_16687 n2_20679_16833 9.269841e-02
R15336 n2_20679_16833 n2_20679_16866 2.095238e-02
R15337 n2_20679_16866 n2_20679_17049 1.161905e-01
R15338 n2_20679_17049 n2_20679_17082 2.095238e-02
R15339 n2_20679_17082 n2_20679_17265 1.161905e-01
R15340 n2_20679_17265 n2_20679_17298 2.095238e-02
R15341 n2_20679_17298 n2_20679_17299 6.349206e-04
R15342 n2_20679_17299 n2_20679_17395 6.095238e-02
R15343 n2_20679_17395 n2_20679_17481 5.460317e-02
R15344 n2_20679_17481 n2_20679_17514 2.095238e-02
R15345 n2_20679_17514 n2_20679_17697 1.161905e-01
R15346 n2_20679_17697 n2_20679_17730 2.095238e-02
R15347 n2_20679_17730 n2_20679_17913 1.161905e-01
R15348 n2_20679_17913 n2_20679_17946 2.095238e-02
R15349 n2_20679_17946 n2_20679_18129 1.161905e-01
R15350 n2_20679_18129 n2_20679_18162 2.095238e-02
R15351 n2_20679_18162 n2_20679_18345 1.161905e-01
R15352 n2_20679_18594 n2_20679_18777 1.161905e-01
R15353 n2_20679_18777 n2_20679_18810 2.095238e-02
R15354 n2_20679_18810 n2_20679_18993 1.161905e-01
R15355 n2_20679_18993 n2_20679_19026 2.095238e-02
R15356 n2_20679_19026 n2_20679_19040 8.888889e-03
R15357 n2_20679_19040 n2_20679_19209 1.073016e-01
R15358 n2_20679_19209 n2_20679_19242 2.095238e-02
R15359 n2_20679_19242 n2_20679_19425 1.161905e-01
R15360 n2_20679_19425 n2_20679_19458 2.095238e-02
R15361 n2_20679_19458 n2_20679_19549 5.777778e-02
R15362 n2_20679_19549 n2_20679_19641 5.841270e-02
R15363 n2_20679_19641 n2_20679_19645 2.539683e-03
R15364 n2_20679_19645 n2_20679_19674 1.841270e-02
R15365 n2_20679_19674 n2_20679_19857 1.161905e-01
R15366 n2_20679_19857 n2_20679_19890 2.095238e-02
R15367 n2_20679_19890 n2_20679_20073 1.161905e-01
R15368 n2_20679_20073 n2_20679_20106 2.095238e-02
R15369 n2_20679_20106 n2_20679_20289 1.161905e-01
R15370 n2_20679_20289 n2_20679_20322 2.095238e-02
R15371 n2_20679_20322 n2_20679_20505 1.161905e-01
R15372 n2_20679_20505 n2_20679_20538 2.095238e-02
R15373 n2_20630_12799 n2_20630_12846 9.400000e-02
R15374 n2_20630_12846 n2_20630_12895 9.800000e-02
R15375 n2_19505_12799 n2_19505_12846 9.400000e-02
R15376 n2_19505_12846 n2_19505_12895 9.800000e-02
R15377 n2_18380_12799 n2_18380_12846 9.400000e-02
R15378 n2_18380_12846 n2_18380_12895 9.800000e-02
R15379 n2_17255_12799 n2_17255_12846 9.400000e-02
R15380 n2_17255_12846 n2_17255_12895 9.800000e-02
R15381 n2_16130_12776 n2_16130_12799 4.600000e-02
R15382 n2_16130_12799 n2_16130_12846 9.400000e-02
R15383 n2_16130_12846 n2_16130_12895 9.800000e-02
R15384 n2_15005_12776 n2_15005_12799 4.600000e-02
R15385 n2_15005_12799 n2_15005_12846 9.400000e-02
R15386 n2_15005_12846 n2_15005_12895 9.800000e-02
R15387 n2_13880_12776 n2_13880_12799 4.600000e-02
R15388 n2_13880_12799 n2_13880_12846 9.400000e-02
R15389 n2_13880_12846 n2_13880_12895 9.800000e-02
R15390 n2_20630_15049 n2_20630_15096 9.400000e-02
R15391 n2_20630_15096 n2_20630_15105 1.800000e-02
R15392 n2_20630_15105 n2_20630_15138 6.600000e-02
R15393 n2_20630_15138 n2_20630_15145 1.400000e-02
R15394 n2_20630_15145 n2_20630_15152 1.400000e-02
R15395 n2_19505_15049 n2_19505_15096 9.400000e-02
R15396 n2_19505_15096 n2_19505_15105 1.800000e-02
R15397 n2_19505_15105 n2_19505_15138 6.600000e-02
R15398 n2_19505_15138 n2_19505_15145 1.400000e-02
R15399 n2_19505_15145 n2_19505_15152 1.400000e-02
R15400 n2_18380_15049 n2_18380_15096 9.400000e-02
R15401 n2_18380_15096 n2_18380_15105 1.800000e-02
R15402 n2_18380_15105 n2_18380_15138 6.600000e-02
R15403 n2_18380_15138 n2_18380_15145 1.400000e-02
R15404 n2_18380_15145 n2_18380_15152 1.400000e-02
R15405 n2_17255_15049 n2_17255_15096 9.400000e-02
R15406 n2_17255_15096 n2_17255_15105 1.800000e-02
R15407 n2_17255_15105 n2_17255_15138 6.600000e-02
R15408 n2_17255_15138 n2_17255_15145 1.400000e-02
R15409 n2_17255_15145 n2_17255_15152 1.400000e-02
R15410 n2_17255_15152 n2_17255_15159 1.400000e-02
R15411 n2_16130_15049 n2_16130_15096 9.400000e-02
R15412 n2_16130_15096 n2_16130_15105 1.800000e-02
R15413 n2_16130_15105 n2_16130_15138 6.600000e-02
R15414 n2_16130_15138 n2_16130_15145 1.400000e-02
R15415 n2_16130_15145 n2_16130_15159 2.800000e-02
R15416 n2_20630_17298 n2_20630_17299 2.000000e-03
R15417 n2_20630_17299 n2_20630_17346 9.400000e-02
R15418 n2_20630_17346 n2_20630_17395 9.800000e-02
R15419 n2_19505_17298 n2_19505_17299 2.000000e-03
R15420 n2_19505_17299 n2_19505_17346 9.400000e-02
R15421 n2_19505_17346 n2_19505_17395 9.800000e-02
R15422 n2_18380_17298 n2_18380_17299 2.000000e-03
R15423 n2_18380_17299 n2_18380_17346 9.400000e-02
R15424 n2_18380_17346 n2_18380_17395 9.800000e-02
R15425 n2_20630_19549 n2_20630_19596 9.400000e-02
R15426 n2_20630_19596 n2_20630_19641 9.000000e-02
R15427 n2_20630_19641 n2_20630_19645 8.000000e-03
R15428 n2_20630_19645 n2_20630_19674 5.800000e-02
R15429 n2_19505_20674 n2_19505_20721 9.400000e-02
R15430 n2_19505_20721 n2_19505_20754 6.600000e-02
R15431 n2_19505_20754 n2_19505_20770 3.200000e-02
R15432 n2_17255_20674 n2_17255_20721 9.400000e-02
R15433 n2_17255_20721 n2_17255_20754 6.600000e-02
R15434 n2_17255_20754 n2_17255_20770 3.200000e-02
R15435 n2_17255_19549 n2_17255_19596 9.400000e-02
R15436 n2_17255_19596 n2_17255_19641 9.000000e-02
R15437 n2_17255_19641 n2_17255_19645 8.000000e-03
R15438 n2_17255_19645 n2_17255_19674 5.800000e-02
R15439 n2_17255_18424 n2_17255_18471 9.400000e-02
R15440 n2_17255_18471 n2_17255_18520 9.800000e-02
R15441 n2_17255_17298 n2_17255_17299 2.000000e-03
R15442 n2_17255_17299 n2_17255_17346 9.400000e-02
R15443 n2_17255_17346 n2_17255_17395 9.800000e-02
R15444 n2_15005_20674 n2_15005_20721 9.400000e-02
R15445 n2_15005_20721 n2_15005_20754 6.600000e-02
R15446 n2_15005_20754 n2_15005_20770 3.200000e-02
R15447 n2_15005_19549 n2_15005_19596 9.400000e-02
R15448 n2_15005_19596 n2_15005_19641 9.000000e-02
R15449 n2_15005_19641 n2_15005_19645 8.000000e-03
R15450 n2_15005_19645 n2_15005_19674 5.800000e-02
R15451 n2_15005_18424 n2_15005_18471 9.400000e-02
R15452 n2_15005_18471 n2_15005_18520 9.800000e-02
R15453 n2_15005_17298 n2_15005_17299 2.000000e-03
R15454 n2_15005_17299 n2_15005_17346 9.400000e-02
R15455 n2_15005_17346 n2_15005_17395 9.800000e-02
R15456 n2_15005_16174 n2_15005_16185 2.200000e-02
R15457 n2_15005_16185 n2_15005_16218 6.600000e-02
R15458 n2_15005_16218 n2_15005_16221 6.000000e-03
R15459 n2_15005_16221 n2_15005_16270 9.800000e-02
R15460 n2_15005_15049 n2_15005_15096 9.400000e-02
R15461 n2_15005_15096 n2_15005_15105 1.800000e-02
R15462 n2_15005_15105 n2_15005_15138 6.600000e-02
R15463 n2_15005_15138 n2_15005_15145 1.400000e-02
R15464 n2_15005_15145 n2_15005_15159 2.800000e-02
R15465 n2_12755_20674 n2_12755_20721 9.400000e-02
R15466 n2_12755_20721 n2_12755_20754 6.600000e-02
R15467 n2_12755_20754 n2_12755_20770 3.200000e-02
R15468 n2_12755_19549 n2_12755_19596 9.400000e-02
R15469 n2_12755_19596 n2_12755_19641 9.000000e-02
R15470 n2_12755_19641 n2_12755_19645 8.000000e-03
R15471 n2_12755_19645 n2_12755_19674 5.800000e-02
R15472 n2_12755_18424 n2_12755_18471 9.400000e-02
R15473 n2_12755_18471 n2_12755_18520 9.800000e-02
R15474 n2_12755_17298 n2_12755_17299 2.000000e-03
R15475 n2_12755_17299 n2_12755_17346 9.400000e-02
R15476 n2_12755_17346 n2_12755_17395 9.800000e-02
R15477 n2_12755_16174 n2_12755_16185 2.200000e-02
R15478 n2_12755_16185 n2_12755_16218 6.600000e-02
R15479 n2_12755_16218 n2_12755_16221 6.000000e-03
R15480 n2_12755_16221 n2_12755_16270 9.800000e-02
R15481 n2_12755_15049 n2_12755_15096 9.400000e-02
R15482 n2_12755_15096 n2_12755_15105 1.800000e-02
R15483 n2_12755_15105 n2_12755_15138 6.600000e-02
R15484 n2_12755_15138 n2_12755_15145 1.400000e-02
R15485 n2_12755_13924 n2_12755_13971 9.400000e-02
R15486 n2_12755_13971 n2_12755_14020 9.800000e-02
R15487 n2_12755_14020 n2_12755_14025 1.000000e-02
R15488 n2_12755_12799 n2_12755_12846 9.400000e-02
R15489 n2_12755_12846 n2_12755_12895 9.800000e-02
R15490 n2_10505_20674 n2_10505_20721 9.400000e-02
R15491 n2_10505_20721 n2_10505_20754 6.600000e-02
R15492 n2_10505_20754 n2_10505_20770 3.200000e-02
R15493 n2_10505_19549 n2_10505_19596 9.400000e-02
R15494 n2_10505_19596 n2_10505_19641 9.000000e-02
R15495 n2_10505_19641 n2_10505_19645 8.000000e-03
R15496 n2_10505_19645 n2_10505_19674 5.800000e-02
R15497 n2_10505_18392 n2_10505_18424 6.400000e-02
R15498 n2_10505_18424 n2_10505_18471 9.400000e-02
R15499 n2_10505_18471 n2_10505_18520 9.800000e-02
R15500 n2_10505_17298 n2_10505_17299 2.000000e-03
R15501 n2_10505_17299 n2_10505_17312 2.600000e-02
R15502 n2_10505_17312 n2_10505_17346 6.800000e-02
R15503 n2_10505_17346 n2_10505_17395 9.800000e-02
R15504 n2_10505_16174 n2_10505_16185 2.200000e-02
R15505 n2_10505_16185 n2_10505_16218 6.600000e-02
R15506 n2_10505_16218 n2_10505_16221 6.000000e-03
R15507 n2_10505_16221 n2_10505_16270 9.800000e-02
R15508 n2_10505_15049 n2_10505_15096 9.400000e-02
R15509 n2_10505_15096 n2_10505_15105 1.800000e-02
R15510 n2_10505_15105 n2_10505_15138 6.600000e-02
R15511 n2_10505_15138 n2_10505_15145 1.400000e-02
R15512 n2_10505_13924 n2_10505_13971 9.400000e-02
R15513 n2_10505_13971 n2_10505_14020 9.800000e-02
R15514 n2_10505_14020 n2_10505_14025 1.000000e-02
R15515 n2_10505_12799 n2_10505_12846 9.400000e-02
R15516 n2_10505_12846 n2_10505_12895 9.800000e-02
R15517 n2_10505_11649 n2_10505_11674 5.000000e-02
R15518 n2_10505_11674 n2_10505_11682 1.600000e-02
R15519 n2_10505_11682 n2_10505_11721 7.800000e-02
R15520 n2_10505_11721 n2_10505_11770 9.800000e-02
R15521 n2_8255_20674 n2_8255_20721 9.400000e-02
R15522 n2_8255_20721 n2_8255_20754 6.600000e-02
R15523 n2_8255_20754 n2_8255_20770 3.200000e-02
R15524 n2_8255_19549 n2_8255_19596 9.400000e-02
R15525 n2_8255_19596 n2_8255_19641 9.000000e-02
R15526 n2_8255_19641 n2_8255_19645 8.000000e-03
R15527 n2_8255_19645 n2_8255_19674 5.800000e-02
R15528 n2_8255_18392 n2_8255_18421 5.800000e-02
R15529 n2_8255_18421 n2_8255_18424 6.000000e-03
R15530 n2_8255_18424 n2_8255_18471 9.400000e-02
R15531 n2_8255_18471 n2_8255_18520 9.800000e-02
R15532 n2_8255_17298 n2_8255_17299 2.000000e-03
R15533 n2_8255_17299 n2_8255_17312 2.600000e-02
R15534 n2_8255_17312 n2_8255_17346 6.800000e-02
R15535 n2_8255_17346 n2_8255_17395 9.800000e-02
R15536 n2_8255_16174 n2_8255_16185 2.200000e-02
R15537 n2_8255_16185 n2_8255_16218 6.600000e-02
R15538 n2_8255_16218 n2_8255_16221 6.000000e-03
R15539 n2_8255_16221 n2_8255_16270 9.800000e-02
R15540 n2_8255_15049 n2_8255_15096 9.400000e-02
R15541 n2_8255_15096 n2_8255_15105 1.800000e-02
R15542 n2_8255_15105 n2_8255_15138 6.600000e-02
R15543 n2_8255_15138 n2_8255_15145 1.400000e-02
R15544 n2_8255_13924 n2_8255_13971 9.400000e-02
R15545 n2_8255_13971 n2_8255_14020 9.800000e-02
R15546 n2_8255_14020 n2_8255_14025 1.000000e-02
R15547 n2_6005_20674 n2_6005_20721 9.400000e-02
R15548 n2_6005_20721 n2_6005_20754 6.600000e-02
R15549 n2_6005_20754 n2_6005_20770 3.200000e-02
R15550 n2_6005_19549 n2_6005_19596 9.400000e-02
R15551 n2_6005_19596 n2_6005_19641 9.000000e-02
R15552 n2_6005_19641 n2_6005_19645 8.000000e-03
R15553 n2_6005_19645 n2_6005_19674 5.800000e-02
R15554 n2_6005_18392 n2_6005_18424 6.400000e-02
R15555 n2_6005_18424 n2_6005_18471 9.400000e-02
R15556 n2_6005_18471 n2_6005_18520 9.800000e-02
R15557 n2_6005_17298 n2_6005_17299 2.000000e-03
R15558 n2_6005_17299 n2_6005_17312 2.600000e-02
R15559 n2_6005_17312 n2_6005_17335 4.600000e-02
R15560 n2_6005_17335 n2_6005_17346 2.200000e-02
R15561 n2_6005_17346 n2_6005_17395 9.800000e-02
R15562 n2_6005_16174 n2_6005_16185 2.200000e-02
R15563 n2_6005_16185 n2_6005_16218 6.600000e-02
R15564 n2_6005_16218 n2_6005_16221 6.000000e-03
R15565 n2_6005_16221 n2_6005_16270 9.800000e-02
R15566 n2_3755_20674 n2_3755_20721 9.400000e-02
R15567 n2_3755_20721 n2_3755_20754 6.600000e-02
R15568 n2_3755_20754 n2_3755_20770 3.200000e-02
R15569 n2_3755_19549 n2_3755_19596 9.400000e-02
R15570 n2_3755_19596 n2_3755_19641 9.000000e-02
R15571 n2_3755_19641 n2_3755_19645 8.000000e-03
R15572 n2_3755_19645 n2_3755_19674 5.800000e-02
R15573 n2_3755_18424 n2_3755_18471 9.400000e-02
R15574 n2_3755_18471 n2_3755_18520 9.800000e-02
R15575 n2_1505_20674 n2_1505_20721 9.400000e-02
R15576 n2_1505_20721 n2_1505_20754 6.600000e-02
R15577 n2_1505_20754 n2_1505_20770 3.200000e-02
R15578 n2_380_19549 n2_380_19596 9.400000e-02
R15579 n2_380_19596 n2_380_19641 9.000000e-02
R15580 n2_380_19641 n2_380_19645 8.000000e-03
R15581 n2_380_19645 n2_380_19674 5.800000e-02
R15582 n2_380_17298 n2_380_17299 2.000000e-03
R15583 n2_380_17299 n2_380_17346 9.400000e-02
R15584 n2_380_17346 n2_380_17395 9.800000e-02
R15585 n2_1505_17298 n2_1505_17299 2.000000e-03
R15586 n2_1505_17299 n2_1505_17346 9.400000e-02
R15587 n2_1505_17346 n2_1505_17395 9.800000e-02
R15588 n2_2630_17298 n2_2630_17299 2.000000e-03
R15589 n2_2630_17299 n2_2630_17346 9.400000e-02
R15590 n2_2630_17346 n2_2630_17395 9.800000e-02
R15591 n2_3755_17298 n2_3755_17299 2.000000e-03
R15592 n2_3755_17299 n2_3755_17335 7.200000e-02
R15593 n2_3755_17335 n2_3755_17346 2.200000e-02
R15594 n2_3755_17346 n2_3755_17395 9.800000e-02
R15595 n2_380_15049 n2_380_15096 9.400000e-02
R15596 n2_380_15096 n2_380_15105 1.800000e-02
R15597 n2_380_15105 n2_380_15138 6.600000e-02
R15598 n2_380_15138 n2_380_15145 1.400000e-02
R15599 n2_1505_15049 n2_1505_15096 9.400000e-02
R15600 n2_1505_15096 n2_1505_15105 1.800000e-02
R15601 n2_1505_15105 n2_1505_15138 6.600000e-02
R15602 n2_1505_15138 n2_1505_15145 1.400000e-02
R15603 n2_2630_15049 n2_2630_15096 9.400000e-02
R15604 n2_2630_15096 n2_2630_15105 1.800000e-02
R15605 n2_2630_15105 n2_2630_15138 6.600000e-02
R15606 n2_2630_15138 n2_2630_15145 1.400000e-02
R15607 n2_3755_15049 n2_3755_15096 9.400000e-02
R15608 n2_3755_15096 n2_3755_15105 1.800000e-02
R15609 n2_3755_15105 n2_3755_15138 6.600000e-02
R15610 n2_3755_15138 n2_3755_15145 1.400000e-02
R15611 n2_4880_15049 n2_4880_15096 9.400000e-02
R15612 n2_4880_15096 n2_4880_15105 1.800000e-02
R15613 n2_4880_15105 n2_4880_15138 6.600000e-02
R15614 n2_4880_15138 n2_4880_15145 1.400000e-02
R15615 n2_6005_15049 n2_6005_15096 9.400000e-02
R15616 n2_6005_15096 n2_6005_15105 1.800000e-02
R15617 n2_6005_15105 n2_6005_15138 6.600000e-02
R15618 n2_6005_15138 n2_6005_15145 1.400000e-02
R15619 n2_380_12799 n2_380_12846 9.400000e-02
R15620 n2_380_12846 n2_380_12895 9.800000e-02
R15621 n2_1505_12799 n2_1505_12846 9.400000e-02
R15622 n2_1505_12846 n2_1505_12895 9.800000e-02
R15623 n2_2630_12799 n2_2630_12846 9.400000e-02
R15624 n2_2630_12846 n2_2630_12895 9.800000e-02
R15625 n2_3755_12799 n2_3755_12846 9.400000e-02
R15626 n2_3755_12846 n2_3755_12895 9.800000e-02
R15627 n2_4880_12799 n2_4880_12846 9.400000e-02
R15628 n2_4880_12846 n2_4880_12895 9.800000e-02
R15629 n2_6005_12799 n2_6005_12846 9.400000e-02
R15630 n2_6005_12846 n2_6005_12895 9.800000e-02
R15631 n2_7130_12799 n2_7130_12846 9.400000e-02
R15632 n2_7130_12846 n2_7130_12895 9.800000e-02
R15633 n2_8255_12799 n2_8255_12846 9.400000e-02
R15634 n2_8255_12846 n2_8255_12895 9.800000e-02
R15635 n2_380_10549 n2_380_10569 4.000000e-02
R15636 n2_380_10569 n2_380_10596 5.400000e-02
R15637 n2_380_10596 n2_380_10602 1.200000e-02
R15638 n2_380_10602 n2_380_10645 8.600000e-02
R15639 n2_1505_10549 n2_1505_10569 4.000000e-02
R15640 n2_1505_10569 n2_1505_10596 5.400000e-02
R15641 n2_1505_10596 n2_1505_10602 1.200000e-02
R15642 n2_1505_10602 n2_1505_10645 8.600000e-02
R15643 n2_2630_10549 n2_2630_10569 4.000000e-02
R15644 n2_2630_10569 n2_2630_10596 5.400000e-02
R15645 n2_2630_10596 n2_2630_10602 1.200000e-02
R15646 n2_2630_10602 n2_2630_10645 8.600000e-02
R15647 n2_3755_10549 n2_3755_10569 4.000000e-02
R15648 n2_3755_10569 n2_3755_10596 5.400000e-02
R15649 n2_3755_10596 n2_3755_10602 1.200000e-02
R15650 n2_3755_10602 n2_3755_10645 8.600000e-02
R15651 n2_4880_10549 n2_4880_10569 4.000000e-02
R15652 n2_4880_10569 n2_4880_10596 5.400000e-02
R15653 n2_4880_10596 n2_4880_10602 1.200000e-02
R15654 n2_4880_10602 n2_4880_10645 8.600000e-02
R15655 n2_6005_10549 n2_6005_10569 4.000000e-02
R15656 n2_6005_10569 n2_6005_10596 5.400000e-02
R15657 n2_6005_10596 n2_6005_10602 1.200000e-02
R15658 n2_6005_10602 n2_6005_10645 8.600000e-02
R15659 n2_7130_10549 n2_7130_10569 4.000000e-02
R15660 n2_7130_10569 n2_7130_10596 5.400000e-02
R15661 n2_7130_10596 n2_7130_10602 1.200000e-02
R15662 n2_7130_10602 n2_7130_10645 8.600000e-02
R15663 n2_8255_10549 n2_8255_10569 4.000000e-02
R15664 n2_8255_10569 n2_8255_10596 5.400000e-02
R15665 n2_8255_10596 n2_8255_10602 1.200000e-02
R15666 n2_8255_10602 n2_8255_10645 8.600000e-02
R15667 n2_9380_10549 n2_9380_10569 4.000000e-02
R15668 n2_9380_10569 n2_9380_10596 5.400000e-02
R15669 n2_9380_10596 n2_9380_10602 1.200000e-02
R15670 n2_9380_10602 n2_9380_10645 8.600000e-02
R15671 n2_12755_417 n2_12755_424 1.400000e-02
R15672 n2_12755_424 n2_12755_450 5.200000e-02
R15673 n2_12755_450 n2_12755_471 4.200000e-02
R15674 n2_12755_471 n2_12755_520 9.800000e-02
R15675 n2_12755_1530 n2_12755_1549 3.800000e-02
R15676 n2_12755_1549 n2_12755_1596 9.400000e-02
R15677 n2_12755_1596 n2_12755_1645 9.800000e-02
R15678 n2_12755_2674 n2_12755_2721 9.400000e-02
R15679 n2_12755_2721 n2_12755_2770 9.800000e-02
R15680 n2_12755_2770 n2_12755_2793 4.600000e-02
R15681 n2_12755_3799 n2_12755_3846 9.400000e-02
R15682 n2_12755_3846 n2_12755_3873 5.400000e-02
R15683 n2_12755_3873 n2_12755_3895 4.400000e-02
R15684 n2_12755_3895 n2_12755_3906 2.200000e-02
R15685 n2_12755_4924 n2_12755_4953 5.800000e-02
R15686 n2_12755_4953 n2_12755_4971 3.600000e-02
R15687 n2_12755_4971 n2_12755_4986 3.000000e-02
R15688 n2_12755_4986 n2_12755_5020 6.800000e-02
R15689 n2_12755_5020 n2_12755_5023 6.000000e-03
R15690 n2_12755_6033 n2_12755_6049 3.200000e-02
R15691 n2_12755_6049 n2_12755_6066 3.400000e-02
R15692 n2_12755_6066 n2_12755_6096 6.000000e-02
R15693 n2_12755_6096 n2_12755_6145 9.800000e-02
R15694 n2_12755_7146 n2_12755_7174 5.600000e-02
R15695 n2_12755_7174 n2_12755_7178 8.000000e-03
R15696 n2_12755_7178 n2_12755_7221 8.600000e-02
R15697 n2_12755_7221 n2_12755_7270 9.800000e-02
R15698 n2_15005_417 n2_15005_424 1.400000e-02
R15699 n2_15005_424 n2_15005_450 5.200000e-02
R15700 n2_15005_450 n2_15005_471 4.200000e-02
R15701 n2_15005_471 n2_15005_520 9.800000e-02
R15702 n2_15005_1530 n2_15005_1549 3.800000e-02
R15703 n2_15005_1549 n2_15005_1596 9.400000e-02
R15704 n2_15005_1596 n2_15005_1645 9.800000e-02
R15705 n2_15005_2674 n2_15005_2721 9.400000e-02
R15706 n2_15005_2721 n2_15005_2770 9.800000e-02
R15707 n2_15005_2770 n2_15005_2793 4.600000e-02
R15708 n2_15005_3799 n2_15005_3846 9.400000e-02
R15709 n2_15005_3846 n2_15005_3873 5.400000e-02
R15710 n2_15005_3873 n2_15005_3895 4.400000e-02
R15711 n2_15005_3895 n2_15005_3906 2.200000e-02
R15712 n2_15005_4924 n2_15005_4953 5.800000e-02
R15713 n2_15005_4953 n2_15005_4971 3.600000e-02
R15714 n2_15005_4971 n2_15005_4986 3.000000e-02
R15715 n2_15005_4986 n2_15005_5020 6.800000e-02
R15716 n2_17255_417 n2_17255_424 1.400000e-02
R15717 n2_17255_424 n2_17255_450 5.200000e-02
R15718 n2_17255_450 n2_17255_471 4.200000e-02
R15719 n2_17255_471 n2_17255_520 9.800000e-02
R15720 n2_17255_1530 n2_17255_1549 3.800000e-02
R15721 n2_17255_1549 n2_17255_1596 9.400000e-02
R15722 n2_17255_1596 n2_17255_1645 9.800000e-02
R15723 n2_17255_2674 n2_17255_2721 9.400000e-02
R15724 n2_17255_2721 n2_17255_2770 9.800000e-02
R15725 n2_17255_2770 n2_17255_2793 4.600000e-02
R15726 n2_19505_417 n2_19505_424 1.400000e-02
R15727 n2_19505_424 n2_19505_450 5.200000e-02
R15728 n2_19505_450 n2_19505_471 4.200000e-02
R15729 n2_19505_471 n2_19505_520 9.800000e-02
R15730 n2_20630_1530 n2_20630_1549 3.800000e-02
R15731 n2_20630_1549 n2_20630_1596 9.400000e-02
R15732 n2_20630_1596 n2_20630_1645 9.800000e-02
R15733 n2_20630_3799 n2_20630_3846 9.400000e-02
R15734 n2_20630_3846 n2_20630_3873 5.400000e-02
R15735 n2_20630_3873 n2_20630_3895 4.400000e-02
R15736 n2_20630_3895 n2_20630_3906 2.200000e-02
R15737 n2_19505_3799 n2_19505_3846 9.400000e-02
R15738 n2_19505_3846 n2_19505_3873 5.400000e-02
R15739 n2_19505_3873 n2_19505_3895 4.400000e-02
R15740 n2_19505_3895 n2_19505_3906 2.200000e-02
R15741 n2_18380_3799 n2_18380_3846 9.400000e-02
R15742 n2_18380_3846 n2_18380_3873 5.400000e-02
R15743 n2_18380_3873 n2_18380_3895 4.400000e-02
R15744 n2_18380_3895 n2_18380_3906 2.200000e-02
R15745 n2_17255_3799 n2_17255_3846 9.400000e-02
R15746 n2_17255_3846 n2_17255_3873 5.400000e-02
R15747 n2_17255_3873 n2_17255_3895 4.400000e-02
R15748 n2_17255_3895 n2_17255_3906 2.200000e-02
R15749 n2_20630_6033 n2_20630_6049 3.200000e-02
R15750 n2_20630_6049 n2_20630_6066 3.400000e-02
R15751 n2_20630_6066 n2_20630_6096 6.000000e-02
R15752 n2_20630_6096 n2_20630_6145 9.800000e-02
R15753 n2_19505_6033 n2_19505_6049 3.200000e-02
R15754 n2_19505_6049 n2_19505_6066 3.400000e-02
R15755 n2_19505_6066 n2_19505_6096 6.000000e-02
R15756 n2_19505_6096 n2_19505_6145 9.800000e-02
R15757 n2_18380_6033 n2_18380_6049 3.200000e-02
R15758 n2_18380_6049 n2_18380_6066 3.400000e-02
R15759 n2_18380_6066 n2_18380_6096 6.000000e-02
R15760 n2_18380_6096 n2_18380_6145 9.800000e-02
R15761 n2_17255_6033 n2_17255_6049 3.200000e-02
R15762 n2_17255_6049 n2_17255_6066 3.400000e-02
R15763 n2_17255_6066 n2_17255_6096 6.000000e-02
R15764 n2_17255_6096 n2_17255_6145 9.800000e-02
R15765 n2_16130_6033 n2_16130_6049 3.200000e-02
R15766 n2_16130_6049 n2_16130_6066 3.400000e-02
R15767 n2_16130_6066 n2_16130_6096 6.000000e-02
R15768 n2_16130_6096 n2_16130_6145 9.800000e-02
R15769 n2_15005_6033 n2_15005_6049 3.200000e-02
R15770 n2_15005_6049 n2_15005_6066 3.400000e-02
R15771 n2_15005_6066 n2_15005_6096 6.000000e-02
R15772 n2_15005_6096 n2_15005_6145 9.800000e-02
R15773 n2_20630_8299 n2_20630_8346 9.400000e-02
R15774 n2_20630_8346 n2_20630_8395 9.800000e-02
R15775 n2_20630_8395 n2_20630_8409 2.800000e-02
R15776 n2_19505_8299 n2_19505_8346 9.400000e-02
R15777 n2_19505_8346 n2_19505_8395 9.800000e-02
R15778 n2_19505_8395 n2_19505_8409 2.800000e-02
R15779 n2_18380_8299 n2_18380_8346 9.400000e-02
R15780 n2_18380_8346 n2_18380_8395 9.800000e-02
R15781 n2_18380_8395 n2_18380_8409 2.800000e-02
R15782 n2_17255_8299 n2_17255_8346 9.400000e-02
R15783 n2_17255_8346 n2_17255_8395 9.800000e-02
R15784 n2_17255_8395 n2_17255_8409 2.800000e-02
R15785 n2_16130_8299 n2_16130_8346 9.400000e-02
R15786 n2_16130_8346 n2_16130_8395 9.800000e-02
R15787 n2_16130_8395 n2_16130_8409 2.800000e-02
R15788 n2_15005_8299 n2_15005_8346 9.400000e-02
R15789 n2_15005_8346 n2_15005_8395 9.800000e-02
R15790 n2_15005_8395 n2_15005_8409 2.800000e-02
R15791 n2_13880_8299 n2_13880_8346 9.400000e-02
R15792 n2_13880_8346 n2_13880_8395 9.800000e-02
R15793 n2_13880_8395 n2_13880_8409 2.800000e-02
R15794 n2_12755_8299 n2_12755_8346 9.400000e-02
R15795 n2_12755_8346 n2_12755_8395 9.800000e-02
R15796 n2_12755_8395 n2_12755_8409 2.800000e-02
R15797 n2_20630_10549 n2_20630_10596 9.400000e-02
R15798 n2_20630_10596 n2_20630_10645 9.800000e-02
R15799 n2_19505_10549 n2_19505_10569 4.000000e-02
R15800 n2_19505_10569 n2_19505_10596 5.400000e-02
R15801 n2_19505_10596 n2_19505_10602 1.200000e-02
R15802 n2_19505_10602 n2_19505_10645 8.600000e-02
R15803 n2_18380_10549 n2_18380_10569 4.000000e-02
R15804 n2_18380_10569 n2_18380_10596 5.400000e-02
R15805 n2_18380_10596 n2_18380_10602 1.200000e-02
R15806 n2_18380_10602 n2_18380_10645 8.600000e-02
R15807 n2_17255_10549 n2_17255_10569 4.000000e-02
R15808 n2_17255_10569 n2_17255_10596 5.400000e-02
R15809 n2_17255_10596 n2_17255_10602 1.200000e-02
R15810 n2_17255_10602 n2_17255_10645 8.600000e-02
R15811 n2_16130_10549 n2_16130_10569 4.000000e-02
R15812 n2_16130_10569 n2_16130_10596 5.400000e-02
R15813 n2_16130_10596 n2_16130_10602 1.200000e-02
R15814 n2_16130_10602 n2_16130_10645 8.600000e-02
R15815 n2_15005_10549 n2_15005_10569 4.000000e-02
R15816 n2_15005_10569 n2_15005_10596 5.400000e-02
R15817 n2_15005_10596 n2_15005_10602 1.200000e-02
R15818 n2_15005_10602 n2_15005_10645 8.600000e-02
R15819 n2_13880_10549 n2_13880_10569 4.000000e-02
R15820 n2_13880_10569 n2_13880_10596 5.400000e-02
R15821 n2_13880_10596 n2_13880_10602 1.200000e-02
R15822 n2_13880_10602 n2_13880_10645 8.600000e-02
R15823 n2_12755_10549 n2_12755_10569 4.000000e-02
R15824 n2_12755_10569 n2_12755_10596 5.400000e-02
R15825 n2_12755_10596 n2_12755_10602 1.200000e-02
R15826 n2_12755_10602 n2_12755_10645 8.600000e-02
R15827 n2_11630_10549 n2_11630_10569 4.000000e-02
R15828 n2_11630_10569 n2_11630_10596 5.400000e-02
R15829 n2_11630_10596 n2_11630_10602 1.200000e-02
R15830 n2_11630_10602 n2_11630_10645 8.600000e-02
R15831 n2_1505_417 n2_1505_424 1.400000e-02
R15832 n2_1505_424 n2_1505_450 5.200000e-02
R15833 n2_1505_450 n2_1505_471 4.200000e-02
R15834 n2_1505_471 n2_1505_520 9.800000e-02
R15835 n2_3755_417 n2_3755_424 1.400000e-02
R15836 n2_3755_424 n2_3755_450 5.200000e-02
R15837 n2_3755_450 n2_3755_471 4.200000e-02
R15838 n2_3755_471 n2_3755_520 9.800000e-02
R15839 n2_3755_1530 n2_3755_1549 3.800000e-02
R15840 n2_3755_1549 n2_3755_1596 9.400000e-02
R15841 n2_3755_1596 n2_3755_1645 9.800000e-02
R15842 n2_3755_1645 n2_3755_1652 1.400000e-02
R15843 n2_3755_2674 n2_3755_2721 9.400000e-02
R15844 n2_3755_2721 n2_3755_2770 9.800000e-02
R15845 n2_3755_2770 n2_3755_2793 4.600000e-02
R15846 n2_3755_3799 n2_3755_3846 9.400000e-02
R15847 n2_3755_3846 n2_3755_3873 5.400000e-02
R15848 n2_3755_3873 n2_3755_3895 4.400000e-02
R15849 n2_3755_3895 n2_3755_3906 2.200000e-02
R15850 n2_3755_3906 n2_3755_3920 2.800000e-02
R15851 n2_6005_417 n2_6005_424 1.400000e-02
R15852 n2_6005_424 n2_6005_450 5.200000e-02
R15853 n2_6005_450 n2_6005_471 4.200000e-02
R15854 n2_6005_471 n2_6005_520 9.800000e-02
R15855 n2_6005_1530 n2_6005_1549 3.800000e-02
R15856 n2_6005_1549 n2_6005_1596 9.400000e-02
R15857 n2_6005_1596 n2_6005_1645 9.800000e-02
R15858 n2_6005_2674 n2_6005_2721 9.400000e-02
R15859 n2_6005_2721 n2_6005_2770 9.800000e-02
R15860 n2_6005_2770 n2_6005_2793 4.600000e-02
R15861 n2_6005_3799 n2_6005_3846 9.400000e-02
R15862 n2_6005_3846 n2_6005_3873 5.400000e-02
R15863 n2_6005_3873 n2_6005_3895 4.400000e-02
R15864 n2_6005_3895 n2_6005_3906 2.200000e-02
R15865 n2_6005_4924 n2_6005_4953 5.800000e-02
R15866 n2_6005_4953 n2_6005_4971 3.600000e-02
R15867 n2_6005_4971 n2_6005_4986 3.000000e-02
R15868 n2_6005_4986 n2_6005_5020 6.800000e-02
R15869 n2_6005_6033 n2_6005_6049 3.200000e-02
R15870 n2_6005_6049 n2_6005_6066 3.400000e-02
R15871 n2_6005_6066 n2_6005_6096 6.000000e-02
R15872 n2_6005_6096 n2_6005_6145 9.800000e-02
R15873 n2_8255_417 n2_8255_424 1.400000e-02
R15874 n2_8255_424 n2_8255_450 5.200000e-02
R15875 n2_8255_450 n2_8255_471 4.200000e-02
R15876 n2_8255_471 n2_8255_520 9.800000e-02
R15877 n2_8255_1530 n2_8255_1549 3.800000e-02
R15878 n2_8255_1549 n2_8255_1596 9.400000e-02
R15879 n2_8255_1596 n2_8255_1645 9.800000e-02
R15880 n2_8255_2674 n2_8255_2721 9.400000e-02
R15881 n2_8255_2721 n2_8255_2770 9.800000e-02
R15882 n2_8255_2770 n2_8255_2793 4.600000e-02
R15883 n2_8255_3799 n2_8255_3846 9.400000e-02
R15884 n2_8255_3846 n2_8255_3873 5.400000e-02
R15885 n2_8255_3873 n2_8255_3895 4.400000e-02
R15886 n2_8255_3895 n2_8255_3906 2.200000e-02
R15887 n2_8255_4924 n2_8255_4953 5.800000e-02
R15888 n2_8255_4953 n2_8255_4971 3.600000e-02
R15889 n2_8255_4971 n2_8255_4986 3.000000e-02
R15890 n2_8255_4986 n2_8255_5020 6.800000e-02
R15891 n2_8255_6033 n2_8255_6049 3.200000e-02
R15892 n2_8255_6049 n2_8255_6066 3.400000e-02
R15893 n2_8255_6066 n2_8255_6096 6.000000e-02
R15894 n2_8255_6096 n2_8255_6145 9.800000e-02
R15895 n2_8255_7146 n2_8255_7160 2.800000e-02
R15896 n2_8255_7160 n2_8255_7174 2.800000e-02
R15897 n2_8255_7174 n2_8255_7221 9.400000e-02
R15898 n2_8255_7221 n2_8255_7270 9.800000e-02
R15899 n2_8255_8299 n2_8255_8346 9.400000e-02
R15900 n2_8255_8346 n2_8255_8395 9.800000e-02
R15901 n2_8255_8395 n2_8255_8409 2.800000e-02
R15902 n2_10505_417 n2_10505_424 1.400000e-02
R15903 n2_10505_424 n2_10505_450 5.200000e-02
R15904 n2_10505_450 n2_10505_471 4.200000e-02
R15905 n2_10505_471 n2_10505_520 9.800000e-02
R15906 n2_10505_1530 n2_10505_1549 3.800000e-02
R15907 n2_10505_1549 n2_10505_1596 9.400000e-02
R15908 n2_10505_1596 n2_10505_1645 9.800000e-02
R15909 n2_10505_2647 n2_10505_2674 5.400000e-02
R15910 n2_10505_2674 n2_10505_2721 9.400000e-02
R15911 n2_10505_2721 n2_10505_2770 9.800000e-02
R15912 n2_10505_2770 n2_10505_2793 4.600000e-02
R15913 n2_10505_3799 n2_10505_3846 9.400000e-02
R15914 n2_10505_3846 n2_10505_3873 5.400000e-02
R15915 n2_10505_3873 n2_10505_3895 4.400000e-02
R15916 n2_10505_3895 n2_10505_3906 2.200000e-02
R15917 n2_10505_4924 n2_10505_4953 5.800000e-02
R15918 n2_10505_4953 n2_10505_4971 3.600000e-02
R15919 n2_10505_4971 n2_10505_4986 3.000000e-02
R15920 n2_10505_4986 n2_10505_5020 6.800000e-02
R15921 n2_10505_6033 n2_10505_6049 3.200000e-02
R15922 n2_10505_6049 n2_10505_6066 3.400000e-02
R15923 n2_10505_6066 n2_10505_6096 6.000000e-02
R15924 n2_10505_6096 n2_10505_6145 9.800000e-02
R15925 n2_10505_7146 n2_10505_7160 2.800000e-02
R15926 n2_10505_7160 n2_10505_7174 2.800000e-02
R15927 n2_10505_7174 n2_10505_7178 8.000000e-03
R15928 n2_10505_7178 n2_10505_7221 8.600000e-02
R15929 n2_10505_7221 n2_10505_7270 9.800000e-02
R15930 n2_10505_8299 n2_10505_8346 9.400000e-02
R15931 n2_10505_8346 n2_10505_8395 9.800000e-02
R15932 n2_10505_8395 n2_10505_8409 2.800000e-02
R15933 n2_10505_9424 n2_10505_9471 9.400000e-02
R15934 n2_10505_9471 n2_10505_9489 3.600000e-02
R15935 n2_10505_9489 n2_10505_9520 6.200000e-02
R15936 n2_10505_9520 n2_10505_9522 4.000000e-03
R15937 n2_10505_10549 n2_10505_10569 4.000000e-02
R15938 n2_10505_10569 n2_10505_10596 5.400000e-02
R15939 n2_10505_10596 n2_10505_10602 1.200000e-02
R15940 n2_10505_10602 n2_10505_10645 8.600000e-02
R15941 n2_380_8299 n2_380_8346 9.400000e-02
R15942 n2_380_8346 n2_380_8395 9.800000e-02
R15943 n2_380_8395 n2_380_8409 2.800000e-02
R15944 n2_1505_8299 n2_1505_8346 9.400000e-02
R15945 n2_1505_8346 n2_1505_8395 9.800000e-02
R15946 n2_1505_8395 n2_1505_8409 2.800000e-02
R15947 n2_2630_8299 n2_2630_8346 9.400000e-02
R15948 n2_2630_8346 n2_2630_8395 9.800000e-02
R15949 n2_2630_8395 n2_2630_8409 2.800000e-02
R15950 n2_3755_8299 n2_3755_8346 9.400000e-02
R15951 n2_3755_8346 n2_3755_8395 9.800000e-02
R15952 n2_3755_8395 n2_3755_8409 2.800000e-02
R15953 n2_4880_8299 n2_4880_8346 9.400000e-02
R15954 n2_4880_8346 n2_4880_8395 9.800000e-02
R15955 n2_4880_8395 n2_4880_8409 2.800000e-02
R15956 n2_6005_8299 n2_6005_8346 9.400000e-02
R15957 n2_6005_8346 n2_6005_8395 9.800000e-02
R15958 n2_6005_8395 n2_6005_8409 2.800000e-02
R15959 n2_7130_8299 n2_7130_8346 9.400000e-02
R15960 n2_7130_8346 n2_7130_8395 9.800000e-02
R15961 n2_7130_8395 n2_7130_8409 2.800000e-02
R15962 n2_380_6033 n2_380_6049 3.200000e-02
R15963 n2_380_6049 n2_380_6066 3.400000e-02
R15964 n2_380_6066 n2_380_6096 6.000000e-02
R15965 n2_380_6096 n2_380_6145 9.800000e-02
R15966 n2_1505_6033 n2_1505_6049 3.200000e-02
R15967 n2_1505_6049 n2_1505_6066 3.400000e-02
R15968 n2_1505_6066 n2_1505_6096 6.000000e-02
R15969 n2_1505_6096 n2_1505_6145 9.800000e-02
R15970 n2_2630_6033 n2_2630_6049 3.200000e-02
R15971 n2_2630_6049 n2_2630_6066 3.400000e-02
R15972 n2_2630_6066 n2_2630_6096 6.000000e-02
R15973 n2_2630_6096 n2_2630_6145 9.800000e-02
R15974 n2_3755_6033 n2_3755_6049 3.200000e-02
R15975 n2_3755_6049 n2_3755_6066 3.400000e-02
R15976 n2_3755_6066 n2_3755_6096 6.000000e-02
R15977 n2_3755_6096 n2_3755_6145 9.800000e-02
R15978 n2_4880_6033 n2_4880_6049 3.200000e-02
R15979 n2_4880_6049 n2_4880_6066 3.400000e-02
R15980 n2_4880_6066 n2_4880_6096 6.000000e-02
R15981 n2_4880_6096 n2_4880_6145 9.800000e-02
R15982 n2_380_3799 n2_380_3846 9.400000e-02
R15983 n2_380_3846 n2_380_3873 5.400000e-02
R15984 n2_380_3873 n2_380_3895 4.400000e-02
R15985 n2_380_3895 n2_380_3906 2.200000e-02
R15986 n2_1505_3799 n2_1505_3846 9.400000e-02
R15987 n2_1505_3846 n2_1505_3873 5.400000e-02
R15988 n2_1505_3873 n2_1505_3895 4.400000e-02
R15989 n2_1505_3895 n2_1505_3906 2.200000e-02
R15990 n2_1505_3906 n2_1505_3920 2.800000e-02
R15991 n2_2630_3799 n2_2630_3846 9.400000e-02
R15992 n2_2630_3846 n2_2630_3873 5.400000e-02
R15993 n2_2630_3873 n2_2630_3895 4.400000e-02
R15994 n2_2630_3895 n2_2630_3906 2.200000e-02
R15995 n2_2630_3906 n2_2630_3920 2.800000e-02
R15996 n2_380_1530 n2_380_1549 3.800000e-02
R15997 n2_380_1549 n2_380_1596 9.400000e-02
R15998 n2_380_1596 n2_380_1645 9.800000e-02
v4f _X_n2_10505_16221 0 0
v99 _X_n2_6005_12846 0 0
rr21e n3_13880_13971 _X_n3_13880_13971 2.500000e-01
v147 _X_n2_2630_8346 0 0
v149 _X_n2_3755_8346 0 0
v151 _X_n2_380_6096 0 0
v5b _X_n2_8255_19596 0 0
* vias from: 0 to 2
V15999 n0_241_633 n2_241_633 0.0
V16000 n0_241_666 n2_241_666 0.0
V16001 n0_241_849 n2_241_849 0.0
V16002 n0_241_882 n2_241_882 0.0
V16003 n0_241_1065 n2_241_1065 0.0
V16004 n0_241_1098 n2_241_1098 0.0
V16005 n0_241_1281 n2_241_1281 0.0
V16006 n0_241_1314 n2_241_1314 0.0
V16007 n0_241_1497 n2_241_1497 0.0
V16008 n0_241_1530 n2_241_1530 0.0
V16009 n0_241_1713 n2_241_1713 0.0
V16010 n0_241_1746 n2_241_1746 0.0
V16011 n0_241_1929 n2_241_1929 0.0
V16012 n0_241_1962 n2_241_1962 0.0
V16013 n0_241_2145 n2_241_2145 0.0
V16014 n0_241_2178 n2_241_2178 0.0
V16015 n0_241_2361 n2_241_2361 0.0
V16016 n0_241_2394 n2_241_2394 0.0
V16017 n0_241_2577 n2_241_2577 0.0
V16018 n0_241_2610 n2_241_2610 0.0
V16019 n0_241_2793 n2_241_2793 0.0
V16020 n0_241_2826 n2_241_2826 0.0
V16021 n0_241_3009 n2_241_3009 0.0
V16022 n0_241_3042 n2_241_3042 0.0
V16023 n0_241_3225 n2_241_3225 0.0
V16024 n0_241_3258 n2_241_3258 0.0
V16025 n0_241_3441 n2_241_3441 0.0
V16026 n0_241_3474 n2_241_3474 0.0
V16027 n0_241_3657 n2_241_3657 0.0
V16028 n0_241_3690 n2_241_3690 0.0
V16029 n0_241_3873 n2_241_3873 0.0
V16030 n0_241_3906 n2_241_3906 0.0
V16031 n0_241_4089 n2_241_4089 0.0
V16032 n0_241_4122 n2_241_4122 0.0
V16033 n0_241_4305 n2_241_4305 0.0
V16034 n0_241_4338 n2_241_4338 0.0
V16035 n0_241_4375 n2_241_4375 0.0
V16036 n0_241_4521 n2_241_4521 0.0
V16037 n0_241_4554 n2_241_4554 0.0
V16038 n0_241_4737 n2_241_4737 0.0
V16039 n0_241_4770 n2_241_4770 0.0
V16040 n0_241_4953 n2_241_4953 0.0
V16041 n0_241_4986 n2_241_4986 0.0
V16042 n0_241_5169 n2_241_5169 0.0
V16043 n0_241_5202 n2_241_5202 0.0
V16044 n0_241_5385 n2_241_5385 0.0
V16045 n0_241_5418 n2_241_5418 0.0
V16046 n0_241_5601 n2_241_5601 0.0
V16047 n0_241_5634 n2_241_5634 0.0
V16048 n0_241_5817 n2_241_5817 0.0
V16049 n0_241_5850 n2_241_5850 0.0
V16050 n0_241_6033 n2_241_6033 0.0
V16051 n0_241_6066 n2_241_6066 0.0
V16052 n0_241_6249 n2_241_6249 0.0
V16053 n0_241_6282 n2_241_6282 0.0
V16054 n0_241_6465 n2_241_6465 0.0
V16055 n0_241_6498 n2_241_6498 0.0
V16056 n0_241_6681 n2_241_6681 0.0
V16057 n0_241_6714 n2_241_6714 0.0
V16058 n0_241_6897 n2_241_6897 0.0
V16059 n0_241_6930 n2_241_6930 0.0
V16060 n0_241_7113 n2_241_7113 0.0
V16061 n0_241_7146 n2_241_7146 0.0
V16062 n0_241_7329 n2_241_7329 0.0
V16063 n0_241_7362 n2_241_7362 0.0
V16064 n0_241_7545 n2_241_7545 0.0
V16065 n0_241_7578 n2_241_7578 0.0
V16066 n0_241_7761 n2_241_7761 0.0
V16067 n0_241_7794 n2_241_7794 0.0
V16068 n0_241_7977 n2_241_7977 0.0
V16069 n0_241_8010 n2_241_8010 0.0
V16070 n0_241_8193 n2_241_8193 0.0
V16071 n0_241_8226 n2_241_8226 0.0
V16072 n0_241_8409 n2_241_8409 0.0
V16073 n0_241_8442 n2_241_8442 0.0
V16074 n0_241_8625 n2_241_8625 0.0
V16075 n0_241_8658 n2_241_8658 0.0
V16076 n0_241_8841 n2_241_8841 0.0
V16077 n0_241_8874 n2_241_8874 0.0
V16078 n0_241_9057 n2_241_9057 0.0
V16079 n0_241_9090 n2_241_9090 0.0
V16080 n0_241_9273 n2_241_9273 0.0
V16081 n0_241_9306 n2_241_9306 0.0
V16082 n0_241_9489 n2_241_9489 0.0
V16083 n0_241_9522 n2_241_9522 0.0
V16084 n0_241_9705 n2_241_9705 0.0
V16085 n0_241_9738 n2_241_9738 0.0
V16086 n0_241_9921 n2_241_9921 0.0
V16087 n0_241_9954 n2_241_9954 0.0
V16088 n0_241_10137 n2_241_10137 0.0
V16089 n0_241_10170 n2_241_10170 0.0
V16090 n0_241_10353 n2_241_10353 0.0
V16091 n0_241_10386 n2_241_10386 0.0
V16092 n0_241_10569 n2_241_10569 0.0
V16093 n0_241_10785 n2_241_10785 0.0
V16094 n0_241_10818 n2_241_10818 0.0
V16095 n0_241_11001 n2_241_11001 0.0
V16096 n0_241_11034 n2_241_11034 0.0
V16097 n0_241_11217 n2_241_11217 0.0
V16098 n0_241_11250 n2_241_11250 0.0
V16099 n0_241_11433 n2_241_11433 0.0
V16100 n0_241_11466 n2_241_11466 0.0
V16101 n0_241_11649 n2_241_11649 0.0
V16102 n0_241_11682 n2_241_11682 0.0
V16103 n0_241_11865 n2_241_11865 0.0
V16104 n0_241_11898 n2_241_11898 0.0
V16105 n0_241_12081 n2_241_12081 0.0
V16106 n0_241_12114 n2_241_12114 0.0
V16107 n0_241_12297 n2_241_12297 0.0
V16108 n0_241_12330 n2_241_12330 0.0
V16109 n0_241_12513 n2_241_12513 0.0
V16110 n0_241_12546 n2_241_12546 0.0
V16111 n0_241_12729 n2_241_12729 0.0
V16112 n0_241_12762 n2_241_12762 0.0
V16113 n0_241_12945 n2_241_12945 0.0
V16114 n0_241_12978 n2_241_12978 0.0
V16115 n0_241_13161 n2_241_13161 0.0
V16116 n0_241_13194 n2_241_13194 0.0
V16117 n0_241_13377 n2_241_13377 0.0
V16118 n0_241_13410 n2_241_13410 0.0
V16119 n0_241_13593 n2_241_13593 0.0
V16120 n0_241_13626 n2_241_13626 0.0
V16121 n0_241_13663 n2_241_13663 0.0
V16122 n0_241_13809 n2_241_13809 0.0
V16123 n0_241_13842 n2_241_13842 0.0
V16124 n0_241_14025 n2_241_14025 0.0
V16125 n0_241_14058 n2_241_14058 0.0
V16126 n0_241_14241 n2_241_14241 0.0
V16127 n0_241_14274 n2_241_14274 0.0
V16128 n0_241_14457 n2_241_14457 0.0
V16129 n0_241_14490 n2_241_14490 0.0
V16130 n0_241_14673 n2_241_14673 0.0
V16131 n0_241_14706 n2_241_14706 0.0
V16132 n0_241_14889 n2_241_14889 0.0
V16133 n0_241_14922 n2_241_14922 0.0
V16134 n0_241_15138 n2_241_15138 0.0
V16135 n0_241_15321 n2_241_15321 0.0
V16136 n0_241_15354 n2_241_15354 0.0
V16137 n0_241_15537 n2_241_15537 0.0
V16138 n0_241_15570 n2_241_15570 0.0
V16139 n0_241_15753 n2_241_15753 0.0
V16140 n0_241_15786 n2_241_15786 0.0
V16141 n0_241_15969 n2_241_15969 0.0
V16142 n0_241_16002 n2_241_16002 0.0
V16143 n0_241_16185 n2_241_16185 0.0
V16144 n0_241_16218 n2_241_16218 0.0
V16145 n0_241_16401 n2_241_16401 0.0
V16146 n0_241_16434 n2_241_16434 0.0
V16147 n0_241_16617 n2_241_16617 0.0
V16148 n0_241_16650 n2_241_16650 0.0
V16149 n0_241_16833 n2_241_16833 0.0
V16150 n0_241_16866 n2_241_16866 0.0
V16151 n0_241_17049 n2_241_17049 0.0
V16152 n0_241_17082 n2_241_17082 0.0
V16153 n0_241_17265 n2_241_17265 0.0
V16154 n0_241_17298 n2_241_17298 0.0
V16155 n0_241_17481 n2_241_17481 0.0
V16156 n0_241_17514 n2_241_17514 0.0
V16157 n0_241_17697 n2_241_17697 0.0
V16158 n0_241_17730 n2_241_17730 0.0
V16159 n0_241_17913 n2_241_17913 0.0
V16160 n0_241_17946 n2_241_17946 0.0
V16161 n0_241_17960 n2_241_17960 0.0
V16162 n0_241_18129 n2_241_18129 0.0
V16163 n0_241_18162 n2_241_18162 0.0
V16164 n0_241_18345 n2_241_18345 0.0
V16165 n0_241_18378 n2_241_18378 0.0
V16166 n0_241_18561 n2_241_18561 0.0
V16167 n0_241_18594 n2_241_18594 0.0
V16168 n0_241_18777 n2_241_18777 0.0
V16169 n0_241_18810 n2_241_18810 0.0
V16170 n0_241_18993 n2_241_18993 0.0
V16171 n0_241_19026 n2_241_19026 0.0
V16172 n0_241_19040 n2_241_19040 0.0
V16173 n0_241_19209 n2_241_19209 0.0
V16174 n0_241_19242 n2_241_19242 0.0
V16175 n0_241_19256 n2_241_19256 0.0
V16176 n0_241_19425 n2_241_19425 0.0
V16177 n0_241_19458 n2_241_19458 0.0
V16178 n0_241_19472 n2_241_19472 0.0
V16179 n0_241_19641 n2_241_19641 0.0
V16180 n0_241_19674 n2_241_19674 0.0
V16181 n0_241_19857 n2_241_19857 0.0
V16182 n0_241_19890 n2_241_19890 0.0
V16183 n0_241_20073 n2_241_20073 0.0
V16184 n0_241_20106 n2_241_20106 0.0
V16185 n0_241_20289 n2_241_20289 0.0
V16186 n0_241_20322 n2_241_20322 0.0
V16187 n0_241_20505 n2_241_20505 0.0
V16188 n0_241_20538 n2_241_20538 0.0
V16189 n0_380_1530 n2_380_1530 0.0
V16190 n0_380_3873 n2_380_3873 0.0
V16191 n0_380_3906 n2_380_3906 0.0
V16192 n0_380_6033 n2_380_6033 0.0
V16193 n0_380_6066 n2_380_6066 0.0
V16194 n0_380_8409 n2_380_8409 0.0
V16195 n0_380_10569 n2_380_10569 0.0
V16196 n0_380_10602 n2_380_10602 0.0
V16197 n0_380_15105 n2_380_15105 0.0
V16198 n0_380_15138 n2_380_15138 0.0
V16199 n0_380_17298 n2_380_17298 0.0
V16200 n0_380_19641 n2_380_19641 0.0
V16201 n0_380_19674 n2_380_19674 0.0
V16202 n0_429_633 n2_429_633 0.0
V16203 n0_429_666 n2_429_666 0.0
V16204 n0_429_849 n2_429_849 0.0
V16205 n0_429_882 n2_429_882 0.0
V16206 n0_429_1065 n2_429_1065 0.0
V16207 n0_429_1098 n2_429_1098 0.0
V16208 n0_429_1281 n2_429_1281 0.0
V16209 n0_429_1314 n2_429_1314 0.0
V16210 n0_429_1497 n2_429_1497 0.0
V16211 n0_429_1530 n2_429_1530 0.0
V16212 n0_429_1713 n2_429_1713 0.0
V16213 n0_429_1746 n2_429_1746 0.0
V16214 n0_429_1929 n2_429_1929 0.0
V16215 n0_429_1962 n2_429_1962 0.0
V16216 n0_429_2145 n2_429_2145 0.0
V16217 n0_429_2178 n2_429_2178 0.0
V16218 n0_429_2361 n2_429_2361 0.0
V16219 n0_429_2394 n2_429_2394 0.0
V16220 n0_429_2577 n2_429_2577 0.0
V16221 n0_429_2610 n2_429_2610 0.0
V16222 n0_429_2826 n2_429_2826 0.0
V16223 n0_429_3009 n2_429_3009 0.0
V16224 n0_429_3042 n2_429_3042 0.0
V16225 n0_429_3225 n2_429_3225 0.0
V16226 n0_429_3258 n2_429_3258 0.0
V16227 n0_429_3441 n2_429_3441 0.0
V16228 n0_429_3474 n2_429_3474 0.0
V16229 n0_429_3657 n2_429_3657 0.0
V16230 n0_429_3690 n2_429_3690 0.0
V16231 n0_429_3873 n2_429_3873 0.0
V16232 n0_429_3906 n2_429_3906 0.0
V16233 n0_429_4089 n2_429_4089 0.0
V16234 n0_429_4122 n2_429_4122 0.0
V16235 n0_429_4305 n2_429_4305 0.0
V16236 n0_429_4338 n2_429_4338 0.0
V16237 n0_429_4375 n2_429_4375 0.0
V16238 n0_429_4521 n2_429_4521 0.0
V16239 n0_429_4554 n2_429_4554 0.0
V16240 n0_429_4737 n2_429_4737 0.0
V16241 n0_429_4770 n2_429_4770 0.0
V16242 n0_429_5169 n2_429_5169 0.0
V16243 n0_429_5202 n2_429_5202 0.0
V16244 n0_429_5385 n2_429_5385 0.0
V16245 n0_429_5418 n2_429_5418 0.0
V16246 n0_429_5601 n2_429_5601 0.0
V16247 n0_429_5634 n2_429_5634 0.0
V16248 n0_429_5817 n2_429_5817 0.0
V16249 n0_429_5850 n2_429_5850 0.0
V16250 n0_429_6033 n2_429_6033 0.0
V16251 n0_429_6066 n2_429_6066 0.0
V16252 n0_429_6249 n2_429_6249 0.0
V16253 n0_429_6282 n2_429_6282 0.0
V16254 n0_429_6465 n2_429_6465 0.0
V16255 n0_429_6498 n2_429_6498 0.0
V16256 n0_429_6681 n2_429_6681 0.0
V16257 n0_429_6714 n2_429_6714 0.0
V16258 n0_429_6897 n2_429_6897 0.0
V16259 n0_429_6930 n2_429_6930 0.0
V16260 n0_429_7113 n2_429_7113 0.0
V16261 n0_429_7329 n2_429_7329 0.0
V16262 n0_429_7362 n2_429_7362 0.0
V16263 n0_429_7545 n2_429_7545 0.0
V16264 n0_429_7578 n2_429_7578 0.0
V16265 n0_429_7761 n2_429_7761 0.0
V16266 n0_429_7794 n2_429_7794 0.0
V16267 n0_429_7977 n2_429_7977 0.0
V16268 n0_429_8010 n2_429_8010 0.0
V16269 n0_429_8193 n2_429_8193 0.0
V16270 n0_429_8226 n2_429_8226 0.0
V16271 n0_429_8409 n2_429_8409 0.0
V16272 n0_429_8442 n2_429_8442 0.0
V16273 n0_429_8625 n2_429_8625 0.0
V16274 n0_429_8658 n2_429_8658 0.0
V16275 n0_429_8841 n2_429_8841 0.0
V16276 n0_429_8874 n2_429_8874 0.0
V16277 n0_429_9057 n2_429_9057 0.0
V16278 n0_429_9090 n2_429_9090 0.0
V16279 n0_429_9273 n2_429_9273 0.0
V16280 n0_429_9306 n2_429_9306 0.0
V16281 n0_429_9705 n2_429_9705 0.0
V16282 n0_429_9738 n2_429_9738 0.0
V16283 n0_429_9921 n2_429_9921 0.0
V16284 n0_429_9954 n2_429_9954 0.0
V16285 n0_429_10137 n2_429_10137 0.0
V16286 n0_429_10170 n2_429_10170 0.0
V16287 n0_429_10353 n2_429_10353 0.0
V16288 n0_429_10386 n2_429_10386 0.0
V16289 n0_429_10569 n2_429_10569 0.0
V16290 n0_429_10602 n2_429_10602 0.0
V16291 n0_429_10785 n2_429_10785 0.0
V16292 n0_429_10818 n2_429_10818 0.0
V16293 n0_429_11001 n2_429_11001 0.0
V16294 n0_429_11034 n2_429_11034 0.0
V16295 n0_429_11217 n2_429_11217 0.0
V16296 n0_429_11250 n2_429_11250 0.0
V16297 n0_429_11433 n2_429_11433 0.0
V16298 n0_429_11466 n2_429_11466 0.0
V16299 n0_429_11865 n2_429_11865 0.0
V16300 n0_429_11898 n2_429_11898 0.0
V16301 n0_429_12081 n2_429_12081 0.0
V16302 n0_429_12114 n2_429_12114 0.0
V16303 n0_429_12297 n2_429_12297 0.0
V16304 n0_429_12330 n2_429_12330 0.0
V16305 n0_429_12513 n2_429_12513 0.0
V16306 n0_429_12546 n2_429_12546 0.0
V16307 n0_429_12729 n2_429_12729 0.0
V16308 n0_429_12762 n2_429_12762 0.0
V16309 n0_429_12945 n2_429_12945 0.0
V16310 n0_429_12978 n2_429_12978 0.0
V16311 n0_429_13161 n2_429_13161 0.0
V16312 n0_429_13194 n2_429_13194 0.0
V16313 n0_429_13377 n2_429_13377 0.0
V16314 n0_429_13410 n2_429_13410 0.0
V16315 n0_429_13593 n2_429_13593 0.0
V16316 n0_429_13626 n2_429_13626 0.0
V16317 n0_429_13663 n2_429_13663 0.0
V16318 n0_429_13809 n2_429_13809 0.0
V16319 n0_429_13842 n2_429_13842 0.0
V16320 n0_429_14241 n2_429_14241 0.0
V16321 n0_429_14274 n2_429_14274 0.0
V16322 n0_429_14457 n2_429_14457 0.0
V16323 n0_429_14490 n2_429_14490 0.0
V16324 n0_429_14673 n2_429_14673 0.0
V16325 n0_429_14706 n2_429_14706 0.0
V16326 n0_429_14889 n2_429_14889 0.0
V16327 n0_429_14922 n2_429_14922 0.0
V16328 n0_429_15105 n2_429_15105 0.0
V16329 n0_429_15138 n2_429_15138 0.0
V16330 n0_429_15321 n2_429_15321 0.0
V16331 n0_429_15354 n2_429_15354 0.0
V16332 n0_429_15537 n2_429_15537 0.0
V16333 n0_429_15570 n2_429_15570 0.0
V16334 n0_429_15753 n2_429_15753 0.0
V16335 n0_429_15786 n2_429_15786 0.0
V16336 n0_429_15969 n2_429_15969 0.0
V16337 n0_429_16002 n2_429_16002 0.0
V16338 n0_429_16401 n2_429_16401 0.0
V16339 n0_429_16434 n2_429_16434 0.0
V16340 n0_429_16617 n2_429_16617 0.0
V16341 n0_429_16650 n2_429_16650 0.0
V16342 n0_429_16833 n2_429_16833 0.0
V16343 n0_429_16866 n2_429_16866 0.0
V16344 n0_429_17049 n2_429_17049 0.0
V16345 n0_429_17082 n2_429_17082 0.0
V16346 n0_429_17265 n2_429_17265 0.0
V16347 n0_429_17298 n2_429_17298 0.0
V16348 n0_429_17481 n2_429_17481 0.0
V16349 n0_429_17514 n2_429_17514 0.0
V16350 n0_429_17697 n2_429_17697 0.0
V16351 n0_429_17730 n2_429_17730 0.0
V16352 n0_429_17913 n2_429_17913 0.0
V16353 n0_429_17946 n2_429_17946 0.0
V16354 n0_429_17960 n2_429_17960 0.0
V16355 n0_429_18129 n2_429_18129 0.0
V16356 n0_429_18162 n2_429_18162 0.0
V16357 n0_429_18345 n2_429_18345 0.0
V16358 n0_429_18594 n2_429_18594 0.0
V16359 n0_429_18777 n2_429_18777 0.0
V16360 n0_429_18810 n2_429_18810 0.0
V16361 n0_429_18993 n2_429_18993 0.0
V16362 n0_429_19026 n2_429_19026 0.0
V16363 n0_429_19040 n2_429_19040 0.0
V16364 n0_429_19209 n2_429_19209 0.0
V16365 n0_429_19242 n2_429_19242 0.0
V16366 n0_429_19256 n2_429_19256 0.0
V16367 n0_429_19425 n2_429_19425 0.0
V16368 n0_429_19458 n2_429_19458 0.0
V16369 n0_429_19472 n2_429_19472 0.0
V16370 n0_429_19641 n2_429_19641 0.0
V16371 n0_429_19674 n2_429_19674 0.0
V16372 n0_429_19857 n2_429_19857 0.0
V16373 n0_429_19890 n2_429_19890 0.0
V16374 n0_429_20073 n2_429_20073 0.0
V16375 n0_429_20106 n2_429_20106 0.0
V16376 n0_429_20289 n2_429_20289 0.0
V16377 n0_429_20322 n2_429_20322 0.0
V16378 n0_429_20505 n2_429_20505 0.0
V16379 n0_429_20538 n2_429_20538 0.0
V16380 n0_1366_201 n2_1366_201 0.0
V16381 n0_1366_234 n2_1366_234 0.0
V16382 n0_1366_417 n2_1366_417 0.0
V16383 n0_1366_450 n2_1366_450 0.0
V16384 n0_1366_633 n2_1366_633 0.0
V16385 n0_1366_666 n2_1366_666 0.0
V16386 n0_1366_849 n2_1366_849 0.0
V16387 n0_1366_882 n2_1366_882 0.0
V16388 n0_1366_1065 n2_1366_1065 0.0
V16389 n0_1366_1098 n2_1366_1098 0.0
V16390 n0_1366_1281 n2_1366_1281 0.0
V16391 n0_1366_1314 n2_1366_1314 0.0
V16392 n0_1366_1497 n2_1366_1497 0.0
V16393 n0_1366_1530 n2_1366_1530 0.0
V16394 n0_1366_1713 n2_1366_1713 0.0
V16395 n0_1366_1746 n2_1366_1746 0.0
V16396 n0_1366_1760 n2_1366_1760 0.0
V16397 n0_1366_1929 n2_1366_1929 0.0
V16398 n0_1366_1962 n2_1366_1962 0.0
V16399 n0_1366_2145 n2_1366_2145 0.0
V16400 n0_1366_2178 n2_1366_2178 0.0
V16401 n0_1366_2361 n2_1366_2361 0.0
V16402 n0_1366_2394 n2_1366_2394 0.0
V16403 n0_1366_2577 n2_1366_2577 0.0
V16404 n0_1366_2610 n2_1366_2610 0.0
V16405 n0_1366_2793 n2_1366_2793 0.0
V16406 n0_1366_2826 n2_1366_2826 0.0
V16407 n0_1366_3009 n2_1366_3009 0.0
V16408 n0_1366_3042 n2_1366_3042 0.0
V16409 n0_1366_3225 n2_1366_3225 0.0
V16410 n0_1366_3258 n2_1366_3258 0.0
V16411 n0_1366_3272 n2_1366_3272 0.0
V16412 n0_1366_3441 n2_1366_3441 0.0
V16413 n0_1366_3474 n2_1366_3474 0.0
V16414 n0_1366_3657 n2_1366_3657 0.0
V16415 n0_1366_3690 n2_1366_3690 0.0
V16416 n0_1366_3704 n2_1366_3704 0.0
V16417 n0_1366_3873 n2_1366_3873 0.0
V16418 n0_1366_3906 n2_1366_3906 0.0
V16419 n0_1366_3920 n2_1366_3920 0.0
V16420 n0_1366_4089 n2_1366_4089 0.0
V16421 n0_1366_4122 n2_1366_4122 0.0
V16422 n0_1366_4159 n2_1366_4159 0.0
V16423 n0_1366_4305 n2_1366_4305 0.0
V16424 n0_1366_4338 n2_1366_4338 0.0
V16425 n0_1366_4352 n2_1366_4352 0.0
V16426 n0_1366_4375 n2_1366_4375 0.0
V16427 n0_1366_4521 n2_1366_4521 0.0
V16428 n0_1366_4554 n2_1366_4554 0.0
V16429 n0_1366_4737 n2_1366_4737 0.0
V16430 n0_1366_4770 n2_1366_4770 0.0
V16431 n0_1366_4953 n2_1366_4953 0.0
V16432 n0_1366_4986 n2_1366_4986 0.0
V16433 n0_1366_5169 n2_1366_5169 0.0
V16434 n0_1366_5202 n2_1366_5202 0.0
V16435 n0_1366_5385 n2_1366_5385 0.0
V16436 n0_1366_5418 n2_1366_5418 0.0
V16437 n0_1366_5432 n2_1366_5432 0.0
V16438 n0_1366_5601 n2_1366_5601 0.0
V16439 n0_1366_5634 n2_1366_5634 0.0
V16440 n0_1366_5817 n2_1366_5817 0.0
V16441 n0_1366_5850 n2_1366_5850 0.0
V16442 n0_1366_6033 n2_1366_6033 0.0
V16443 n0_1366_6066 n2_1366_6066 0.0
V16444 n0_1366_6249 n2_1366_6249 0.0
V16445 n0_1366_6282 n2_1366_6282 0.0
V16446 n0_1366_6465 n2_1366_6465 0.0
V16447 n0_1366_6498 n2_1366_6498 0.0
V16448 n0_1366_6535 n2_1366_6535 0.0
V16449 n0_1366_6681 n2_1366_6681 0.0
V16450 n0_1366_6714 n2_1366_6714 0.0
V16451 n0_1366_6897 n2_1366_6897 0.0
V16452 n0_1366_6930 n2_1366_6930 0.0
V16453 n0_1366_7113 n2_1366_7113 0.0
V16454 n0_1366_7146 n2_1366_7146 0.0
V16455 n0_1366_7329 n2_1366_7329 0.0
V16456 n0_1366_7362 n2_1366_7362 0.0
V16457 n0_1366_7545 n2_1366_7545 0.0
V16458 n0_1366_7578 n2_1366_7578 0.0
V16459 n0_1366_7761 n2_1366_7761 0.0
V16460 n0_1366_7794 n2_1366_7794 0.0
V16461 n0_1366_7808 n2_1366_7808 0.0
V16462 n0_1366_7977 n2_1366_7977 0.0
V16463 n0_1366_8010 n2_1366_8010 0.0
V16464 n0_1366_8193 n2_1366_8193 0.0
V16465 n0_1366_8226 n2_1366_8226 0.0
V16466 n0_1366_8409 n2_1366_8409 0.0
V16467 n0_1366_8442 n2_1366_8442 0.0
V16468 n0_1366_8625 n2_1366_8625 0.0
V16469 n0_1366_8658 n2_1366_8658 0.0
V16470 n0_1366_8841 n2_1366_8841 0.0
V16471 n0_1366_8874 n2_1366_8874 0.0
V16472 n0_1366_8888 n2_1366_8888 0.0
V16473 n0_1366_8911 n2_1366_8911 0.0
V16474 n0_1366_9057 n2_1366_9057 0.0
V16475 n0_1366_9090 n2_1366_9090 0.0
V16476 n0_1366_9273 n2_1366_9273 0.0
V16477 n0_1366_9306 n2_1366_9306 0.0
V16478 n0_1366_9489 n2_1366_9489 0.0
V16479 n0_1366_9522 n2_1366_9522 0.0
V16480 n0_1366_9705 n2_1366_9705 0.0
V16481 n0_1366_9738 n2_1366_9738 0.0
V16482 n0_1366_9921 n2_1366_9921 0.0
V16483 n0_1366_9954 n2_1366_9954 0.0
V16484 n0_1366_9968 n2_1366_9968 0.0
V16485 n0_1366_10137 n2_1366_10137 0.0
V16486 n0_1366_10170 n2_1366_10170 0.0
V16487 n0_1366_10353 n2_1366_10353 0.0
V16488 n0_1366_10386 n2_1366_10386 0.0
V16489 n0_1366_10569 n2_1366_10569 0.0
V16490 n0_1366_10785 n2_1366_10785 0.0
V16491 n0_1366_10818 n2_1366_10818 0.0
V16492 n0_1366_11001 n2_1366_11001 0.0
V16493 n0_1366_11034 n2_1366_11034 0.0
V16494 n0_1366_11048 n2_1366_11048 0.0
V16495 n0_1366_11071 n2_1366_11071 0.0
V16496 n0_1366_11217 n2_1366_11217 0.0
V16497 n0_1366_11250 n2_1366_11250 0.0
V16498 n0_1366_11433 n2_1366_11433 0.0
V16499 n0_1366_11466 n2_1366_11466 0.0
V16500 n0_1366_11649 n2_1366_11649 0.0
V16501 n0_1366_11682 n2_1366_11682 0.0
V16502 n0_1366_11865 n2_1366_11865 0.0
V16503 n0_1366_11898 n2_1366_11898 0.0
V16504 n0_1366_12081 n2_1366_12081 0.0
V16505 n0_1366_12114 n2_1366_12114 0.0
V16506 n0_1366_12128 n2_1366_12128 0.0
V16507 n0_1366_12297 n2_1366_12297 0.0
V16508 n0_1366_12330 n2_1366_12330 0.0
V16509 n0_1366_12513 n2_1366_12513 0.0
V16510 n0_1366_12546 n2_1366_12546 0.0
V16511 n0_1366_12729 n2_1366_12729 0.0
V16512 n0_1366_12762 n2_1366_12762 0.0
V16513 n0_1366_12945 n2_1366_12945 0.0
V16514 n0_1366_12978 n2_1366_12978 0.0
V16515 n0_1366_13161 n2_1366_13161 0.0
V16516 n0_1366_13194 n2_1366_13194 0.0
V16517 n0_1366_13377 n2_1366_13377 0.0
V16518 n0_1366_13410 n2_1366_13410 0.0
V16519 n0_1366_13447 n2_1366_13447 0.0
V16520 n0_1366_13593 n2_1366_13593 0.0
V16521 n0_1366_13626 n2_1366_13626 0.0
V16522 n0_1366_13663 n2_1366_13663 0.0
V16523 n0_1366_13809 n2_1366_13809 0.0
V16524 n0_1366_13842 n2_1366_13842 0.0
V16525 n0_1366_14025 n2_1366_14025 0.0
V16526 n0_1366_14058 n2_1366_14058 0.0
V16527 n0_1366_14241 n2_1366_14241 0.0
V16528 n0_1366_14274 n2_1366_14274 0.0
V16529 n0_1366_14457 n2_1366_14457 0.0
V16530 n0_1366_14490 n2_1366_14490 0.0
V16531 n0_1366_14504 n2_1366_14504 0.0
V16532 n0_1366_14673 n2_1366_14673 0.0
V16533 n0_1366_14706 n2_1366_14706 0.0
V16534 n0_1366_14889 n2_1366_14889 0.0
V16535 n0_1366_14922 n2_1366_14922 0.0
V16536 n0_1366_15138 n2_1366_15138 0.0
V16537 n0_1366_15321 n2_1366_15321 0.0
V16538 n0_1366_15354 n2_1366_15354 0.0
V16539 n0_1366_15368 n2_1366_15368 0.0
V16540 n0_1366_15537 n2_1366_15537 0.0
V16541 n0_1366_15570 n2_1366_15570 0.0
V16542 n0_1366_15753 n2_1366_15753 0.0
V16543 n0_1366_15786 n2_1366_15786 0.0
V16544 n0_1366_15969 n2_1366_15969 0.0
V16545 n0_1366_16002 n2_1366_16002 0.0
V16546 n0_1366_16185 n2_1366_16185 0.0
V16547 n0_1366_16218 n2_1366_16218 0.0
V16548 n0_1366_16401 n2_1366_16401 0.0
V16549 n0_1366_16434 n2_1366_16434 0.0
V16550 n0_1366_16471 n2_1366_16471 0.0
V16551 n0_1366_16617 n2_1366_16617 0.0
V16552 n0_1366_16650 n2_1366_16650 0.0
V16553 n0_1366_16687 n2_1366_16687 0.0
V16554 n0_1366_16833 n2_1366_16833 0.0
V16555 n0_1366_16866 n2_1366_16866 0.0
V16556 n0_1366_16880 n2_1366_16880 0.0
V16557 n0_1366_17049 n2_1366_17049 0.0
V16558 n0_1366_17082 n2_1366_17082 0.0
V16559 n0_1366_17265 n2_1366_17265 0.0
V16560 n0_1366_17298 n2_1366_17298 0.0
V16561 n0_1366_17481 n2_1366_17481 0.0
V16562 n0_1366_17514 n2_1366_17514 0.0
V16563 n0_1366_17528 n2_1366_17528 0.0
V16564 n0_1366_17697 n2_1366_17697 0.0
V16565 n0_1366_17730 n2_1366_17730 0.0
V16566 n0_1366_17913 n2_1366_17913 0.0
V16567 n0_1366_17946 n2_1366_17946 0.0
V16568 n0_1366_17960 n2_1366_17960 0.0
V16569 n0_1366_18129 n2_1366_18129 0.0
V16570 n0_1366_18162 n2_1366_18162 0.0
V16571 n0_1366_18345 n2_1366_18345 0.0
V16572 n0_1366_18378 n2_1366_18378 0.0
V16573 n0_1366_18561 n2_1366_18561 0.0
V16574 n0_1366_18594 n2_1366_18594 0.0
V16575 n0_1366_18777 n2_1366_18777 0.0
V16576 n0_1366_18810 n2_1366_18810 0.0
V16577 n0_1366_18993 n2_1366_18993 0.0
V16578 n0_1366_19026 n2_1366_19026 0.0
V16579 n0_1366_19040 n2_1366_19040 0.0
V16580 n0_1366_19209 n2_1366_19209 0.0
V16581 n0_1366_19242 n2_1366_19242 0.0
V16582 n0_1366_19256 n2_1366_19256 0.0
V16583 n0_1366_19425 n2_1366_19425 0.0
V16584 n0_1366_19458 n2_1366_19458 0.0
V16585 n0_1366_19472 n2_1366_19472 0.0
V16586 n0_1366_19641 n2_1366_19641 0.0
V16587 n0_1366_19674 n2_1366_19674 0.0
V16588 n0_1366_19857 n2_1366_19857 0.0
V16589 n0_1366_19890 n2_1366_19890 0.0
V16590 n0_1366_20073 n2_1366_20073 0.0
V16591 n0_1366_20106 n2_1366_20106 0.0
V16592 n0_1366_20289 n2_1366_20289 0.0
V16593 n0_1366_20322 n2_1366_20322 0.0
V16594 n0_1366_20505 n2_1366_20505 0.0
V16595 n0_1366_20538 n2_1366_20538 0.0
V16596 n0_1366_20754 n2_1366_20754 0.0
V16597 n0_1366_20937 n2_1366_20937 0.0
V16598 n0_1366_20970 n2_1366_20970 0.0
V16599 n0_1458_201 n2_1458_201 0.0
V16600 n0_1458_234 n2_1458_234 0.0
V16601 n0_1458_417 n2_1458_417 0.0
V16602 n0_1458_450 n2_1458_450 0.0
V16603 n0_1458_633 n2_1458_633 0.0
V16604 n0_1458_666 n2_1458_666 0.0
V16605 n0_1458_849 n2_1458_849 0.0
V16606 n0_1458_882 n2_1458_882 0.0
V16607 n0_1458_1065 n2_1458_1065 0.0
V16608 n0_1458_1098 n2_1458_1098 0.0
V16609 n0_1458_1281 n2_1458_1281 0.0
V16610 n0_1458_1314 n2_1458_1314 0.0
V16611 n0_1458_1497 n2_1458_1497 0.0
V16612 n0_1458_19857 n2_1458_19857 0.0
V16613 n0_1458_19890 n2_1458_19890 0.0
V16614 n0_1458_20073 n2_1458_20073 0.0
V16615 n0_1458_20106 n2_1458_20106 0.0
V16616 n0_1458_20289 n2_1458_20289 0.0
V16617 n0_1458_20322 n2_1458_20322 0.0
V16618 n0_1458_20505 n2_1458_20505 0.0
V16619 n0_1458_20538 n2_1458_20538 0.0
V16620 n0_1458_20721 n2_1458_20721 0.0
V16621 n0_1458_20754 n2_1458_20754 0.0
V16622 n0_1458_20937 n2_1458_20937 0.0
V16623 n0_1458_20970 n2_1458_20970 0.0
V16624 n0_1505_417 n2_1505_417 0.0
V16625 n0_1505_450 n2_1505_450 0.0
V16626 n0_1505_3873 n2_1505_3873 0.0
V16627 n0_1505_3906 n2_1505_3906 0.0
V16628 n0_1505_3920 n2_1505_3920 0.0
V16629 n0_1505_6033 n2_1505_6033 0.0
V16630 n0_1505_6066 n2_1505_6066 0.0
V16631 n0_1505_8409 n2_1505_8409 0.0
V16632 n0_1505_10569 n2_1505_10569 0.0
V16633 n0_1505_10602 n2_1505_10602 0.0
V16634 n0_1505_15105 n2_1505_15105 0.0
V16635 n0_1505_15138 n2_1505_15138 0.0
V16636 n0_1505_17298 n2_1505_17298 0.0
V16637 n0_1505_20721 n2_1505_20721 0.0
V16638 n0_1505_20754 n2_1505_20754 0.0
V16639 n0_1554_201 n2_1554_201 0.0
V16640 n0_1554_234 n2_1554_234 0.0
V16641 n0_1554_417 n2_1554_417 0.0
V16642 n0_1554_450 n2_1554_450 0.0
V16643 n0_1554_633 n2_1554_633 0.0
V16644 n0_1554_666 n2_1554_666 0.0
V16645 n0_1554_849 n2_1554_849 0.0
V16646 n0_1554_882 n2_1554_882 0.0
V16647 n0_1554_1065 n2_1554_1065 0.0
V16648 n0_1554_1098 n2_1554_1098 0.0
V16649 n0_1554_1281 n2_1554_1281 0.0
V16650 n0_1554_1314 n2_1554_1314 0.0
V16651 n0_1554_1497 n2_1554_1497 0.0
V16652 n0_1554_1713 n2_1554_1713 0.0
V16653 n0_1554_1746 n2_1554_1746 0.0
V16654 n0_1554_1760 n2_1554_1760 0.0
V16655 n0_1554_1929 n2_1554_1929 0.0
V16656 n0_1554_1962 n2_1554_1962 0.0
V16657 n0_1554_2145 n2_1554_2145 0.0
V16658 n0_1554_2178 n2_1554_2178 0.0
V16659 n0_1554_2361 n2_1554_2361 0.0
V16660 n0_1554_2394 n2_1554_2394 0.0
V16661 n0_1554_2577 n2_1554_2577 0.0
V16662 n0_1554_2610 n2_1554_2610 0.0
V16663 n0_1554_2826 n2_1554_2826 0.0
V16664 n0_1554_3009 n2_1554_3009 0.0
V16665 n0_1554_3042 n2_1554_3042 0.0
V16666 n0_1554_3225 n2_1554_3225 0.0
V16667 n0_1554_3258 n2_1554_3258 0.0
V16668 n0_1554_3272 n2_1554_3272 0.0
V16669 n0_1554_3441 n2_1554_3441 0.0
V16670 n0_1554_3474 n2_1554_3474 0.0
V16671 n0_1554_3657 n2_1554_3657 0.0
V16672 n0_1554_3690 n2_1554_3690 0.0
V16673 n0_1554_3704 n2_1554_3704 0.0
V16674 n0_1554_3873 n2_1554_3873 0.0
V16675 n0_1554_3906 n2_1554_3906 0.0
V16676 n0_1554_3920 n2_1554_3920 0.0
V16677 n0_1554_4089 n2_1554_4089 0.0
V16678 n0_1554_4122 n2_1554_4122 0.0
V16679 n0_1554_4159 n2_1554_4159 0.0
V16680 n0_1554_4305 n2_1554_4305 0.0
V16681 n0_1554_4338 n2_1554_4338 0.0
V16682 n0_1554_4352 n2_1554_4352 0.0
V16683 n0_1554_4375 n2_1554_4375 0.0
V16684 n0_1554_4521 n2_1554_4521 0.0
V16685 n0_1554_4554 n2_1554_4554 0.0
V16686 n0_1554_4737 n2_1554_4737 0.0
V16687 n0_1554_4770 n2_1554_4770 0.0
V16688 n0_1554_5169 n2_1554_5169 0.0
V16689 n0_1554_5202 n2_1554_5202 0.0
V16690 n0_1554_5385 n2_1554_5385 0.0
V16691 n0_1554_5418 n2_1554_5418 0.0
V16692 n0_1554_5432 n2_1554_5432 0.0
V16693 n0_1554_5534 n2_1554_5534 0.0
V16694 n0_1554_5601 n2_1554_5601 0.0
V16695 n0_1554_5634 n2_1554_5634 0.0
V16696 n0_1554_5817 n2_1554_5817 0.0
V16697 n0_1554_5850 n2_1554_5850 0.0
V16698 n0_1554_6033 n2_1554_6033 0.0
V16699 n0_1554_6066 n2_1554_6066 0.0
V16700 n0_1554_6249 n2_1554_6249 0.0
V16701 n0_1554_6282 n2_1554_6282 0.0
V16702 n0_1554_6465 n2_1554_6465 0.0
V16703 n0_1554_6498 n2_1554_6498 0.0
V16704 n0_1554_6535 n2_1554_6535 0.0
V16705 n0_1554_6681 n2_1554_6681 0.0
V16706 n0_1554_6714 n2_1554_6714 0.0
V16707 n0_1554_6897 n2_1554_6897 0.0
V16708 n0_1554_6930 n2_1554_6930 0.0
V16709 n0_1554_7113 n2_1554_7113 0.0
V16710 n0_1554_7329 n2_1554_7329 0.0
V16711 n0_1554_7362 n2_1554_7362 0.0
V16712 n0_1554_7545 n2_1554_7545 0.0
V16713 n0_1554_7578 n2_1554_7578 0.0
V16714 n0_1554_7761 n2_1554_7761 0.0
V16715 n0_1554_7794 n2_1554_7794 0.0
V16716 n0_1554_7808 n2_1554_7808 0.0
V16717 n0_1554_7977 n2_1554_7977 0.0
V16718 n0_1554_8010 n2_1554_8010 0.0
V16719 n0_1554_8193 n2_1554_8193 0.0
V16720 n0_1554_8226 n2_1554_8226 0.0
V16721 n0_1554_8409 n2_1554_8409 0.0
V16722 n0_1554_8442 n2_1554_8442 0.0
V16723 n0_1554_8625 n2_1554_8625 0.0
V16724 n0_1554_8658 n2_1554_8658 0.0
V16725 n0_1554_8841 n2_1554_8841 0.0
V16726 n0_1554_8874 n2_1554_8874 0.0
V16727 n0_1554_8888 n2_1554_8888 0.0
V16728 n0_1554_8911 n2_1554_8911 0.0
V16729 n0_1554_9057 n2_1554_9057 0.0
V16730 n0_1554_9090 n2_1554_9090 0.0
V16731 n0_1554_9273 n2_1554_9273 0.0
V16732 n0_1554_9306 n2_1554_9306 0.0
V16733 n0_1554_9705 n2_1554_9705 0.0
V16734 n0_1554_9738 n2_1554_9738 0.0
V16735 n0_1554_9921 n2_1554_9921 0.0
V16736 n0_1554_9954 n2_1554_9954 0.0
V16737 n0_1554_9968 n2_1554_9968 0.0
V16738 n0_1554_10137 n2_1554_10137 0.0
V16739 n0_1554_10170 n2_1554_10170 0.0
V16740 n0_1554_10353 n2_1554_10353 0.0
V16741 n0_1554_10386 n2_1554_10386 0.0
V16742 n0_1554_10569 n2_1554_10569 0.0
V16743 n0_1554_10602 n2_1554_10602 0.0
V16744 n0_1554_10785 n2_1554_10785 0.0
V16745 n0_1554_10818 n2_1554_10818 0.0
V16746 n0_1554_11001 n2_1554_11001 0.0
V16747 n0_1554_11034 n2_1554_11034 0.0
V16748 n0_1554_11048 n2_1554_11048 0.0
V16749 n0_1554_11071 n2_1554_11071 0.0
V16750 n0_1554_11217 n2_1554_11217 0.0
V16751 n0_1554_11250 n2_1554_11250 0.0
V16752 n0_1554_11433 n2_1554_11433 0.0
V16753 n0_1554_11466 n2_1554_11466 0.0
V16754 n0_1554_11865 n2_1554_11865 0.0
V16755 n0_1554_11898 n2_1554_11898 0.0
V16756 n0_1554_12081 n2_1554_12081 0.0
V16757 n0_1554_12114 n2_1554_12114 0.0
V16758 n0_1554_12128 n2_1554_12128 0.0
V16759 n0_1554_12297 n2_1554_12297 0.0
V16760 n0_1554_12330 n2_1554_12330 0.0
V16761 n0_1554_12513 n2_1554_12513 0.0
V16762 n0_1554_12546 n2_1554_12546 0.0
V16763 n0_1554_12729 n2_1554_12729 0.0
V16764 n0_1554_12762 n2_1554_12762 0.0
V16765 n0_1554_12945 n2_1554_12945 0.0
V16766 n0_1554_12978 n2_1554_12978 0.0
V16767 n0_1554_13161 n2_1554_13161 0.0
V16768 n0_1554_13194 n2_1554_13194 0.0
V16769 n0_1554_13377 n2_1554_13377 0.0
V16770 n0_1554_13410 n2_1554_13410 0.0
V16771 n0_1554_13447 n2_1554_13447 0.0
V16772 n0_1554_13593 n2_1554_13593 0.0
V16773 n0_1554_13626 n2_1554_13626 0.0
V16774 n0_1554_13663 n2_1554_13663 0.0
V16775 n0_1554_13809 n2_1554_13809 0.0
V16776 n0_1554_13842 n2_1554_13842 0.0
V16777 n0_1554_14241 n2_1554_14241 0.0
V16778 n0_1554_14274 n2_1554_14274 0.0
V16779 n0_1554_14457 n2_1554_14457 0.0
V16780 n0_1554_14490 n2_1554_14490 0.0
V16781 n0_1554_14504 n2_1554_14504 0.0
V16782 n0_1554_14673 n2_1554_14673 0.0
V16783 n0_1554_14706 n2_1554_14706 0.0
V16784 n0_1554_14889 n2_1554_14889 0.0
V16785 n0_1554_14922 n2_1554_14922 0.0
V16786 n0_1554_15105 n2_1554_15105 0.0
V16787 n0_1554_15138 n2_1554_15138 0.0
V16788 n0_1554_15321 n2_1554_15321 0.0
V16789 n0_1554_15354 n2_1554_15354 0.0
V16790 n0_1554_15368 n2_1554_15368 0.0
V16791 n0_1554_15537 n2_1554_15537 0.0
V16792 n0_1554_15570 n2_1554_15570 0.0
V16793 n0_1554_15753 n2_1554_15753 0.0
V16794 n0_1554_15786 n2_1554_15786 0.0
V16795 n0_1554_15969 n2_1554_15969 0.0
V16796 n0_1554_16002 n2_1554_16002 0.0
V16797 n0_1554_16401 n2_1554_16401 0.0
V16798 n0_1554_16434 n2_1554_16434 0.0
V16799 n0_1554_16471 n2_1554_16471 0.0
V16800 n0_1554_16617 n2_1554_16617 0.0
V16801 n0_1554_16650 n2_1554_16650 0.0
V16802 n0_1554_16687 n2_1554_16687 0.0
V16803 n0_1554_16833 n2_1554_16833 0.0
V16804 n0_1554_16866 n2_1554_16866 0.0
V16805 n0_1554_16880 n2_1554_16880 0.0
V16806 n0_1554_17049 n2_1554_17049 0.0
V16807 n0_1554_17082 n2_1554_17082 0.0
V16808 n0_1554_17265 n2_1554_17265 0.0
V16809 n0_1554_17298 n2_1554_17298 0.0
V16810 n0_1554_17481 n2_1554_17481 0.0
V16811 n0_1554_17514 n2_1554_17514 0.0
V16812 n0_1554_17528 n2_1554_17528 0.0
V16813 n0_1554_17697 n2_1554_17697 0.0
V16814 n0_1554_17730 n2_1554_17730 0.0
V16815 n0_1554_17913 n2_1554_17913 0.0
V16816 n0_1554_17946 n2_1554_17946 0.0
V16817 n0_1554_17960 n2_1554_17960 0.0
V16818 n0_1554_18129 n2_1554_18129 0.0
V16819 n0_1554_18162 n2_1554_18162 0.0
V16820 n0_1554_18345 n2_1554_18345 0.0
V16821 n0_1554_18594 n2_1554_18594 0.0
V16822 n0_1554_18777 n2_1554_18777 0.0
V16823 n0_1554_18810 n2_1554_18810 0.0
V16824 n0_1554_18993 n2_1554_18993 0.0
V16825 n0_1554_19026 n2_1554_19026 0.0
V16826 n0_1554_19040 n2_1554_19040 0.0
V16827 n0_1554_19209 n2_1554_19209 0.0
V16828 n0_1554_19242 n2_1554_19242 0.0
V16829 n0_1554_19256 n2_1554_19256 0.0
V16830 n0_1554_19425 n2_1554_19425 0.0
V16831 n0_1554_19458 n2_1554_19458 0.0
V16832 n0_1554_19472 n2_1554_19472 0.0
V16833 n0_1554_19857 n2_1554_19857 0.0
V16834 n0_1554_19890 n2_1554_19890 0.0
V16835 n0_1554_20073 n2_1554_20073 0.0
V16836 n0_1554_20106 n2_1554_20106 0.0
V16837 n0_1554_20289 n2_1554_20289 0.0
V16838 n0_1554_20322 n2_1554_20322 0.0
V16839 n0_1554_20505 n2_1554_20505 0.0
V16840 n0_1554_20538 n2_1554_20538 0.0
V16841 n0_1554_20721 n2_1554_20721 0.0
V16842 n0_1554_20754 n2_1554_20754 0.0
V16843 n0_1554_20937 n2_1554_20937 0.0
V16844 n0_1554_20970 n2_1554_20970 0.0
V16845 n0_1646_201 n2_1646_201 0.0
V16846 n0_1646_234 n2_1646_234 0.0
V16847 n0_1646_417 n2_1646_417 0.0
V16848 n0_1646_450 n2_1646_450 0.0
V16849 n0_1646_633 n2_1646_633 0.0
V16850 n0_1646_666 n2_1646_666 0.0
V16851 n0_1646_849 n2_1646_849 0.0
V16852 n0_1646_882 n2_1646_882 0.0
V16853 n0_1646_1065 n2_1646_1065 0.0
V16854 n0_1646_1098 n2_1646_1098 0.0
V16855 n0_1646_1281 n2_1646_1281 0.0
V16856 n0_1646_1314 n2_1646_1314 0.0
V16857 n0_1646_1497 n2_1646_1497 0.0
V16858 n0_1646_1530 n2_1646_1530 0.0
V16859 n0_1646_19641 n2_1646_19641 0.0
V16860 n0_1646_19674 n2_1646_19674 0.0
V16861 n0_1646_19857 n2_1646_19857 0.0
V16862 n0_1646_19890 n2_1646_19890 0.0
V16863 n0_1646_20073 n2_1646_20073 0.0
V16864 n0_1646_20106 n2_1646_20106 0.0
V16865 n0_1646_20289 n2_1646_20289 0.0
V16866 n0_1646_20322 n2_1646_20322 0.0
V16867 n0_1646_20505 n2_1646_20505 0.0
V16868 n0_1646_20538 n2_1646_20538 0.0
V16869 n0_1646_20754 n2_1646_20754 0.0
V16870 n0_1646_20937 n2_1646_20937 0.0
V16871 n0_1646_20970 n2_1646_20970 0.0
V16872 n0_2491_2793 n2_2491_2793 0.0
V16873 n0_2491_2826 n2_2491_2826 0.0
V16874 n0_2491_3009 n2_2491_3009 0.0
V16875 n0_2491_3042 n2_2491_3042 0.0
V16876 n0_2491_3225 n2_2491_3225 0.0
V16877 n0_2491_3258 n2_2491_3258 0.0
V16878 n0_2491_3272 n2_2491_3272 0.0
V16879 n0_2491_3441 n2_2491_3441 0.0
V16880 n0_2491_3474 n2_2491_3474 0.0
V16881 n0_2491_3657 n2_2491_3657 0.0
V16882 n0_2491_3690 n2_2491_3690 0.0
V16883 n0_2491_3704 n2_2491_3704 0.0
V16884 n0_2491_3873 n2_2491_3873 0.0
V16885 n0_2491_3906 n2_2491_3906 0.0
V16886 n0_2491_3920 n2_2491_3920 0.0
V16887 n0_2491_4089 n2_2491_4089 0.0
V16888 n0_2491_4122 n2_2491_4122 0.0
V16889 n0_2491_4159 n2_2491_4159 0.0
V16890 n0_2491_4305 n2_2491_4305 0.0
V16891 n0_2491_4338 n2_2491_4338 0.0
V16892 n0_2491_4352 n2_2491_4352 0.0
V16893 n0_2491_4521 n2_2491_4521 0.0
V16894 n0_2491_4554 n2_2491_4554 0.0
V16895 n0_2491_4737 n2_2491_4737 0.0
V16896 n0_2491_4770 n2_2491_4770 0.0
V16897 n0_2491_4953 n2_2491_4953 0.0
V16898 n0_2491_4986 n2_2491_4986 0.0
V16899 n0_2491_5169 n2_2491_5169 0.0
V16900 n0_2491_5202 n2_2491_5202 0.0
V16901 n0_2491_5385 n2_2491_5385 0.0
V16902 n0_2491_5418 n2_2491_5418 0.0
V16903 n0_2491_5432 n2_2491_5432 0.0
V16904 n0_2491_5601 n2_2491_5601 0.0
V16905 n0_2491_5634 n2_2491_5634 0.0
V16906 n0_2491_5817 n2_2491_5817 0.0
V16907 n0_2491_5850 n2_2491_5850 0.0
V16908 n0_2491_6033 n2_2491_6033 0.0
V16909 n0_2491_6066 n2_2491_6066 0.0
V16910 n0_2491_6249 n2_2491_6249 0.0
V16911 n0_2491_6282 n2_2491_6282 0.0
V16912 n0_2491_6465 n2_2491_6465 0.0
V16913 n0_2491_6498 n2_2491_6498 0.0
V16914 n0_2491_6535 n2_2491_6535 0.0
V16915 n0_2491_6681 n2_2491_6681 0.0
V16916 n0_2491_6714 n2_2491_6714 0.0
V16917 n0_2491_6897 n2_2491_6897 0.0
V16918 n0_2491_6930 n2_2491_6930 0.0
V16919 n0_2491_7113 n2_2491_7113 0.0
V16920 n0_2491_7146 n2_2491_7146 0.0
V16921 n0_2491_7329 n2_2491_7329 0.0
V16922 n0_2491_7362 n2_2491_7362 0.0
V16923 n0_2491_7545 n2_2491_7545 0.0
V16924 n0_2491_7578 n2_2491_7578 0.0
V16925 n0_2491_7761 n2_2491_7761 0.0
V16926 n0_2491_7794 n2_2491_7794 0.0
V16927 n0_2491_7808 n2_2491_7808 0.0
V16928 n0_2491_7977 n2_2491_7977 0.0
V16929 n0_2491_8010 n2_2491_8010 0.0
V16930 n0_2491_8193 n2_2491_8193 0.0
V16931 n0_2491_8226 n2_2491_8226 0.0
V16932 n0_2491_8409 n2_2491_8409 0.0
V16933 n0_2491_8442 n2_2491_8442 0.0
V16934 n0_2491_8625 n2_2491_8625 0.0
V16935 n0_2491_8658 n2_2491_8658 0.0
V16936 n0_2491_8841 n2_2491_8841 0.0
V16937 n0_2491_8874 n2_2491_8874 0.0
V16938 n0_2491_8888 n2_2491_8888 0.0
V16939 n0_2491_8911 n2_2491_8911 0.0
V16940 n0_2491_9057 n2_2491_9057 0.0
V16941 n0_2491_9090 n2_2491_9090 0.0
V16942 n0_2491_9273 n2_2491_9273 0.0
V16943 n0_2491_9306 n2_2491_9306 0.0
V16944 n0_2491_9489 n2_2491_9489 0.0
V16945 n0_2491_9522 n2_2491_9522 0.0
V16946 n0_2491_9705 n2_2491_9705 0.0
V16947 n0_2491_9738 n2_2491_9738 0.0
V16948 n0_2491_9921 n2_2491_9921 0.0
V16949 n0_2491_9954 n2_2491_9954 0.0
V16950 n0_2491_9968 n2_2491_9968 0.0
V16951 n0_2491_10137 n2_2491_10137 0.0
V16952 n0_2491_10170 n2_2491_10170 0.0
V16953 n0_2491_10353 n2_2491_10353 0.0
V16954 n0_2491_10386 n2_2491_10386 0.0
V16955 n0_2491_10569 n2_2491_10569 0.0
V16956 n0_2491_10785 n2_2491_10785 0.0
V16957 n0_2491_10818 n2_2491_10818 0.0
V16958 n0_2491_11001 n2_2491_11001 0.0
V16959 n0_2491_11034 n2_2491_11034 0.0
V16960 n0_2491_11048 n2_2491_11048 0.0
V16961 n0_2491_11071 n2_2491_11071 0.0
V16962 n0_2491_11217 n2_2491_11217 0.0
V16963 n0_2491_11250 n2_2491_11250 0.0
V16964 n0_2491_11433 n2_2491_11433 0.0
V16965 n0_2491_11466 n2_2491_11466 0.0
V16966 n0_2491_11649 n2_2491_11649 0.0
V16967 n0_2491_11682 n2_2491_11682 0.0
V16968 n0_2491_11865 n2_2491_11865 0.0
V16969 n0_2491_11898 n2_2491_11898 0.0
V16970 n0_2491_12081 n2_2491_12081 0.0
V16971 n0_2491_12114 n2_2491_12114 0.0
V16972 n0_2491_12128 n2_2491_12128 0.0
V16973 n0_2491_12151 n2_2491_12151 0.0
V16974 n0_2491_12297 n2_2491_12297 0.0
V16975 n0_2491_12330 n2_2491_12330 0.0
V16976 n0_2491_12513 n2_2491_12513 0.0
V16977 n0_2491_12546 n2_2491_12546 0.0
V16978 n0_2491_12729 n2_2491_12729 0.0
V16979 n0_2491_12762 n2_2491_12762 0.0
V16980 n0_2491_12945 n2_2491_12945 0.0
V16981 n0_2491_12978 n2_2491_12978 0.0
V16982 n0_2491_13161 n2_2491_13161 0.0
V16983 n0_2491_13194 n2_2491_13194 0.0
V16984 n0_2491_13377 n2_2491_13377 0.0
V16985 n0_2491_13410 n2_2491_13410 0.0
V16986 n0_2491_13424 n2_2491_13424 0.0
V16987 n0_2491_13447 n2_2491_13447 0.0
V16988 n0_2491_13593 n2_2491_13593 0.0
V16989 n0_2491_13626 n2_2491_13626 0.0
V16990 n0_2491_13640 n2_2491_13640 0.0
V16991 n0_2491_13809 n2_2491_13809 0.0
V16992 n0_2491_13842 n2_2491_13842 0.0
V16993 n0_2491_13879 n2_2491_13879 0.0
V16994 n0_2491_14025 n2_2491_14025 0.0
V16995 n0_2491_14058 n2_2491_14058 0.0
V16996 n0_2491_14100 n2_2491_14100 0.0
V16997 n0_2491_14241 n2_2491_14241 0.0
V16998 n0_2491_14274 n2_2491_14274 0.0
V16999 n0_2491_14457 n2_2491_14457 0.0
V17000 n0_2491_14490 n2_2491_14490 0.0
V17001 n0_2491_14504 n2_2491_14504 0.0
V17002 n0_2491_14536 n2_2491_14536 0.0
V17003 n0_2491_14673 n2_2491_14673 0.0
V17004 n0_2491_14706 n2_2491_14706 0.0
V17005 n0_2491_14889 n2_2491_14889 0.0
V17006 n0_2491_14922 n2_2491_14922 0.0
V17007 n0_2491_15138 n2_2491_15138 0.0
V17008 n0_2491_15321 n2_2491_15321 0.0
V17009 n0_2491_15354 n2_2491_15354 0.0
V17010 n0_2491_15368 n2_2491_15368 0.0
V17011 n0_2491_15537 n2_2491_15537 0.0
V17012 n0_2491_15570 n2_2491_15570 0.0
V17013 n0_2491_15584 n2_2491_15584 0.0
V17014 n0_2491_15753 n2_2491_15753 0.0
V17015 n0_2491_15786 n2_2491_15786 0.0
V17016 n0_2491_15969 n2_2491_15969 0.0
V17017 n0_2491_16002 n2_2491_16002 0.0
V17018 n0_2491_16185 n2_2491_16185 0.0
V17019 n0_2491_16218 n2_2491_16218 0.0
V17020 n0_2491_16401 n2_2491_16401 0.0
V17021 n0_2491_16434 n2_2491_16434 0.0
V17022 n0_2491_16471 n2_2491_16471 0.0
V17023 n0_2491_16617 n2_2491_16617 0.0
V17024 n0_2491_16650 n2_2491_16650 0.0
V17025 n0_2491_16664 n2_2491_16664 0.0
V17026 n0_2491_16687 n2_2491_16687 0.0
V17027 n0_2491_16833 n2_2491_16833 0.0
V17028 n0_2491_16866 n2_2491_16866 0.0
V17029 n0_2491_16880 n2_2491_16880 0.0
V17030 n0_2491_17049 n2_2491_17049 0.0
V17031 n0_2491_17082 n2_2491_17082 0.0
V17032 n0_2491_17265 n2_2491_17265 0.0
V17033 n0_2491_17298 n2_2491_17298 0.0
V17034 n0_2491_17481 n2_2491_17481 0.0
V17035 n0_2491_17514 n2_2491_17514 0.0
V17036 n0_2491_17528 n2_2491_17528 0.0
V17037 n0_2491_17551 n2_2491_17551 0.0
V17038 n0_2491_17697 n2_2491_17697 0.0
V17039 n0_2491_17730 n2_2491_17730 0.0
V17040 n0_2491_17913 n2_2491_17913 0.0
V17041 n0_2491_17946 n2_2491_17946 0.0
V17042 n0_2491_17960 n2_2491_17960 0.0
V17043 n0_2491_18129 n2_2491_18129 0.0
V17044 n0_2491_18162 n2_2491_18162 0.0
V17045 n0_2491_18345 n2_2491_18345 0.0
V17046 n0_2491_18378 n2_2491_18378 0.0
V17047 n0_2630_3873 n2_2630_3873 0.0
V17048 n0_2630_3906 n2_2630_3906 0.0
V17049 n0_2630_3920 n2_2630_3920 0.0
V17050 n0_2630_6033 n2_2630_6033 0.0
V17051 n0_2630_6066 n2_2630_6066 0.0
V17052 n0_2630_8409 n2_2630_8409 0.0
V17053 n0_2630_10569 n2_2630_10569 0.0
V17054 n0_2630_10602 n2_2630_10602 0.0
V17055 n0_2630_15105 n2_2630_15105 0.0
V17056 n0_2630_15138 n2_2630_15138 0.0
V17057 n0_2630_17298 n2_2630_17298 0.0
V17058 n0_2679_2826 n2_2679_2826 0.0
V17059 n0_2679_3009 n2_2679_3009 0.0
V17060 n0_2679_3042 n2_2679_3042 0.0
V17061 n0_2679_3225 n2_2679_3225 0.0
V17062 n0_2679_3258 n2_2679_3258 0.0
V17063 n0_2679_3272 n2_2679_3272 0.0
V17064 n0_2679_3441 n2_2679_3441 0.0
V17065 n0_2679_3474 n2_2679_3474 0.0
V17066 n0_2679_3657 n2_2679_3657 0.0
V17067 n0_2679_3690 n2_2679_3690 0.0
V17068 n0_2679_3704 n2_2679_3704 0.0
V17069 n0_2679_3873 n2_2679_3873 0.0
V17070 n0_2679_3906 n2_2679_3906 0.0
V17071 n0_2679_3920 n2_2679_3920 0.0
V17072 n0_2679_4089 n2_2679_4089 0.0
V17073 n0_2679_4122 n2_2679_4122 0.0
V17074 n0_2679_4159 n2_2679_4159 0.0
V17075 n0_2679_4305 n2_2679_4305 0.0
V17076 n0_2679_4338 n2_2679_4338 0.0
V17077 n0_2679_4352 n2_2679_4352 0.0
V17078 n0_2679_4521 n2_2679_4521 0.0
V17079 n0_2679_4554 n2_2679_4554 0.0
V17080 n0_2679_4737 n2_2679_4737 0.0
V17081 n0_2679_4770 n2_2679_4770 0.0
V17082 n0_2679_5169 n2_2679_5169 0.0
V17083 n0_2679_5202 n2_2679_5202 0.0
V17084 n0_2679_5385 n2_2679_5385 0.0
V17085 n0_2679_5418 n2_2679_5418 0.0
V17086 n0_2679_5432 n2_2679_5432 0.0
V17087 n0_2679_5601 n2_2679_5601 0.0
V17088 n0_2679_5634 n2_2679_5634 0.0
V17089 n0_2679_5817 n2_2679_5817 0.0
V17090 n0_2679_5850 n2_2679_5850 0.0
V17091 n0_2679_6033 n2_2679_6033 0.0
V17092 n0_2679_6066 n2_2679_6066 0.0
V17093 n0_2679_6249 n2_2679_6249 0.0
V17094 n0_2679_6282 n2_2679_6282 0.0
V17095 n0_2679_6465 n2_2679_6465 0.0
V17096 n0_2679_6498 n2_2679_6498 0.0
V17097 n0_2679_6535 n2_2679_6535 0.0
V17098 n0_2679_6681 n2_2679_6681 0.0
V17099 n0_2679_6714 n2_2679_6714 0.0
V17100 n0_2679_6897 n2_2679_6897 0.0
V17101 n0_2679_6930 n2_2679_6930 0.0
V17102 n0_2679_7113 n2_2679_7113 0.0
V17103 n0_2679_7329 n2_2679_7329 0.0
V17104 n0_2679_7362 n2_2679_7362 0.0
V17105 n0_2679_7545 n2_2679_7545 0.0
V17106 n0_2679_7578 n2_2679_7578 0.0
V17107 n0_2679_7761 n2_2679_7761 0.0
V17108 n0_2679_7794 n2_2679_7794 0.0
V17109 n0_2679_7808 n2_2679_7808 0.0
V17110 n0_2679_7977 n2_2679_7977 0.0
V17111 n0_2679_8010 n2_2679_8010 0.0
V17112 n0_2679_8193 n2_2679_8193 0.0
V17113 n0_2679_8226 n2_2679_8226 0.0
V17114 n0_2679_8409 n2_2679_8409 0.0
V17115 n0_2679_8442 n2_2679_8442 0.0
V17116 n0_2679_8625 n2_2679_8625 0.0
V17117 n0_2679_8658 n2_2679_8658 0.0
V17118 n0_2679_8841 n2_2679_8841 0.0
V17119 n0_2679_8874 n2_2679_8874 0.0
V17120 n0_2679_8888 n2_2679_8888 0.0
V17121 n0_2679_8911 n2_2679_8911 0.0
V17122 n0_2679_9057 n2_2679_9057 0.0
V17123 n0_2679_9090 n2_2679_9090 0.0
V17124 n0_2679_9273 n2_2679_9273 0.0
V17125 n0_2679_9306 n2_2679_9306 0.0
V17126 n0_2679_9705 n2_2679_9705 0.0
V17127 n0_2679_9738 n2_2679_9738 0.0
V17128 n0_2679_9921 n2_2679_9921 0.0
V17129 n0_2679_9954 n2_2679_9954 0.0
V17130 n0_2679_9968 n2_2679_9968 0.0
V17131 n0_2679_10137 n2_2679_10137 0.0
V17132 n0_2679_10170 n2_2679_10170 0.0
V17133 n0_2679_10353 n2_2679_10353 0.0
V17134 n0_2679_10386 n2_2679_10386 0.0
V17135 n0_2679_10569 n2_2679_10569 0.0
V17136 n0_2679_10602 n2_2679_10602 0.0
V17137 n0_2679_10785 n2_2679_10785 0.0
V17138 n0_2679_10818 n2_2679_10818 0.0
V17139 n0_2679_11001 n2_2679_11001 0.0
V17140 n0_2679_11034 n2_2679_11034 0.0
V17141 n0_2679_11048 n2_2679_11048 0.0
V17142 n0_2679_11071 n2_2679_11071 0.0
V17143 n0_2679_11217 n2_2679_11217 0.0
V17144 n0_2679_11250 n2_2679_11250 0.0
V17145 n0_2679_11433 n2_2679_11433 0.0
V17146 n0_2679_11466 n2_2679_11466 0.0
V17147 n0_2679_11865 n2_2679_11865 0.0
V17148 n0_2679_11898 n2_2679_11898 0.0
V17149 n0_2679_12081 n2_2679_12081 0.0
V17150 n0_2679_12114 n2_2679_12114 0.0
V17151 n0_2679_12128 n2_2679_12128 0.0
V17152 n0_2679_12151 n2_2679_12151 0.0
V17153 n0_2679_12297 n2_2679_12297 0.0
V17154 n0_2679_12330 n2_2679_12330 0.0
V17155 n0_2679_12513 n2_2679_12513 0.0
V17156 n0_2679_12546 n2_2679_12546 0.0
V17157 n0_2679_12729 n2_2679_12729 0.0
V17158 n0_2679_12762 n2_2679_12762 0.0
V17159 n0_2679_12945 n2_2679_12945 0.0
V17160 n0_2679_12978 n2_2679_12978 0.0
V17161 n0_2679_13161 n2_2679_13161 0.0
V17162 n0_2679_13194 n2_2679_13194 0.0
V17163 n0_2679_13377 n2_2679_13377 0.0
V17164 n0_2679_13410 n2_2679_13410 0.0
V17165 n0_2679_13424 n2_2679_13424 0.0
V17166 n0_2679_13447 n2_2679_13447 0.0
V17167 n0_2679_13593 n2_2679_13593 0.0
V17168 n0_2679_13626 n2_2679_13626 0.0
V17169 n0_2679_13640 n2_2679_13640 0.0
V17170 n0_2679_13809 n2_2679_13809 0.0
V17171 n0_2679_13842 n2_2679_13842 0.0
V17172 n0_2679_14100 n2_2679_14100 0.0
V17173 n0_2679_14241 n2_2679_14241 0.0
V17174 n0_2679_14274 n2_2679_14274 0.0
V17175 n0_2679_14457 n2_2679_14457 0.0
V17176 n0_2679_14490 n2_2679_14490 0.0
V17177 n0_2679_14504 n2_2679_14504 0.0
V17178 n0_2679_14536 n2_2679_14536 0.0
V17179 n0_2679_14673 n2_2679_14673 0.0
V17180 n0_2679_14706 n2_2679_14706 0.0
V17181 n0_2679_14889 n2_2679_14889 0.0
V17182 n0_2679_14922 n2_2679_14922 0.0
V17183 n0_2679_15105 n2_2679_15105 0.0
V17184 n0_2679_15138 n2_2679_15138 0.0
V17185 n0_2679_15321 n2_2679_15321 0.0
V17186 n0_2679_15354 n2_2679_15354 0.0
V17187 n0_2679_15368 n2_2679_15368 0.0
V17188 n0_2679_15537 n2_2679_15537 0.0
V17189 n0_2679_15570 n2_2679_15570 0.0
V17190 n0_2679_15584 n2_2679_15584 0.0
V17191 n0_2679_15753 n2_2679_15753 0.0
V17192 n0_2679_15786 n2_2679_15786 0.0
V17193 n0_2679_15969 n2_2679_15969 0.0
V17194 n0_2679_16002 n2_2679_16002 0.0
V17195 n0_2679_16401 n2_2679_16401 0.0
V17196 n0_2679_16434 n2_2679_16434 0.0
V17197 n0_2679_16471 n2_2679_16471 0.0
V17198 n0_2679_16617 n2_2679_16617 0.0
V17199 n0_2679_16650 n2_2679_16650 0.0
V17200 n0_2679_16664 n2_2679_16664 0.0
V17201 n0_2679_16687 n2_2679_16687 0.0
V17202 n0_2679_16833 n2_2679_16833 0.0
V17203 n0_2679_16866 n2_2679_16866 0.0
V17204 n0_2679_16880 n2_2679_16880 0.0
V17205 n0_2679_17049 n2_2679_17049 0.0
V17206 n0_2679_17082 n2_2679_17082 0.0
V17207 n0_2679_17265 n2_2679_17265 0.0
V17208 n0_2679_17298 n2_2679_17298 0.0
V17209 n0_2679_17481 n2_2679_17481 0.0
V17210 n0_2679_17514 n2_2679_17514 0.0
V17211 n0_2679_17528 n2_2679_17528 0.0
V17212 n0_2679_17551 n2_2679_17551 0.0
V17213 n0_2679_17697 n2_2679_17697 0.0
V17214 n0_2679_17730 n2_2679_17730 0.0
V17215 n0_2679_17913 n2_2679_17913 0.0
V17216 n0_2679_17946 n2_2679_17946 0.0
V17217 n0_2679_17960 n2_2679_17960 0.0
V17218 n0_2679_18129 n2_2679_18129 0.0
V17219 n0_2679_18162 n2_2679_18162 0.0
V17220 n0_2679_18345 n2_2679_18345 0.0
V17221 n0_3616_201 n2_3616_201 0.0
V17222 n0_3616_234 n2_3616_234 0.0
V17223 n0_3616_356 n2_3616_356 0.0
V17224 n0_3616_417 n2_3616_417 0.0
V17225 n0_3616_450 n2_3616_450 0.0
V17226 n0_3616_633 n2_3616_633 0.0
V17227 n0_3616_666 n2_3616_666 0.0
V17228 n0_3616_788 n2_3616_788 0.0
V17229 n0_3616_849 n2_3616_849 0.0
V17230 n0_3616_882 n2_3616_882 0.0
V17231 n0_3616_1065 n2_3616_1065 0.0
V17232 n0_3616_1098 n2_3616_1098 0.0
V17233 n0_3616_1281 n2_3616_1281 0.0
V17234 n0_3616_1314 n2_3616_1314 0.0
V17235 n0_3616_1497 n2_3616_1497 0.0
V17236 n0_3616_1530 n2_3616_1530 0.0
V17237 n0_3616_1652 n2_3616_1652 0.0
V17238 n0_3616_1713 n2_3616_1713 0.0
V17239 n0_3616_1746 n2_3616_1746 0.0
V17240 n0_3616_1929 n2_3616_1929 0.0
V17241 n0_3616_1962 n2_3616_1962 0.0
V17242 n0_3616_1976 n2_3616_1976 0.0
V17243 n0_3616_2145 n2_3616_2145 0.0
V17244 n0_3616_2178 n2_3616_2178 0.0
V17245 n0_3616_2361 n2_3616_2361 0.0
V17246 n0_3616_2394 n2_3616_2394 0.0
V17247 n0_3616_2577 n2_3616_2577 0.0
V17248 n0_3616_2610 n2_3616_2610 0.0
V17249 n0_3616_2793 n2_3616_2793 0.0
V17250 n0_3616_2826 n2_3616_2826 0.0
V17251 n0_3616_3009 n2_3616_3009 0.0
V17252 n0_3616_3042 n2_3616_3042 0.0
V17253 n0_3616_3225 n2_3616_3225 0.0
V17254 n0_3616_3258 n2_3616_3258 0.0
V17255 n0_3616_3441 n2_3616_3441 0.0
V17256 n0_3616_3474 n2_3616_3474 0.0
V17257 n0_3616_3657 n2_3616_3657 0.0
V17258 n0_3616_3690 n2_3616_3690 0.0
V17259 n0_3616_3704 n2_3616_3704 0.0
V17260 n0_3616_3873 n2_3616_3873 0.0
V17261 n0_3616_3906 n2_3616_3906 0.0
V17262 n0_3616_3920 n2_3616_3920 0.0
V17263 n0_3616_4089 n2_3616_4089 0.0
V17264 n0_3616_4122 n2_3616_4122 0.0
V17265 n0_3616_4136 n2_3616_4136 0.0
V17266 n0_3616_4159 n2_3616_4159 0.0
V17267 n0_3616_4305 n2_3616_4305 0.0
V17268 n0_3616_4338 n2_3616_4338 0.0
V17269 n0_3616_4352 n2_3616_4352 0.0
V17270 n0_3616_4375 n2_3616_4375 0.0
V17271 n0_3616_4521 n2_3616_4521 0.0
V17272 n0_3616_4554 n2_3616_4554 0.0
V17273 n0_3616_4737 n2_3616_4737 0.0
V17274 n0_3616_4770 n2_3616_4770 0.0
V17275 n0_3616_4953 n2_3616_4953 0.0
V17276 n0_3616_4986 n2_3616_4986 0.0
V17277 n0_3616_5169 n2_3616_5169 0.0
V17278 n0_3616_5202 n2_3616_5202 0.0
V17279 n0_3616_5385 n2_3616_5385 0.0
V17280 n0_3616_5418 n2_3616_5418 0.0
V17281 n0_3616_5432 n2_3616_5432 0.0
V17282 n0_3616_5601 n2_3616_5601 0.0
V17283 n0_3616_5634 n2_3616_5634 0.0
V17284 n0_3616_5817 n2_3616_5817 0.0
V17285 n0_3616_5850 n2_3616_5850 0.0
V17286 n0_3616_6033 n2_3616_6033 0.0
V17287 n0_3616_6066 n2_3616_6066 0.0
V17288 n0_3616_6249 n2_3616_6249 0.0
V17289 n0_3616_6282 n2_3616_6282 0.0
V17290 n0_3616_6465 n2_3616_6465 0.0
V17291 n0_3616_6498 n2_3616_6498 0.0
V17292 n0_3616_6535 n2_3616_6535 0.0
V17293 n0_3616_6681 n2_3616_6681 0.0
V17294 n0_3616_6714 n2_3616_6714 0.0
V17295 n0_3616_6897 n2_3616_6897 0.0
V17296 n0_3616_6930 n2_3616_6930 0.0
V17297 n0_3616_7113 n2_3616_7113 0.0
V17298 n0_3616_7146 n2_3616_7146 0.0
V17299 n0_3616_7329 n2_3616_7329 0.0
V17300 n0_3616_7362 n2_3616_7362 0.0
V17301 n0_3616_7545 n2_3616_7545 0.0
V17302 n0_3616_7578 n2_3616_7578 0.0
V17303 n0_3616_7761 n2_3616_7761 0.0
V17304 n0_3616_7794 n2_3616_7794 0.0
V17305 n0_3616_7808 n2_3616_7808 0.0
V17306 n0_3616_7977 n2_3616_7977 0.0
V17307 n0_3616_8010 n2_3616_8010 0.0
V17308 n0_3616_8193 n2_3616_8193 0.0
V17309 n0_3616_8226 n2_3616_8226 0.0
V17310 n0_3616_8409 n2_3616_8409 0.0
V17311 n0_3616_8442 n2_3616_8442 0.0
V17312 n0_3616_8625 n2_3616_8625 0.0
V17313 n0_3616_8658 n2_3616_8658 0.0
V17314 n0_3616_8841 n2_3616_8841 0.0
V17315 n0_3616_8874 n2_3616_8874 0.0
V17316 n0_3616_8888 n2_3616_8888 0.0
V17317 n0_3616_8911 n2_3616_8911 0.0
V17318 n0_3616_9057 n2_3616_9057 0.0
V17319 n0_3616_9090 n2_3616_9090 0.0
V17320 n0_3616_9273 n2_3616_9273 0.0
V17321 n0_3616_9306 n2_3616_9306 0.0
V17322 n0_3616_9489 n2_3616_9489 0.0
V17323 n0_3616_9522 n2_3616_9522 0.0
V17324 n0_3616_9705 n2_3616_9705 0.0
V17325 n0_3616_9738 n2_3616_9738 0.0
V17326 n0_3616_9921 n2_3616_9921 0.0
V17327 n0_3616_9954 n2_3616_9954 0.0
V17328 n0_3616_9968 n2_3616_9968 0.0
V17329 n0_3616_10137 n2_3616_10137 0.0
V17330 n0_3616_10170 n2_3616_10170 0.0
V17331 n0_3616_10353 n2_3616_10353 0.0
V17332 n0_3616_10386 n2_3616_10386 0.0
V17333 n0_3616_10569 n2_3616_10569 0.0
V17334 n0_3616_10785 n2_3616_10785 0.0
V17335 n0_3616_10818 n2_3616_10818 0.0
V17336 n0_3616_11001 n2_3616_11001 0.0
V17337 n0_3616_11034 n2_3616_11034 0.0
V17338 n0_3616_11048 n2_3616_11048 0.0
V17339 n0_3616_11217 n2_3616_11217 0.0
V17340 n0_3616_11250 n2_3616_11250 0.0
V17341 n0_3616_11433 n2_3616_11433 0.0
V17342 n0_3616_11466 n2_3616_11466 0.0
V17343 n0_3616_11649 n2_3616_11649 0.0
V17344 n0_3616_11682 n2_3616_11682 0.0
V17345 n0_3616_11865 n2_3616_11865 0.0
V17346 n0_3616_11898 n2_3616_11898 0.0
V17347 n0_3616_12081 n2_3616_12081 0.0
V17348 n0_3616_12114 n2_3616_12114 0.0
V17349 n0_3616_12128 n2_3616_12128 0.0
V17350 n0_3616_12151 n2_3616_12151 0.0
V17351 n0_3616_12297 n2_3616_12297 0.0
V17352 n0_3616_12330 n2_3616_12330 0.0
V17353 n0_3616_12513 n2_3616_12513 0.0
V17354 n0_3616_12546 n2_3616_12546 0.0
V17355 n0_3616_12729 n2_3616_12729 0.0
V17356 n0_3616_12762 n2_3616_12762 0.0
V17357 n0_3616_12945 n2_3616_12945 0.0
V17358 n0_3616_12978 n2_3616_12978 0.0
V17359 n0_3616_13161 n2_3616_13161 0.0
V17360 n0_3616_13194 n2_3616_13194 0.0
V17361 n0_3616_13377 n2_3616_13377 0.0
V17362 n0_3616_13410 n2_3616_13410 0.0
V17363 n0_3616_13424 n2_3616_13424 0.0
V17364 n0_3616_13593 n2_3616_13593 0.0
V17365 n0_3616_13626 n2_3616_13626 0.0
V17366 n0_3616_13640 n2_3616_13640 0.0
V17367 n0_3616_13809 n2_3616_13809 0.0
V17368 n0_3616_13842 n2_3616_13842 0.0
V17369 n0_3616_13879 n2_3616_13879 0.0
V17370 n0_3616_14025 n2_3616_14025 0.0
V17371 n0_3616_14058 n2_3616_14058 0.0
V17372 n0_3616_14100 n2_3616_14100 0.0
V17373 n0_3616_14241 n2_3616_14241 0.0
V17374 n0_3616_14274 n2_3616_14274 0.0
V17375 n0_3616_14457 n2_3616_14457 0.0
V17376 n0_3616_14490 n2_3616_14490 0.0
V17377 n0_3616_14536 n2_3616_14536 0.0
V17378 n0_3616_14673 n2_3616_14673 0.0
V17379 n0_3616_14706 n2_3616_14706 0.0
V17380 n0_3616_14889 n2_3616_14889 0.0
V17381 n0_3616_14922 n2_3616_14922 0.0
V17382 n0_3616_15138 n2_3616_15138 0.0
V17383 n0_3616_15321 n2_3616_15321 0.0
V17384 n0_3616_15354 n2_3616_15354 0.0
V17385 n0_3616_15368 n2_3616_15368 0.0
V17386 n0_3616_15537 n2_3616_15537 0.0
V17387 n0_3616_15570 n2_3616_15570 0.0
V17388 n0_3616_15584 n2_3616_15584 0.0
V17389 n0_3616_15753 n2_3616_15753 0.0
V17390 n0_3616_15786 n2_3616_15786 0.0
V17391 n0_3616_15969 n2_3616_15969 0.0
V17392 n0_3616_16002 n2_3616_16002 0.0
V17393 n0_3616_16185 n2_3616_16185 0.0
V17394 n0_3616_16218 n2_3616_16218 0.0
V17395 n0_3616_16401 n2_3616_16401 0.0
V17396 n0_3616_16434 n2_3616_16434 0.0
V17397 n0_3616_16471 n2_3616_16471 0.0
V17398 n0_3616_16617 n2_3616_16617 0.0
V17399 n0_3616_16650 n2_3616_16650 0.0
V17400 n0_3616_16664 n2_3616_16664 0.0
V17401 n0_3616_16833 n2_3616_16833 0.0
V17402 n0_3616_16866 n2_3616_16866 0.0
V17403 n0_3616_16880 n2_3616_16880 0.0
V17404 n0_3616_17049 n2_3616_17049 0.0
V17405 n0_3616_17082 n2_3616_17082 0.0
V17406 n0_3616_17265 n2_3616_17265 0.0
V17407 n0_3616_17298 n2_3616_17298 0.0
V17408 n0_3616_17481 n2_3616_17481 0.0
V17409 n0_3616_17514 n2_3616_17514 0.0
V17410 n0_3616_17528 n2_3616_17528 0.0
V17411 n0_3616_17551 n2_3616_17551 0.0
V17412 n0_3616_17697 n2_3616_17697 0.0
V17413 n0_3616_17730 n2_3616_17730 0.0
V17414 n0_3616_17913 n2_3616_17913 0.0
V17415 n0_3616_17946 n2_3616_17946 0.0
V17416 n0_3616_18129 n2_3616_18129 0.0
V17417 n0_3616_18162 n2_3616_18162 0.0
V17418 n0_3616_18345 n2_3616_18345 0.0
V17419 n0_3616_18378 n2_3616_18378 0.0
V17420 n0_3616_18561 n2_3616_18561 0.0
V17421 n0_3616_18594 n2_3616_18594 0.0
V17422 n0_3616_18777 n2_3616_18777 0.0
V17423 n0_3616_18810 n2_3616_18810 0.0
V17424 n0_3616_18993 n2_3616_18993 0.0
V17425 n0_3616_19026 n2_3616_19026 0.0
V17426 n0_3616_19209 n2_3616_19209 0.0
V17427 n0_3616_19242 n2_3616_19242 0.0
V17428 n0_3616_19425 n2_3616_19425 0.0
V17429 n0_3616_19458 n2_3616_19458 0.0
V17430 n0_3616_19641 n2_3616_19641 0.0
V17431 n0_3616_19674 n2_3616_19674 0.0
V17432 n0_3616_19857 n2_3616_19857 0.0
V17433 n0_3616_19890 n2_3616_19890 0.0
V17434 n0_3616_20073 n2_3616_20073 0.0
V17435 n0_3616_20106 n2_3616_20106 0.0
V17436 n0_3616_20289 n2_3616_20289 0.0
V17437 n0_3616_20322 n2_3616_20322 0.0
V17438 n0_3616_20505 n2_3616_20505 0.0
V17439 n0_3616_20538 n2_3616_20538 0.0
V17440 n0_3616_20754 n2_3616_20754 0.0
V17441 n0_3616_20937 n2_3616_20937 0.0
V17442 n0_3616_20970 n2_3616_20970 0.0
V17443 n0_3708_201 n2_3708_201 0.0
V17444 n0_3708_234 n2_3708_234 0.0
V17445 n0_3708_356 n2_3708_356 0.0
V17446 n0_3708_417 n2_3708_417 0.0
V17447 n0_3708_450 n2_3708_450 0.0
V17448 n0_3708_633 n2_3708_633 0.0
V17449 n0_3708_666 n2_3708_666 0.0
V17450 n0_3708_788 n2_3708_788 0.0
V17451 n0_3708_849 n2_3708_849 0.0
V17452 n0_3708_882 n2_3708_882 0.0
V17453 n0_3708_1065 n2_3708_1065 0.0
V17454 n0_3708_1098 n2_3708_1098 0.0
V17455 n0_3708_1281 n2_3708_1281 0.0
V17456 n0_3708_1314 n2_3708_1314 0.0
V17457 n0_3708_1497 n2_3708_1497 0.0
V17458 n0_3708_1530 n2_3708_1530 0.0
V17459 n0_3708_1652 n2_3708_1652 0.0
V17460 n0_3708_1713 n2_3708_1713 0.0
V17461 n0_3708_1746 n2_3708_1746 0.0
V17462 n0_3708_1929 n2_3708_1929 0.0
V17463 n0_3708_1962 n2_3708_1962 0.0
V17464 n0_3708_1976 n2_3708_1976 0.0
V17465 n0_3708_2145 n2_3708_2145 0.0
V17466 n0_3708_2178 n2_3708_2178 0.0
V17467 n0_3708_2361 n2_3708_2361 0.0
V17468 n0_3708_2394 n2_3708_2394 0.0
V17469 n0_3708_2577 n2_3708_2577 0.0
V17470 n0_3708_2610 n2_3708_2610 0.0
V17471 n0_3708_2793 n2_3708_2793 0.0
V17472 n0_3708_2826 n2_3708_2826 0.0
V17473 n0_3708_3009 n2_3708_3009 0.0
V17474 n0_3708_3042 n2_3708_3042 0.0
V17475 n0_3708_3225 n2_3708_3225 0.0
V17476 n0_3708_3258 n2_3708_3258 0.0
V17477 n0_3708_3441 n2_3708_3441 0.0
V17478 n0_3708_3474 n2_3708_3474 0.0
V17479 n0_3708_3657 n2_3708_3657 0.0
V17480 n0_3708_3690 n2_3708_3690 0.0
V17481 n0_3708_3704 n2_3708_3704 0.0
V17482 n0_3708_3873 n2_3708_3873 0.0
V17483 n0_3708_3906 n2_3708_3906 0.0
V17484 n0_3708_3920 n2_3708_3920 0.0
V17485 n0_3708_17265 n2_3708_17265 0.0
V17486 n0_3708_17298 n2_3708_17298 0.0
V17487 n0_3708_17335 n2_3708_17335 0.0
V17488 n0_3708_17481 n2_3708_17481 0.0
V17489 n0_3708_17514 n2_3708_17514 0.0
V17490 n0_3708_17528 n2_3708_17528 0.0
V17491 n0_3708_17551 n2_3708_17551 0.0
V17492 n0_3708_17697 n2_3708_17697 0.0
V17493 n0_3708_17730 n2_3708_17730 0.0
V17494 n0_3708_17913 n2_3708_17913 0.0
V17495 n0_3708_17946 n2_3708_17946 0.0
V17496 n0_3708_18129 n2_3708_18129 0.0
V17497 n0_3708_18162 n2_3708_18162 0.0
V17498 n0_3708_18345 n2_3708_18345 0.0
V17499 n0_3708_18378 n2_3708_18378 0.0
V17500 n0_3708_18561 n2_3708_18561 0.0
V17501 n0_3708_18594 n2_3708_18594 0.0
V17502 n0_3708_18777 n2_3708_18777 0.0
V17503 n0_3708_18810 n2_3708_18810 0.0
V17504 n0_3708_18993 n2_3708_18993 0.0
V17505 n0_3708_19026 n2_3708_19026 0.0
V17506 n0_3708_19209 n2_3708_19209 0.0
V17507 n0_3708_19242 n2_3708_19242 0.0
V17508 n0_3708_19425 n2_3708_19425 0.0
V17509 n0_3708_19458 n2_3708_19458 0.0
V17510 n0_3708_19641 n2_3708_19641 0.0
V17511 n0_3708_19674 n2_3708_19674 0.0
V17512 n0_3708_19857 n2_3708_19857 0.0
V17513 n0_3708_19890 n2_3708_19890 0.0
V17514 n0_3708_20073 n2_3708_20073 0.0
V17515 n0_3708_20106 n2_3708_20106 0.0
V17516 n0_3708_20289 n2_3708_20289 0.0
V17517 n0_3708_20322 n2_3708_20322 0.0
V17518 n0_3708_20505 n2_3708_20505 0.0
V17519 n0_3708_20538 n2_3708_20538 0.0
V17520 n0_3708_20721 n2_3708_20721 0.0
V17521 n0_3708_20754 n2_3708_20754 0.0
V17522 n0_3708_20937 n2_3708_20937 0.0
V17523 n0_3708_20970 n2_3708_20970 0.0
V17524 n0_3755_417 n2_3755_417 0.0
V17525 n0_3755_450 n2_3755_450 0.0
V17526 n0_3755_1530 n2_3755_1530 0.0
V17527 n0_3755_1652 n2_3755_1652 0.0
V17528 n0_3755_2793 n2_3755_2793 0.0
V17529 n0_3755_3873 n2_3755_3873 0.0
V17530 n0_3755_3906 n2_3755_3906 0.0
V17531 n0_3755_3920 n2_3755_3920 0.0
V17532 n0_3755_6033 n2_3755_6033 0.0
V17533 n0_3755_6066 n2_3755_6066 0.0
V17534 n0_3755_8409 n2_3755_8409 0.0
V17535 n0_3755_10569 n2_3755_10569 0.0
V17536 n0_3755_10602 n2_3755_10602 0.0
V17537 n0_3755_15105 n2_3755_15105 0.0
V17538 n0_3755_15138 n2_3755_15138 0.0
V17539 n0_3755_17298 n2_3755_17298 0.0
V17540 n0_3755_17335 n2_3755_17335 0.0
V17541 n0_3755_19641 n2_3755_19641 0.0
V17542 n0_3755_19674 n2_3755_19674 0.0
V17543 n0_3755_20721 n2_3755_20721 0.0
V17544 n0_3755_20754 n2_3755_20754 0.0
V17545 n0_3804_201 n2_3804_201 0.0
V17546 n0_3804_234 n2_3804_234 0.0
V17547 n0_3804_356 n2_3804_356 0.0
V17548 n0_3804_417 n2_3804_417 0.0
V17549 n0_3804_450 n2_3804_450 0.0
V17550 n0_3804_633 n2_3804_633 0.0
V17551 n0_3804_666 n2_3804_666 0.0
V17552 n0_3804_788 n2_3804_788 0.0
V17553 n0_3804_849 n2_3804_849 0.0
V17554 n0_3804_882 n2_3804_882 0.0
V17555 n0_3804_1065 n2_3804_1065 0.0
V17556 n0_3804_1098 n2_3804_1098 0.0
V17557 n0_3804_1281 n2_3804_1281 0.0
V17558 n0_3804_1314 n2_3804_1314 0.0
V17559 n0_3804_1497 n2_3804_1497 0.0
V17560 n0_3804_1530 n2_3804_1530 0.0
V17561 n0_3804_1652 n2_3804_1652 0.0
V17562 n0_3804_1713 n2_3804_1713 0.0
V17563 n0_3804_1746 n2_3804_1746 0.0
V17564 n0_3804_1929 n2_3804_1929 0.0
V17565 n0_3804_1962 n2_3804_1962 0.0
V17566 n0_3804_1976 n2_3804_1976 0.0
V17567 n0_3804_2145 n2_3804_2145 0.0
V17568 n0_3804_2178 n2_3804_2178 0.0
V17569 n0_3804_2361 n2_3804_2361 0.0
V17570 n0_3804_2394 n2_3804_2394 0.0
V17571 n0_3804_2577 n2_3804_2577 0.0
V17572 n0_3804_2610 n2_3804_2610 0.0
V17573 n0_3804_2793 n2_3804_2793 0.0
V17574 n0_3804_2826 n2_3804_2826 0.0
V17575 n0_3804_3009 n2_3804_3009 0.0
V17576 n0_3804_3042 n2_3804_3042 0.0
V17577 n0_3804_3225 n2_3804_3225 0.0
V17578 n0_3804_3258 n2_3804_3258 0.0
V17579 n0_3804_3441 n2_3804_3441 0.0
V17580 n0_3804_3474 n2_3804_3474 0.0
V17581 n0_3804_3657 n2_3804_3657 0.0
V17582 n0_3804_3690 n2_3804_3690 0.0
V17583 n0_3804_3704 n2_3804_3704 0.0
V17584 n0_3804_3873 n2_3804_3873 0.0
V17585 n0_3804_3906 n2_3804_3906 0.0
V17586 n0_3804_3920 n2_3804_3920 0.0
V17587 n0_3804_4089 n2_3804_4089 0.0
V17588 n0_3804_4122 n2_3804_4122 0.0
V17589 n0_3804_4136 n2_3804_4136 0.0
V17590 n0_3804_4159 n2_3804_4159 0.0
V17591 n0_3804_4305 n2_3804_4305 0.0
V17592 n0_3804_4338 n2_3804_4338 0.0
V17593 n0_3804_4352 n2_3804_4352 0.0
V17594 n0_3804_4375 n2_3804_4375 0.0
V17595 n0_3804_4521 n2_3804_4521 0.0
V17596 n0_3804_4554 n2_3804_4554 0.0
V17597 n0_3804_4737 n2_3804_4737 0.0
V17598 n0_3804_4770 n2_3804_4770 0.0
V17599 n0_3804_5169 n2_3804_5169 0.0
V17600 n0_3804_5202 n2_3804_5202 0.0
V17601 n0_3804_5385 n2_3804_5385 0.0
V17602 n0_3804_5418 n2_3804_5418 0.0
V17603 n0_3804_5432 n2_3804_5432 0.0
V17604 n0_3804_5601 n2_3804_5601 0.0
V17605 n0_3804_5634 n2_3804_5634 0.0
V17606 n0_3804_5817 n2_3804_5817 0.0
V17607 n0_3804_5850 n2_3804_5850 0.0
V17608 n0_3804_6033 n2_3804_6033 0.0
V17609 n0_3804_6066 n2_3804_6066 0.0
V17610 n0_3804_6249 n2_3804_6249 0.0
V17611 n0_3804_6282 n2_3804_6282 0.0
V17612 n0_3804_6465 n2_3804_6465 0.0
V17613 n0_3804_6498 n2_3804_6498 0.0
V17614 n0_3804_6535 n2_3804_6535 0.0
V17615 n0_3804_6681 n2_3804_6681 0.0
V17616 n0_3804_6714 n2_3804_6714 0.0
V17617 n0_3804_6897 n2_3804_6897 0.0
V17618 n0_3804_6930 n2_3804_6930 0.0
V17619 n0_3804_7113 n2_3804_7113 0.0
V17620 n0_3804_7329 n2_3804_7329 0.0
V17621 n0_3804_7362 n2_3804_7362 0.0
V17622 n0_3804_7545 n2_3804_7545 0.0
V17623 n0_3804_7578 n2_3804_7578 0.0
V17624 n0_3804_7761 n2_3804_7761 0.0
V17625 n0_3804_7794 n2_3804_7794 0.0
V17626 n0_3804_7808 n2_3804_7808 0.0
V17627 n0_3804_7977 n2_3804_7977 0.0
V17628 n0_3804_8010 n2_3804_8010 0.0
V17629 n0_3804_8193 n2_3804_8193 0.0
V17630 n0_3804_8226 n2_3804_8226 0.0
V17631 n0_3804_8409 n2_3804_8409 0.0
V17632 n0_3804_8442 n2_3804_8442 0.0
V17633 n0_3804_8625 n2_3804_8625 0.0
V17634 n0_3804_8658 n2_3804_8658 0.0
V17635 n0_3804_8841 n2_3804_8841 0.0
V17636 n0_3804_8874 n2_3804_8874 0.0
V17637 n0_3804_8888 n2_3804_8888 0.0
V17638 n0_3804_8911 n2_3804_8911 0.0
V17639 n0_3804_9057 n2_3804_9057 0.0
V17640 n0_3804_9090 n2_3804_9090 0.0
V17641 n0_3804_9273 n2_3804_9273 0.0
V17642 n0_3804_9306 n2_3804_9306 0.0
V17643 n0_3804_9705 n2_3804_9705 0.0
V17644 n0_3804_9738 n2_3804_9738 0.0
V17645 n0_3804_9921 n2_3804_9921 0.0
V17646 n0_3804_9954 n2_3804_9954 0.0
V17647 n0_3804_9968 n2_3804_9968 0.0
V17648 n0_3804_10137 n2_3804_10137 0.0
V17649 n0_3804_10170 n2_3804_10170 0.0
V17650 n0_3804_10353 n2_3804_10353 0.0
V17651 n0_3804_10386 n2_3804_10386 0.0
V17652 n0_3804_10569 n2_3804_10569 0.0
V17653 n0_3804_10602 n2_3804_10602 0.0
V17654 n0_3804_10785 n2_3804_10785 0.0
V17655 n0_3804_10818 n2_3804_10818 0.0
V17656 n0_3804_11001 n2_3804_11001 0.0
V17657 n0_3804_11034 n2_3804_11034 0.0
V17658 n0_3804_11048 n2_3804_11048 0.0
V17659 n0_3804_11217 n2_3804_11217 0.0
V17660 n0_3804_11250 n2_3804_11250 0.0
V17661 n0_3804_11433 n2_3804_11433 0.0
V17662 n0_3804_11466 n2_3804_11466 0.0
V17663 n0_3804_11865 n2_3804_11865 0.0
V17664 n0_3804_11898 n2_3804_11898 0.0
V17665 n0_3804_12081 n2_3804_12081 0.0
V17666 n0_3804_12114 n2_3804_12114 0.0
V17667 n0_3804_12128 n2_3804_12128 0.0
V17668 n0_3804_12151 n2_3804_12151 0.0
V17669 n0_3804_12297 n2_3804_12297 0.0
V17670 n0_3804_12330 n2_3804_12330 0.0
V17671 n0_3804_12513 n2_3804_12513 0.0
V17672 n0_3804_12546 n2_3804_12546 0.0
V17673 n0_3804_12729 n2_3804_12729 0.0
V17674 n0_3804_12762 n2_3804_12762 0.0
V17675 n0_3804_12945 n2_3804_12945 0.0
V17676 n0_3804_12978 n2_3804_12978 0.0
V17677 n0_3804_13161 n2_3804_13161 0.0
V17678 n0_3804_13194 n2_3804_13194 0.0
V17679 n0_3804_13377 n2_3804_13377 0.0
V17680 n0_3804_13410 n2_3804_13410 0.0
V17681 n0_3804_13424 n2_3804_13424 0.0
V17682 n0_3804_13593 n2_3804_13593 0.0
V17683 n0_3804_13626 n2_3804_13626 0.0
V17684 n0_3804_13640 n2_3804_13640 0.0
V17685 n0_3804_13809 n2_3804_13809 0.0
V17686 n0_3804_13842 n2_3804_13842 0.0
V17687 n0_3804_14100 n2_3804_14100 0.0
V17688 n0_3804_14241 n2_3804_14241 0.0
V17689 n0_3804_14274 n2_3804_14274 0.0
V17690 n0_3804_14457 n2_3804_14457 0.0
V17691 n0_3804_14490 n2_3804_14490 0.0
V17692 n0_3804_14536 n2_3804_14536 0.0
V17693 n0_3804_14673 n2_3804_14673 0.0
V17694 n0_3804_14706 n2_3804_14706 0.0
V17695 n0_3804_14889 n2_3804_14889 0.0
V17696 n0_3804_14922 n2_3804_14922 0.0
V17697 n0_3804_15105 n2_3804_15105 0.0
V17698 n0_3804_15138 n2_3804_15138 0.0
V17699 n0_3804_15321 n2_3804_15321 0.0
V17700 n0_3804_15354 n2_3804_15354 0.0
V17701 n0_3804_15368 n2_3804_15368 0.0
V17702 n0_3804_15537 n2_3804_15537 0.0
V17703 n0_3804_15570 n2_3804_15570 0.0
V17704 n0_3804_15584 n2_3804_15584 0.0
V17705 n0_3804_15753 n2_3804_15753 0.0
V17706 n0_3804_15786 n2_3804_15786 0.0
V17707 n0_3804_15969 n2_3804_15969 0.0
V17708 n0_3804_16002 n2_3804_16002 0.0
V17709 n0_3804_16401 n2_3804_16401 0.0
V17710 n0_3804_16434 n2_3804_16434 0.0
V17711 n0_3804_16471 n2_3804_16471 0.0
V17712 n0_3804_16617 n2_3804_16617 0.0
V17713 n0_3804_16650 n2_3804_16650 0.0
V17714 n0_3804_16664 n2_3804_16664 0.0
V17715 n0_3804_16833 n2_3804_16833 0.0
V17716 n0_3804_16866 n2_3804_16866 0.0
V17717 n0_3804_16880 n2_3804_16880 0.0
V17718 n0_3804_17049 n2_3804_17049 0.0
V17719 n0_3804_17082 n2_3804_17082 0.0
V17720 n0_3804_17265 n2_3804_17265 0.0
V17721 n0_3804_17298 n2_3804_17298 0.0
V17722 n0_3804_17335 n2_3804_17335 0.0
V17723 n0_3804_17481 n2_3804_17481 0.0
V17724 n0_3804_17514 n2_3804_17514 0.0
V17725 n0_3804_17528 n2_3804_17528 0.0
V17726 n0_3804_17551 n2_3804_17551 0.0
V17727 n0_3804_17697 n2_3804_17697 0.0
V17728 n0_3804_17730 n2_3804_17730 0.0
V17729 n0_3804_17913 n2_3804_17913 0.0
V17730 n0_3804_17946 n2_3804_17946 0.0
V17731 n0_3804_18129 n2_3804_18129 0.0
V17732 n0_3804_18162 n2_3804_18162 0.0
V17733 n0_3804_18345 n2_3804_18345 0.0
V17734 n0_3804_18378 n2_3804_18378 0.0
V17735 n0_3804_18561 n2_3804_18561 0.0
V17736 n0_3804_18594 n2_3804_18594 0.0
V17737 n0_3804_18777 n2_3804_18777 0.0
V17738 n0_3804_18810 n2_3804_18810 0.0
V17739 n0_3804_18993 n2_3804_18993 0.0
V17740 n0_3804_19026 n2_3804_19026 0.0
V17741 n0_3804_19209 n2_3804_19209 0.0
V17742 n0_3804_19242 n2_3804_19242 0.0
V17743 n0_3804_19425 n2_3804_19425 0.0
V17744 n0_3804_19458 n2_3804_19458 0.0
V17745 n0_3804_19641 n2_3804_19641 0.0
V17746 n0_3804_19674 n2_3804_19674 0.0
V17747 n0_3804_19857 n2_3804_19857 0.0
V17748 n0_3804_19890 n2_3804_19890 0.0
V17749 n0_3804_20073 n2_3804_20073 0.0
V17750 n0_3804_20106 n2_3804_20106 0.0
V17751 n0_3804_20289 n2_3804_20289 0.0
V17752 n0_3804_20322 n2_3804_20322 0.0
V17753 n0_3804_20505 n2_3804_20505 0.0
V17754 n0_3804_20538 n2_3804_20538 0.0
V17755 n0_3804_20721 n2_3804_20721 0.0
V17756 n0_3804_20754 n2_3804_20754 0.0
V17757 n0_3804_20937 n2_3804_20937 0.0
V17758 n0_3804_20970 n2_3804_20970 0.0
V17759 n0_3896_201 n2_3896_201 0.0
V17760 n0_3896_234 n2_3896_234 0.0
V17761 n0_3896_356 n2_3896_356 0.0
V17762 n0_3896_417 n2_3896_417 0.0
V17763 n0_3896_450 n2_3896_450 0.0
V17764 n0_3896_633 n2_3896_633 0.0
V17765 n0_3896_666 n2_3896_666 0.0
V17766 n0_3896_788 n2_3896_788 0.0
V17767 n0_3896_849 n2_3896_849 0.0
V17768 n0_3896_882 n2_3896_882 0.0
V17769 n0_3896_1065 n2_3896_1065 0.0
V17770 n0_3896_1098 n2_3896_1098 0.0
V17771 n0_3896_1281 n2_3896_1281 0.0
V17772 n0_3896_1314 n2_3896_1314 0.0
V17773 n0_3896_1497 n2_3896_1497 0.0
V17774 n0_3896_1530 n2_3896_1530 0.0
V17775 n0_3896_1652 n2_3896_1652 0.0
V17776 n0_3896_1713 n2_3896_1713 0.0
V17777 n0_3896_1746 n2_3896_1746 0.0
V17778 n0_3896_1929 n2_3896_1929 0.0
V17779 n0_3896_1962 n2_3896_1962 0.0
V17780 n0_3896_1976 n2_3896_1976 0.0
V17781 n0_3896_2145 n2_3896_2145 0.0
V17782 n0_3896_2178 n2_3896_2178 0.0
V17783 n0_3896_2361 n2_3896_2361 0.0
V17784 n0_3896_2394 n2_3896_2394 0.0
V17785 n0_3896_2577 n2_3896_2577 0.0
V17786 n0_3896_2610 n2_3896_2610 0.0
V17787 n0_3896_2793 n2_3896_2793 0.0
V17788 n0_3896_2826 n2_3896_2826 0.0
V17789 n0_3896_3009 n2_3896_3009 0.0
V17790 n0_3896_3042 n2_3896_3042 0.0
V17791 n0_3896_3225 n2_3896_3225 0.0
V17792 n0_3896_3258 n2_3896_3258 0.0
V17793 n0_3896_3441 n2_3896_3441 0.0
V17794 n0_3896_3474 n2_3896_3474 0.0
V17795 n0_3896_3657 n2_3896_3657 0.0
V17796 n0_3896_3690 n2_3896_3690 0.0
V17797 n0_3896_3704 n2_3896_3704 0.0
V17798 n0_3896_17481 n2_3896_17481 0.0
V17799 n0_3896_17514 n2_3896_17514 0.0
V17800 n0_3896_17528 n2_3896_17528 0.0
V17801 n0_3896_17551 n2_3896_17551 0.0
V17802 n0_3896_17697 n2_3896_17697 0.0
V17803 n0_3896_17730 n2_3896_17730 0.0
V17804 n0_3896_17913 n2_3896_17913 0.0
V17805 n0_3896_17946 n2_3896_17946 0.0
V17806 n0_3896_18129 n2_3896_18129 0.0
V17807 n0_3896_18162 n2_3896_18162 0.0
V17808 n0_3896_18345 n2_3896_18345 0.0
V17809 n0_3896_18378 n2_3896_18378 0.0
V17810 n0_3896_18561 n2_3896_18561 0.0
V17811 n0_3896_18594 n2_3896_18594 0.0
V17812 n0_3896_18777 n2_3896_18777 0.0
V17813 n0_3896_18810 n2_3896_18810 0.0
V17814 n0_3896_18993 n2_3896_18993 0.0
V17815 n0_3896_19026 n2_3896_19026 0.0
V17816 n0_3896_19209 n2_3896_19209 0.0
V17817 n0_3896_19242 n2_3896_19242 0.0
V17818 n0_3896_19425 n2_3896_19425 0.0
V17819 n0_3896_19458 n2_3896_19458 0.0
V17820 n0_3896_19641 n2_3896_19641 0.0
V17821 n0_3896_19674 n2_3896_19674 0.0
V17822 n0_3896_19857 n2_3896_19857 0.0
V17823 n0_3896_19890 n2_3896_19890 0.0
V17824 n0_3896_20073 n2_3896_20073 0.0
V17825 n0_3896_20106 n2_3896_20106 0.0
V17826 n0_3896_20289 n2_3896_20289 0.0
V17827 n0_3896_20322 n2_3896_20322 0.0
V17828 n0_3896_20505 n2_3896_20505 0.0
V17829 n0_3896_20538 n2_3896_20538 0.0
V17830 n0_3896_20754 n2_3896_20754 0.0
V17831 n0_3896_20937 n2_3896_20937 0.0
V17832 n0_3896_20970 n2_3896_20970 0.0
V17833 n0_4741_5169 n2_4741_5169 0.0
V17834 n0_4741_5202 n2_4741_5202 0.0
V17835 n0_4741_5385 n2_4741_5385 0.0
V17836 n0_4741_5418 n2_4741_5418 0.0
V17837 n0_4741_5432 n2_4741_5432 0.0
V17838 n0_4741_5601 n2_4741_5601 0.0
V17839 n0_4741_5634 n2_4741_5634 0.0
V17840 n0_4741_5817 n2_4741_5817 0.0
V17841 n0_4741_5850 n2_4741_5850 0.0
V17842 n0_4741_6033 n2_4741_6033 0.0
V17843 n0_4741_6066 n2_4741_6066 0.0
V17844 n0_4741_6249 n2_4741_6249 0.0
V17845 n0_4741_6282 n2_4741_6282 0.0
V17846 n0_4741_6465 n2_4741_6465 0.0
V17847 n0_4741_6498 n2_4741_6498 0.0
V17848 n0_4741_6535 n2_4741_6535 0.0
V17849 n0_4741_6681 n2_4741_6681 0.0
V17850 n0_4741_6714 n2_4741_6714 0.0
V17851 n0_4741_6897 n2_4741_6897 0.0
V17852 n0_4741_6930 n2_4741_6930 0.0
V17853 n0_4741_7113 n2_4741_7113 0.0
V17854 n0_4741_7146 n2_4741_7146 0.0
V17855 n0_4741_7329 n2_4741_7329 0.0
V17856 n0_4741_7362 n2_4741_7362 0.0
V17857 n0_4741_7545 n2_4741_7545 0.0
V17858 n0_4741_7578 n2_4741_7578 0.0
V17859 n0_4741_7761 n2_4741_7761 0.0
V17860 n0_4741_7794 n2_4741_7794 0.0
V17861 n0_4741_7808 n2_4741_7808 0.0
V17862 n0_4741_7977 n2_4741_7977 0.0
V17863 n0_4741_8010 n2_4741_8010 0.0
V17864 n0_4741_8193 n2_4741_8193 0.0
V17865 n0_4741_8226 n2_4741_8226 0.0
V17866 n0_4741_8409 n2_4741_8409 0.0
V17867 n0_4741_8442 n2_4741_8442 0.0
V17868 n0_4741_8625 n2_4741_8625 0.0
V17869 n0_4741_8658 n2_4741_8658 0.0
V17870 n0_4741_8841 n2_4741_8841 0.0
V17871 n0_4741_8874 n2_4741_8874 0.0
V17872 n0_4741_8888 n2_4741_8888 0.0
V17873 n0_4741_8911 n2_4741_8911 0.0
V17874 n0_4741_9057 n2_4741_9057 0.0
V17875 n0_4741_9090 n2_4741_9090 0.0
V17876 n0_4741_9273 n2_4741_9273 0.0
V17877 n0_4741_9306 n2_4741_9306 0.0
V17878 n0_4741_9489 n2_4741_9489 0.0
V17879 n0_4741_9522 n2_4741_9522 0.0
V17880 n0_4741_9705 n2_4741_9705 0.0
V17881 n0_4741_9738 n2_4741_9738 0.0
V17882 n0_4741_9921 n2_4741_9921 0.0
V17883 n0_4741_9954 n2_4741_9954 0.0
V17884 n0_4741_9968 n2_4741_9968 0.0
V17885 n0_4741_10137 n2_4741_10137 0.0
V17886 n0_4741_10170 n2_4741_10170 0.0
V17887 n0_4741_10353 n2_4741_10353 0.0
V17888 n0_4741_10386 n2_4741_10386 0.0
V17889 n0_4741_10569 n2_4741_10569 0.0
V17890 n0_4741_10785 n2_4741_10785 0.0
V17891 n0_4741_10818 n2_4741_10818 0.0
V17892 n0_4741_11001 n2_4741_11001 0.0
V17893 n0_4741_11034 n2_4741_11034 0.0
V17894 n0_4741_11048 n2_4741_11048 0.0
V17895 n0_4741_11071 n2_4741_11071 0.0
V17896 n0_4741_11217 n2_4741_11217 0.0
V17897 n0_4741_11250 n2_4741_11250 0.0
V17898 n0_4741_11433 n2_4741_11433 0.0
V17899 n0_4741_11466 n2_4741_11466 0.0
V17900 n0_4741_11649 n2_4741_11649 0.0
V17901 n0_4741_11682 n2_4741_11682 0.0
V17902 n0_4741_11865 n2_4741_11865 0.0
V17903 n0_4741_11898 n2_4741_11898 0.0
V17904 n0_4741_12081 n2_4741_12081 0.0
V17905 n0_4741_12114 n2_4741_12114 0.0
V17906 n0_4741_12128 n2_4741_12128 0.0
V17907 n0_4741_12297 n2_4741_12297 0.0
V17908 n0_4741_12330 n2_4741_12330 0.0
V17909 n0_4741_12513 n2_4741_12513 0.0
V17910 n0_4741_12546 n2_4741_12546 0.0
V17911 n0_4741_12729 n2_4741_12729 0.0
V17912 n0_4741_12762 n2_4741_12762 0.0
V17913 n0_4741_12945 n2_4741_12945 0.0
V17914 n0_4741_12978 n2_4741_12978 0.0
V17915 n0_4741_13161 n2_4741_13161 0.0
V17916 n0_4741_13194 n2_4741_13194 0.0
V17917 n0_4741_13377 n2_4741_13377 0.0
V17918 n0_4741_13410 n2_4741_13410 0.0
V17919 n0_4741_13424 n2_4741_13424 0.0
V17920 n0_4741_13593 n2_4741_13593 0.0
V17921 n0_4741_13626 n2_4741_13626 0.0
V17922 n0_4741_13809 n2_4741_13809 0.0
V17923 n0_4741_13842 n2_4741_13842 0.0
V17924 n0_4741_13879 n2_4741_13879 0.0
V17925 n0_4741_14025 n2_4741_14025 0.0
V17926 n0_4741_14058 n2_4741_14058 0.0
V17927 n0_4741_14100 n2_4741_14100 0.0
V17928 n0_4741_14241 n2_4741_14241 0.0
V17929 n0_4741_14274 n2_4741_14274 0.0
V17930 n0_4741_14457 n2_4741_14457 0.0
V17931 n0_4741_14490 n2_4741_14490 0.0
V17932 n0_4741_14536 n2_4741_14536 0.0
V17933 n0_4741_14673 n2_4741_14673 0.0
V17934 n0_4741_14706 n2_4741_14706 0.0
V17935 n0_4741_14889 n2_4741_14889 0.0
V17936 n0_4741_14922 n2_4741_14922 0.0
V17937 n0_4741_15138 n2_4741_15138 0.0
V17938 n0_4741_15321 n2_4741_15321 0.0
V17939 n0_4741_15354 n2_4741_15354 0.0
V17940 n0_4741_15368 n2_4741_15368 0.0
V17941 n0_4741_15537 n2_4741_15537 0.0
V17942 n0_4741_15570 n2_4741_15570 0.0
V17943 n0_4741_15584 n2_4741_15584 0.0
V17944 n0_4741_15753 n2_4741_15753 0.0
V17945 n0_4741_15786 n2_4741_15786 0.0
V17946 n0_4741_15969 n2_4741_15969 0.0
V17947 n0_4741_16002 n2_4741_16002 0.0
V17948 n0_4741_16016 n2_4741_16016 0.0
V17949 n0_4741_16185 n2_4741_16185 0.0
V17950 n0_4880_6033 n2_4880_6033 0.0
V17951 n0_4880_6066 n2_4880_6066 0.0
V17952 n0_4880_8409 n2_4880_8409 0.0
V17953 n0_4880_10569 n2_4880_10569 0.0
V17954 n0_4880_10602 n2_4880_10602 0.0
V17955 n0_4880_15105 n2_4880_15105 0.0
V17956 n0_4880_15138 n2_4880_15138 0.0
V17957 n0_4929_5169 n2_4929_5169 0.0
V17958 n0_4929_5202 n2_4929_5202 0.0
V17959 n0_4929_5385 n2_4929_5385 0.0
V17960 n0_4929_5418 n2_4929_5418 0.0
V17961 n0_4929_5432 n2_4929_5432 0.0
V17962 n0_4929_5601 n2_4929_5601 0.0
V17963 n0_4929_5634 n2_4929_5634 0.0
V17964 n0_4929_5817 n2_4929_5817 0.0
V17965 n0_4929_5850 n2_4929_5850 0.0
V17966 n0_4929_6033 n2_4929_6033 0.0
V17967 n0_4929_6066 n2_4929_6066 0.0
V17968 n0_4929_6249 n2_4929_6249 0.0
V17969 n0_4929_6282 n2_4929_6282 0.0
V17970 n0_4929_6465 n2_4929_6465 0.0
V17971 n0_4929_6498 n2_4929_6498 0.0
V17972 n0_4929_6535 n2_4929_6535 0.0
V17973 n0_4929_6681 n2_4929_6681 0.0
V17974 n0_4929_6714 n2_4929_6714 0.0
V17975 n0_4929_6897 n2_4929_6897 0.0
V17976 n0_4929_6930 n2_4929_6930 0.0
V17977 n0_4929_7113 n2_4929_7113 0.0
V17978 n0_4929_7329 n2_4929_7329 0.0
V17979 n0_4929_7362 n2_4929_7362 0.0
V17980 n0_4929_7545 n2_4929_7545 0.0
V17981 n0_4929_7578 n2_4929_7578 0.0
V17982 n0_4929_7761 n2_4929_7761 0.0
V17983 n0_4929_7794 n2_4929_7794 0.0
V17984 n0_4929_7808 n2_4929_7808 0.0
V17985 n0_4929_7977 n2_4929_7977 0.0
V17986 n0_4929_8010 n2_4929_8010 0.0
V17987 n0_4929_8193 n2_4929_8193 0.0
V17988 n0_4929_8226 n2_4929_8226 0.0
V17989 n0_4929_8409 n2_4929_8409 0.0
V17990 n0_4929_8442 n2_4929_8442 0.0
V17991 n0_4929_8625 n2_4929_8625 0.0
V17992 n0_4929_8658 n2_4929_8658 0.0
V17993 n0_4929_8841 n2_4929_8841 0.0
V17994 n0_4929_8874 n2_4929_8874 0.0
V17995 n0_4929_8888 n2_4929_8888 0.0
V17996 n0_4929_8911 n2_4929_8911 0.0
V17997 n0_4929_9057 n2_4929_9057 0.0
V17998 n0_4929_9090 n2_4929_9090 0.0
V17999 n0_4929_9273 n2_4929_9273 0.0
V18000 n0_4929_9306 n2_4929_9306 0.0
V18001 n0_4929_9705 n2_4929_9705 0.0
V18002 n0_4929_9738 n2_4929_9738 0.0
V18003 n0_4929_9921 n2_4929_9921 0.0
V18004 n0_4929_9954 n2_4929_9954 0.0
V18005 n0_4929_9968 n2_4929_9968 0.0
V18006 n0_4929_10137 n2_4929_10137 0.0
V18007 n0_4929_10170 n2_4929_10170 0.0
V18008 n0_4929_10353 n2_4929_10353 0.0
V18009 n0_4929_10386 n2_4929_10386 0.0
V18010 n0_4929_10569 n2_4929_10569 0.0
V18011 n0_4929_10602 n2_4929_10602 0.0
V18012 n0_4929_10785 n2_4929_10785 0.0
V18013 n0_4929_10818 n2_4929_10818 0.0
V18014 n0_4929_11001 n2_4929_11001 0.0
V18015 n0_4929_11034 n2_4929_11034 0.0
V18016 n0_4929_11048 n2_4929_11048 0.0
V18017 n0_4929_11071 n2_4929_11071 0.0
V18018 n0_4929_11217 n2_4929_11217 0.0
V18019 n0_4929_11250 n2_4929_11250 0.0
V18020 n0_4929_11433 n2_4929_11433 0.0
V18021 n0_4929_11466 n2_4929_11466 0.0
V18022 n0_4929_11865 n2_4929_11865 0.0
V18023 n0_4929_11898 n2_4929_11898 0.0
V18024 n0_4929_12081 n2_4929_12081 0.0
V18025 n0_4929_12114 n2_4929_12114 0.0
V18026 n0_4929_12128 n2_4929_12128 0.0
V18027 n0_4929_12297 n2_4929_12297 0.0
V18028 n0_4929_12330 n2_4929_12330 0.0
V18029 n0_4929_12513 n2_4929_12513 0.0
V18030 n0_4929_12546 n2_4929_12546 0.0
V18031 n0_4929_12729 n2_4929_12729 0.0
V18032 n0_4929_12762 n2_4929_12762 0.0
V18033 n0_4929_12945 n2_4929_12945 0.0
V18034 n0_4929_12978 n2_4929_12978 0.0
V18035 n0_4929_13161 n2_4929_13161 0.0
V18036 n0_4929_13194 n2_4929_13194 0.0
V18037 n0_4929_13377 n2_4929_13377 0.0
V18038 n0_4929_13410 n2_4929_13410 0.0
V18039 n0_4929_13424 n2_4929_13424 0.0
V18040 n0_4929_13593 n2_4929_13593 0.0
V18041 n0_4929_13626 n2_4929_13626 0.0
V18042 n0_4929_13809 n2_4929_13809 0.0
V18043 n0_4929_13842 n2_4929_13842 0.0
V18044 n0_4929_14100 n2_4929_14100 0.0
V18045 n0_4929_14241 n2_4929_14241 0.0
V18046 n0_4929_14274 n2_4929_14274 0.0
V18047 n0_4929_14457 n2_4929_14457 0.0
V18048 n0_4929_14490 n2_4929_14490 0.0
V18049 n0_4929_14536 n2_4929_14536 0.0
V18050 n0_4929_14673 n2_4929_14673 0.0
V18051 n0_4929_14706 n2_4929_14706 0.0
V18052 n0_4929_14889 n2_4929_14889 0.0
V18053 n0_4929_14922 n2_4929_14922 0.0
V18054 n0_4929_15105 n2_4929_15105 0.0
V18055 n0_4929_15138 n2_4929_15138 0.0
V18056 n0_4929_15321 n2_4929_15321 0.0
V18057 n0_4929_15354 n2_4929_15354 0.0
V18058 n0_4929_15368 n2_4929_15368 0.0
V18059 n0_4929_15537 n2_4929_15537 0.0
V18060 n0_4929_15570 n2_4929_15570 0.0
V18061 n0_4929_15584 n2_4929_15584 0.0
V18062 n0_4929_15753 n2_4929_15753 0.0
V18063 n0_4929_15786 n2_4929_15786 0.0
V18064 n0_4929_15969 n2_4929_15969 0.0
V18065 n0_4929_16002 n2_4929_16002 0.0
V18066 n0_4929_16016 n2_4929_16016 0.0
V18067 n0_5866_201 n2_5866_201 0.0
V18068 n0_5866_234 n2_5866_234 0.0
V18069 n0_5866_356 n2_5866_356 0.0
V18070 n0_5866_417 n2_5866_417 0.0
V18071 n0_5866_450 n2_5866_450 0.0
V18072 n0_5866_633 n2_5866_633 0.0
V18073 n0_5866_666 n2_5866_666 0.0
V18074 n0_5866_788 n2_5866_788 0.0
V18075 n0_5866_849 n2_5866_849 0.0
V18076 n0_5866_882 n2_5866_882 0.0
V18077 n0_5866_1065 n2_5866_1065 0.0
V18078 n0_5866_1098 n2_5866_1098 0.0
V18079 n0_5866_1281 n2_5866_1281 0.0
V18080 n0_5866_1314 n2_5866_1314 0.0
V18081 n0_5866_1497 n2_5866_1497 0.0
V18082 n0_5866_1530 n2_5866_1530 0.0
V18083 n0_5866_1713 n2_5866_1713 0.0
V18084 n0_5866_1746 n2_5866_1746 0.0
V18085 n0_5866_1760 n2_5866_1760 0.0
V18086 n0_5866_1929 n2_5866_1929 0.0
V18087 n0_5866_1962 n2_5866_1962 0.0
V18088 n0_5866_2145 n2_5866_2145 0.0
V18089 n0_5866_2178 n2_5866_2178 0.0
V18090 n0_5866_2361 n2_5866_2361 0.0
V18091 n0_5866_2394 n2_5866_2394 0.0
V18092 n0_5866_2408 n2_5866_2408 0.0
V18093 n0_5866_2577 n2_5866_2577 0.0
V18094 n0_5866_2610 n2_5866_2610 0.0
V18095 n0_5866_2793 n2_5866_2793 0.0
V18096 n0_5866_2826 n2_5866_2826 0.0
V18097 n0_5866_2840 n2_5866_2840 0.0
V18098 n0_5866_3009 n2_5866_3009 0.0
V18099 n0_5866_3042 n2_5866_3042 0.0
V18100 n0_5866_3056 n2_5866_3056 0.0
V18101 n0_5866_3225 n2_5866_3225 0.0
V18102 n0_5866_3258 n2_5866_3258 0.0
V18103 n0_5866_3441 n2_5866_3441 0.0
V18104 n0_5866_3474 n2_5866_3474 0.0
V18105 n0_5866_3488 n2_5866_3488 0.0
V18106 n0_5866_3657 n2_5866_3657 0.0
V18107 n0_5866_3690 n2_5866_3690 0.0
V18108 n0_5866_3873 n2_5866_3873 0.0
V18109 n0_5866_3906 n2_5866_3906 0.0
V18110 n0_5866_4089 n2_5866_4089 0.0
V18111 n0_5866_4122 n2_5866_4122 0.0
V18112 n0_5866_4136 n2_5866_4136 0.0
V18113 n0_5866_4305 n2_5866_4305 0.0
V18114 n0_5866_4338 n2_5866_4338 0.0
V18115 n0_5866_4352 n2_5866_4352 0.0
V18116 n0_5866_4375 n2_5866_4375 0.0
V18117 n0_5866_4521 n2_5866_4521 0.0
V18118 n0_5866_4554 n2_5866_4554 0.0
V18119 n0_5866_4568 n2_5866_4568 0.0
V18120 n0_5866_4737 n2_5866_4737 0.0
V18121 n0_5866_4770 n2_5866_4770 0.0
V18122 n0_5866_4953 n2_5866_4953 0.0
V18123 n0_5866_5169 n2_5866_5169 0.0
V18124 n0_5866_5202 n2_5866_5202 0.0
V18125 n0_5866_5216 n2_5866_5216 0.0
V18126 n0_5866_5385 n2_5866_5385 0.0
V18127 n0_5866_5418 n2_5866_5418 0.0
V18128 n0_5866_5432 n2_5866_5432 0.0
V18129 n0_5866_5455 n2_5866_5455 0.0
V18130 n0_5866_5601 n2_5866_5601 0.0
V18131 n0_5866_5634 n2_5866_5634 0.0
V18132 n0_5866_5817 n2_5866_5817 0.0
V18133 n0_5866_5850 n2_5866_5850 0.0
V18134 n0_5866_6033 n2_5866_6033 0.0
V18135 n0_5866_6066 n2_5866_6066 0.0
V18136 n0_5866_6249 n2_5866_6249 0.0
V18137 n0_5866_6282 n2_5866_6282 0.0
V18138 n0_5866_6465 n2_5866_6465 0.0
V18139 n0_5866_6498 n2_5866_6498 0.0
V18140 n0_5866_6535 n2_5866_6535 0.0
V18141 n0_5866_6681 n2_5866_6681 0.0
V18142 n0_5866_6714 n2_5866_6714 0.0
V18143 n0_5866_6897 n2_5866_6897 0.0
V18144 n0_5866_6930 n2_5866_6930 0.0
V18145 n0_5866_7113 n2_5866_7113 0.0
V18146 n0_5866_7146 n2_5866_7146 0.0
V18147 n0_5866_7329 n2_5866_7329 0.0
V18148 n0_5866_7362 n2_5866_7362 0.0
V18149 n0_5866_7545 n2_5866_7545 0.0
V18150 n0_5866_7578 n2_5866_7578 0.0
V18151 n0_5866_7761 n2_5866_7761 0.0
V18152 n0_5866_7794 n2_5866_7794 0.0
V18153 n0_5866_7808 n2_5866_7808 0.0
V18154 n0_5866_7977 n2_5866_7977 0.0
V18155 n0_5866_8010 n2_5866_8010 0.0
V18156 n0_5866_8193 n2_5866_8193 0.0
V18157 n0_5866_8226 n2_5866_8226 0.0
V18158 n0_5866_8409 n2_5866_8409 0.0
V18159 n0_5866_8442 n2_5866_8442 0.0
V18160 n0_5866_8625 n2_5866_8625 0.0
V18161 n0_5866_8658 n2_5866_8658 0.0
V18162 n0_5866_8841 n2_5866_8841 0.0
V18163 n0_5866_8874 n2_5866_8874 0.0
V18164 n0_5866_8888 n2_5866_8888 0.0
V18165 n0_5866_8911 n2_5866_8911 0.0
V18166 n0_5866_9057 n2_5866_9057 0.0
V18167 n0_5866_9090 n2_5866_9090 0.0
V18168 n0_5866_9273 n2_5866_9273 0.0
V18169 n0_5866_9306 n2_5866_9306 0.0
V18170 n0_5866_9489 n2_5866_9489 0.0
V18171 n0_5866_9522 n2_5866_9522 0.0
V18172 n0_5866_9705 n2_5866_9705 0.0
V18173 n0_5866_9738 n2_5866_9738 0.0
V18174 n0_5866_9921 n2_5866_9921 0.0
V18175 n0_5866_9954 n2_5866_9954 0.0
V18176 n0_5866_9968 n2_5866_9968 0.0
V18177 n0_5866_10137 n2_5866_10137 0.0
V18178 n0_5866_10170 n2_5866_10170 0.0
V18179 n0_5866_10353 n2_5866_10353 0.0
V18180 n0_5866_10386 n2_5866_10386 0.0
V18181 n0_5866_10569 n2_5866_10569 0.0
V18182 n0_5866_10785 n2_5866_10785 0.0
V18183 n0_5866_10818 n2_5866_10818 0.0
V18184 n0_5866_11001 n2_5866_11001 0.0
V18185 n0_5866_11034 n2_5866_11034 0.0
V18186 n0_5866_11048 n2_5866_11048 0.0
V18187 n0_5866_11071 n2_5866_11071 0.0
V18188 n0_5866_11217 n2_5866_11217 0.0
V18189 n0_5866_11250 n2_5866_11250 0.0
V18190 n0_5866_11433 n2_5866_11433 0.0
V18191 n0_5866_11466 n2_5866_11466 0.0
V18192 n0_5866_11649 n2_5866_11649 0.0
V18193 n0_5866_11682 n2_5866_11682 0.0
V18194 n0_5866_11865 n2_5866_11865 0.0
V18195 n0_5866_11898 n2_5866_11898 0.0
V18196 n0_5866_12081 n2_5866_12081 0.0
V18197 n0_5866_12114 n2_5866_12114 0.0
V18198 n0_5866_12128 n2_5866_12128 0.0
V18199 n0_5866_12297 n2_5866_12297 0.0
V18200 n0_5866_12330 n2_5866_12330 0.0
V18201 n0_5866_12513 n2_5866_12513 0.0
V18202 n0_5866_12546 n2_5866_12546 0.0
V18203 n0_5866_12729 n2_5866_12729 0.0
V18204 n0_5866_12762 n2_5866_12762 0.0
V18205 n0_5866_12945 n2_5866_12945 0.0
V18206 n0_5866_12978 n2_5866_12978 0.0
V18207 n0_5866_13161 n2_5866_13161 0.0
V18208 n0_5866_13194 n2_5866_13194 0.0
V18209 n0_5866_13377 n2_5866_13377 0.0
V18210 n0_5866_13410 n2_5866_13410 0.0
V18211 n0_5866_13424 n2_5866_13424 0.0
V18212 n0_5866_13593 n2_5866_13593 0.0
V18213 n0_5866_13626 n2_5866_13626 0.0
V18214 n0_5866_13809 n2_5866_13809 0.0
V18215 n0_5866_13842 n2_5866_13842 0.0
V18216 n0_5866_13879 n2_5866_13879 0.0
V18217 n0_5866_14025 n2_5866_14025 0.0
V18218 n0_5866_14058 n2_5866_14058 0.0
V18219 n0_5866_14241 n2_5866_14241 0.0
V18220 n0_5866_14274 n2_5866_14274 0.0
V18221 n0_5866_14457 n2_5866_14457 0.0
V18222 n0_5866_14490 n2_5866_14490 0.0
V18223 n0_5866_14536 n2_5866_14536 0.0
V18224 n0_5866_14673 n2_5866_14673 0.0
V18225 n0_5866_14706 n2_5866_14706 0.0
V18226 n0_5866_14889 n2_5866_14889 0.0
V18227 n0_5866_14922 n2_5866_14922 0.0
V18228 n0_5866_15138 n2_5866_15138 0.0
V18229 n0_5866_15321 n2_5866_15321 0.0
V18230 n0_5866_15354 n2_5866_15354 0.0
V18231 n0_5866_15537 n2_5866_15537 0.0
V18232 n0_5866_15570 n2_5866_15570 0.0
V18233 n0_5866_15584 n2_5866_15584 0.0
V18234 n0_5866_15753 n2_5866_15753 0.0
V18235 n0_5866_15786 n2_5866_15786 0.0
V18236 n0_5866_15800 n2_5866_15800 0.0
V18237 n0_5866_15969 n2_5866_15969 0.0
V18238 n0_5866_16002 n2_5866_16002 0.0
V18239 n0_5866_16016 n2_5866_16016 0.0
V18240 n0_5866_16185 n2_5866_16185 0.0
V18241 n0_5866_16401 n2_5866_16401 0.0
V18242 n0_5866_16434 n2_5866_16434 0.0
V18243 n0_5866_16617 n2_5866_16617 0.0
V18244 n0_5866_16650 n2_5866_16650 0.0
V18245 n0_5866_16833 n2_5866_16833 0.0
V18246 n0_5866_16866 n2_5866_16866 0.0
V18247 n0_5866_17049 n2_5866_17049 0.0
V18248 n0_5866_17082 n2_5866_17082 0.0
V18249 n0_5866_17096 n2_5866_17096 0.0
V18250 n0_5866_17119 n2_5866_17119 0.0
V18251 n0_5866_17265 n2_5866_17265 0.0
V18252 n0_5866_17298 n2_5866_17298 0.0
V18253 n0_5866_17312 n2_5866_17312 0.0
V18254 n0_5866_17481 n2_5866_17481 0.0
V18255 n0_5866_17514 n2_5866_17514 0.0
V18256 n0_5866_17528 n2_5866_17528 0.0
V18257 n0_5866_17697 n2_5866_17697 0.0
V18258 n0_5866_17730 n2_5866_17730 0.0
V18259 n0_5866_17913 n2_5866_17913 0.0
V18260 n0_5866_17946 n2_5866_17946 0.0
V18261 n0_5866_18129 n2_5866_18129 0.0
V18262 n0_5866_18162 n2_5866_18162 0.0
V18263 n0_5866_18345 n2_5866_18345 0.0
V18264 n0_5866_18378 n2_5866_18378 0.0
V18265 n0_5866_18392 n2_5866_18392 0.0
V18266 n0_5866_18561 n2_5866_18561 0.0
V18267 n0_5866_18594 n2_5866_18594 0.0
V18268 n0_5866_18608 n2_5866_18608 0.0
V18269 n0_5866_18777 n2_5866_18777 0.0
V18270 n0_5866_18810 n2_5866_18810 0.0
V18271 n0_5866_18824 n2_5866_18824 0.0
V18272 n0_5866_18993 n2_5866_18993 0.0
V18273 n0_5866_19026 n2_5866_19026 0.0
V18274 n0_5866_19040 n2_5866_19040 0.0
V18275 n0_5866_19209 n2_5866_19209 0.0
V18276 n0_5866_19242 n2_5866_19242 0.0
V18277 n0_5866_19425 n2_5866_19425 0.0
V18278 n0_5866_19458 n2_5866_19458 0.0
V18279 n0_5866_19472 n2_5866_19472 0.0
V18280 n0_5866_19641 n2_5866_19641 0.0
V18281 n0_5866_19674 n2_5866_19674 0.0
V18282 n0_5866_19857 n2_5866_19857 0.0
V18283 n0_5866_19890 n2_5866_19890 0.0
V18284 n0_5866_20073 n2_5866_20073 0.0
V18285 n0_5866_20106 n2_5866_20106 0.0
V18286 n0_5866_20289 n2_5866_20289 0.0
V18287 n0_5866_20322 n2_5866_20322 0.0
V18288 n0_5866_20505 n2_5866_20505 0.0
V18289 n0_5866_20538 n2_5866_20538 0.0
V18290 n0_5866_20754 n2_5866_20754 0.0
V18291 n0_5866_20937 n2_5866_20937 0.0
V18292 n0_5866_20970 n2_5866_20970 0.0
V18293 n0_5958_201 n2_5958_201 0.0
V18294 n0_5958_234 n2_5958_234 0.0
V18295 n0_5958_356 n2_5958_356 0.0
V18296 n0_5958_417 n2_5958_417 0.0
V18297 n0_5958_450 n2_5958_450 0.0
V18298 n0_5958_633 n2_5958_633 0.0
V18299 n0_5958_666 n2_5958_666 0.0
V18300 n0_5958_788 n2_5958_788 0.0
V18301 n0_5958_849 n2_5958_849 0.0
V18302 n0_5958_882 n2_5958_882 0.0
V18303 n0_5958_1065 n2_5958_1065 0.0
V18304 n0_5958_1098 n2_5958_1098 0.0
V18305 n0_5958_1281 n2_5958_1281 0.0
V18306 n0_5958_1314 n2_5958_1314 0.0
V18307 n0_5958_1497 n2_5958_1497 0.0
V18308 n0_5958_1530 n2_5958_1530 0.0
V18309 n0_5958_1713 n2_5958_1713 0.0
V18310 n0_5958_1746 n2_5958_1746 0.0
V18311 n0_5958_1760 n2_5958_1760 0.0
V18312 n0_5958_1929 n2_5958_1929 0.0
V18313 n0_5958_1962 n2_5958_1962 0.0
V18314 n0_5958_2145 n2_5958_2145 0.0
V18315 n0_5958_2178 n2_5958_2178 0.0
V18316 n0_5958_2361 n2_5958_2361 0.0
V18317 n0_5958_2394 n2_5958_2394 0.0
V18318 n0_5958_2408 n2_5958_2408 0.0
V18319 n0_5958_2577 n2_5958_2577 0.0
V18320 n0_5958_2610 n2_5958_2610 0.0
V18321 n0_5958_2793 n2_5958_2793 0.0
V18322 n0_5958_2826 n2_5958_2826 0.0
V18323 n0_5958_2840 n2_5958_2840 0.0
V18324 n0_5958_3009 n2_5958_3009 0.0
V18325 n0_5958_3042 n2_5958_3042 0.0
V18326 n0_5958_3056 n2_5958_3056 0.0
V18327 n0_5958_3225 n2_5958_3225 0.0
V18328 n0_5958_3258 n2_5958_3258 0.0
V18329 n0_5958_3441 n2_5958_3441 0.0
V18330 n0_5958_3474 n2_5958_3474 0.0
V18331 n0_5958_3488 n2_5958_3488 0.0
V18332 n0_5958_3657 n2_5958_3657 0.0
V18333 n0_5958_3690 n2_5958_3690 0.0
V18334 n0_5958_3873 n2_5958_3873 0.0
V18335 n0_5958_3906 n2_5958_3906 0.0
V18336 n0_5958_4089 n2_5958_4089 0.0
V18337 n0_5958_4122 n2_5958_4122 0.0
V18338 n0_5958_4136 n2_5958_4136 0.0
V18339 n0_5958_4305 n2_5958_4305 0.0
V18340 n0_5958_4338 n2_5958_4338 0.0
V18341 n0_5958_4352 n2_5958_4352 0.0
V18342 n0_5958_4375 n2_5958_4375 0.0
V18343 n0_5958_4521 n2_5958_4521 0.0
V18344 n0_5958_4554 n2_5958_4554 0.0
V18345 n0_5958_4568 n2_5958_4568 0.0
V18346 n0_5958_4737 n2_5958_4737 0.0
V18347 n0_5958_4770 n2_5958_4770 0.0
V18348 n0_5958_4953 n2_5958_4953 0.0
V18349 n0_5958_4986 n2_5958_4986 0.0
V18350 n0_5958_5169 n2_5958_5169 0.0
V18351 n0_5958_5202 n2_5958_5202 0.0
V18352 n0_5958_5216 n2_5958_5216 0.0
V18353 n0_5958_5385 n2_5958_5385 0.0
V18354 n0_5958_5418 n2_5958_5418 0.0
V18355 n0_5958_5432 n2_5958_5432 0.0
V18356 n0_5958_5455 n2_5958_5455 0.0
V18357 n0_5958_5601 n2_5958_5601 0.0
V18358 n0_5958_5634 n2_5958_5634 0.0
V18359 n0_5958_5817 n2_5958_5817 0.0
V18360 n0_5958_5850 n2_5958_5850 0.0
V18361 n0_5958_6033 n2_5958_6033 0.0
V18362 n0_5958_6066 n2_5958_6066 0.0
V18363 n0_5958_15105 n2_5958_15105 0.0
V18364 n0_5958_15138 n2_5958_15138 0.0
V18365 n0_5958_15321 n2_5958_15321 0.0
V18366 n0_5958_15354 n2_5958_15354 0.0
V18367 n0_5958_15537 n2_5958_15537 0.0
V18368 n0_5958_15570 n2_5958_15570 0.0
V18369 n0_5958_15584 n2_5958_15584 0.0
V18370 n0_5958_15753 n2_5958_15753 0.0
V18371 n0_5958_15786 n2_5958_15786 0.0
V18372 n0_5958_15800 n2_5958_15800 0.0
V18373 n0_5958_15969 n2_5958_15969 0.0
V18374 n0_5958_16002 n2_5958_16002 0.0
V18375 n0_5958_16016 n2_5958_16016 0.0
V18376 n0_5958_16185 n2_5958_16185 0.0
V18377 n0_5958_16218 n2_5958_16218 0.0
V18378 n0_5958_16401 n2_5958_16401 0.0
V18379 n0_5958_16434 n2_5958_16434 0.0
V18380 n0_5958_16617 n2_5958_16617 0.0
V18381 n0_5958_16650 n2_5958_16650 0.0
V18382 n0_5958_16833 n2_5958_16833 0.0
V18383 n0_5958_16866 n2_5958_16866 0.0
V18384 n0_5958_17049 n2_5958_17049 0.0
V18385 n0_5958_17082 n2_5958_17082 0.0
V18386 n0_5958_17096 n2_5958_17096 0.0
V18387 n0_5958_17119 n2_5958_17119 0.0
V18388 n0_5958_17265 n2_5958_17265 0.0
V18389 n0_5958_17298 n2_5958_17298 0.0
V18390 n0_5958_17312 n2_5958_17312 0.0
V18391 n0_5958_17335 n2_5958_17335 0.0
V18392 n0_5958_17481 n2_5958_17481 0.0
V18393 n0_5958_17514 n2_5958_17514 0.0
V18394 n0_5958_17528 n2_5958_17528 0.0
V18395 n0_5958_17697 n2_5958_17697 0.0
V18396 n0_5958_17730 n2_5958_17730 0.0
V18397 n0_5958_17913 n2_5958_17913 0.0
V18398 n0_5958_17946 n2_5958_17946 0.0
V18399 n0_5958_18129 n2_5958_18129 0.0
V18400 n0_5958_18162 n2_5958_18162 0.0
V18401 n0_5958_18345 n2_5958_18345 0.0
V18402 n0_5958_18378 n2_5958_18378 0.0
V18403 n0_5958_18392 n2_5958_18392 0.0
V18404 n0_5958_18561 n2_5958_18561 0.0
V18405 n0_5958_18594 n2_5958_18594 0.0
V18406 n0_5958_18608 n2_5958_18608 0.0
V18407 n0_5958_18777 n2_5958_18777 0.0
V18408 n0_5958_18810 n2_5958_18810 0.0
V18409 n0_5958_18824 n2_5958_18824 0.0
V18410 n0_5958_18993 n2_5958_18993 0.0
V18411 n0_5958_19026 n2_5958_19026 0.0
V18412 n0_5958_19040 n2_5958_19040 0.0
V18413 n0_5958_19209 n2_5958_19209 0.0
V18414 n0_5958_19242 n2_5958_19242 0.0
V18415 n0_5958_19425 n2_5958_19425 0.0
V18416 n0_5958_19458 n2_5958_19458 0.0
V18417 n0_5958_19472 n2_5958_19472 0.0
V18418 n0_5958_19641 n2_5958_19641 0.0
V18419 n0_5958_19674 n2_5958_19674 0.0
V18420 n0_5958_19857 n2_5958_19857 0.0
V18421 n0_5958_19890 n2_5958_19890 0.0
V18422 n0_5958_20073 n2_5958_20073 0.0
V18423 n0_5958_20106 n2_5958_20106 0.0
V18424 n0_5958_20289 n2_5958_20289 0.0
V18425 n0_5958_20322 n2_5958_20322 0.0
V18426 n0_5958_20505 n2_5958_20505 0.0
V18427 n0_5958_20538 n2_5958_20538 0.0
V18428 n0_5958_20721 n2_5958_20721 0.0
V18429 n0_5958_20754 n2_5958_20754 0.0
V18430 n0_5958_20937 n2_5958_20937 0.0
V18431 n0_5958_20970 n2_5958_20970 0.0
V18432 n0_6005_417 n2_6005_417 0.0
V18433 n0_6005_450 n2_6005_450 0.0
V18434 n0_6005_1530 n2_6005_1530 0.0
V18435 n0_6005_2793 n2_6005_2793 0.0
V18436 n0_6005_3873 n2_6005_3873 0.0
V18437 n0_6005_3906 n2_6005_3906 0.0
V18438 n0_6005_4953 n2_6005_4953 0.0
V18439 n0_6005_4986 n2_6005_4986 0.0
V18440 n0_6005_6033 n2_6005_6033 0.0
V18441 n0_6005_6066 n2_6005_6066 0.0
V18442 n0_6005_8409 n2_6005_8409 0.0
V18443 n0_6005_10569 n2_6005_10569 0.0
V18444 n0_6005_10602 n2_6005_10602 0.0
V18445 n0_6005_15105 n2_6005_15105 0.0
V18446 n0_6005_15138 n2_6005_15138 0.0
V18447 n0_6005_16185 n2_6005_16185 0.0
V18448 n0_6005_16218 n2_6005_16218 0.0
V18449 n0_6005_17298 n2_6005_17298 0.0
V18450 n0_6005_17312 n2_6005_17312 0.0
V18451 n0_6005_17335 n2_6005_17335 0.0
V18452 n0_6005_18392 n2_6005_18392 0.0
V18453 n0_6005_19641 n2_6005_19641 0.0
V18454 n0_6005_19674 n2_6005_19674 0.0
V18455 n0_6005_20721 n2_6005_20721 0.0
V18456 n0_6005_20754 n2_6005_20754 0.0
V18457 n0_6054_201 n2_6054_201 0.0
V18458 n0_6054_234 n2_6054_234 0.0
V18459 n0_6054_356 n2_6054_356 0.0
V18460 n0_6054_417 n2_6054_417 0.0
V18461 n0_6054_450 n2_6054_450 0.0
V18462 n0_6054_633 n2_6054_633 0.0
V18463 n0_6054_666 n2_6054_666 0.0
V18464 n0_6054_788 n2_6054_788 0.0
V18465 n0_6054_849 n2_6054_849 0.0
V18466 n0_6054_882 n2_6054_882 0.0
V18467 n0_6054_1065 n2_6054_1065 0.0
V18468 n0_6054_1098 n2_6054_1098 0.0
V18469 n0_6054_1281 n2_6054_1281 0.0
V18470 n0_6054_1314 n2_6054_1314 0.0
V18471 n0_6054_1497 n2_6054_1497 0.0
V18472 n0_6054_1530 n2_6054_1530 0.0
V18473 n0_6054_1713 n2_6054_1713 0.0
V18474 n0_6054_1746 n2_6054_1746 0.0
V18475 n0_6054_1760 n2_6054_1760 0.0
V18476 n0_6054_1929 n2_6054_1929 0.0
V18477 n0_6054_1962 n2_6054_1962 0.0
V18478 n0_6054_2145 n2_6054_2145 0.0
V18479 n0_6054_2178 n2_6054_2178 0.0
V18480 n0_6054_2361 n2_6054_2361 0.0
V18481 n0_6054_2394 n2_6054_2394 0.0
V18482 n0_6054_2408 n2_6054_2408 0.0
V18483 n0_6054_2577 n2_6054_2577 0.0
V18484 n0_6054_2610 n2_6054_2610 0.0
V18485 n0_6054_2793 n2_6054_2793 0.0
V18486 n0_6054_2826 n2_6054_2826 0.0
V18487 n0_6054_2840 n2_6054_2840 0.0
V18488 n0_6054_3009 n2_6054_3009 0.0
V18489 n0_6054_3042 n2_6054_3042 0.0
V18490 n0_6054_3056 n2_6054_3056 0.0
V18491 n0_6054_3225 n2_6054_3225 0.0
V18492 n0_6054_3258 n2_6054_3258 0.0
V18493 n0_6054_3441 n2_6054_3441 0.0
V18494 n0_6054_3474 n2_6054_3474 0.0
V18495 n0_6054_3488 n2_6054_3488 0.0
V18496 n0_6054_3657 n2_6054_3657 0.0
V18497 n0_6054_3690 n2_6054_3690 0.0
V18498 n0_6054_3873 n2_6054_3873 0.0
V18499 n0_6054_3906 n2_6054_3906 0.0
V18500 n0_6054_4089 n2_6054_4089 0.0
V18501 n0_6054_4122 n2_6054_4122 0.0
V18502 n0_6054_4136 n2_6054_4136 0.0
V18503 n0_6054_4305 n2_6054_4305 0.0
V18504 n0_6054_4338 n2_6054_4338 0.0
V18505 n0_6054_4352 n2_6054_4352 0.0
V18506 n0_6054_4375 n2_6054_4375 0.0
V18507 n0_6054_4521 n2_6054_4521 0.0
V18508 n0_6054_4554 n2_6054_4554 0.0
V18509 n0_6054_4568 n2_6054_4568 0.0
V18510 n0_6054_4737 n2_6054_4737 0.0
V18511 n0_6054_4770 n2_6054_4770 0.0
V18512 n0_6054_4953 n2_6054_4953 0.0
V18513 n0_6054_4986 n2_6054_4986 0.0
V18514 n0_6054_5169 n2_6054_5169 0.0
V18515 n0_6054_5202 n2_6054_5202 0.0
V18516 n0_6054_5216 n2_6054_5216 0.0
V18517 n0_6054_5385 n2_6054_5385 0.0
V18518 n0_6054_5418 n2_6054_5418 0.0
V18519 n0_6054_5432 n2_6054_5432 0.0
V18520 n0_6054_5455 n2_6054_5455 0.0
V18521 n0_6054_5601 n2_6054_5601 0.0
V18522 n0_6054_5634 n2_6054_5634 0.0
V18523 n0_6054_5817 n2_6054_5817 0.0
V18524 n0_6054_5850 n2_6054_5850 0.0
V18525 n0_6054_6033 n2_6054_6033 0.0
V18526 n0_6054_6066 n2_6054_6066 0.0
V18527 n0_6054_6249 n2_6054_6249 0.0
V18528 n0_6054_6282 n2_6054_6282 0.0
V18529 n0_6054_6465 n2_6054_6465 0.0
V18530 n0_6054_6498 n2_6054_6498 0.0
V18531 n0_6054_6535 n2_6054_6535 0.0
V18532 n0_6054_6681 n2_6054_6681 0.0
V18533 n0_6054_6714 n2_6054_6714 0.0
V18534 n0_6054_6897 n2_6054_6897 0.0
V18535 n0_6054_6930 n2_6054_6930 0.0
V18536 n0_6054_7113 n2_6054_7113 0.0
V18537 n0_6054_7329 n2_6054_7329 0.0
V18538 n0_6054_7362 n2_6054_7362 0.0
V18539 n0_6054_7545 n2_6054_7545 0.0
V18540 n0_6054_7578 n2_6054_7578 0.0
V18541 n0_6054_7761 n2_6054_7761 0.0
V18542 n0_6054_7794 n2_6054_7794 0.0
V18543 n0_6054_7808 n2_6054_7808 0.0
V18544 n0_6054_7977 n2_6054_7977 0.0
V18545 n0_6054_8010 n2_6054_8010 0.0
V18546 n0_6054_8193 n2_6054_8193 0.0
V18547 n0_6054_8226 n2_6054_8226 0.0
V18548 n0_6054_8409 n2_6054_8409 0.0
V18549 n0_6054_8442 n2_6054_8442 0.0
V18550 n0_6054_8625 n2_6054_8625 0.0
V18551 n0_6054_8658 n2_6054_8658 0.0
V18552 n0_6054_8841 n2_6054_8841 0.0
V18553 n0_6054_8874 n2_6054_8874 0.0
V18554 n0_6054_8888 n2_6054_8888 0.0
V18555 n0_6054_8911 n2_6054_8911 0.0
V18556 n0_6054_9057 n2_6054_9057 0.0
V18557 n0_6054_9090 n2_6054_9090 0.0
V18558 n0_6054_9273 n2_6054_9273 0.0
V18559 n0_6054_9306 n2_6054_9306 0.0
V18560 n0_6054_9705 n2_6054_9705 0.0
V18561 n0_6054_9738 n2_6054_9738 0.0
V18562 n0_6054_9921 n2_6054_9921 0.0
V18563 n0_6054_9954 n2_6054_9954 0.0
V18564 n0_6054_9968 n2_6054_9968 0.0
V18565 n0_6054_10137 n2_6054_10137 0.0
V18566 n0_6054_10170 n2_6054_10170 0.0
V18567 n0_6054_10353 n2_6054_10353 0.0
V18568 n0_6054_10386 n2_6054_10386 0.0
V18569 n0_6054_10569 n2_6054_10569 0.0
V18570 n0_6054_10602 n2_6054_10602 0.0
V18571 n0_6054_10785 n2_6054_10785 0.0
V18572 n0_6054_10818 n2_6054_10818 0.0
V18573 n0_6054_11001 n2_6054_11001 0.0
V18574 n0_6054_11034 n2_6054_11034 0.0
V18575 n0_6054_11048 n2_6054_11048 0.0
V18576 n0_6054_11071 n2_6054_11071 0.0
V18577 n0_6054_11217 n2_6054_11217 0.0
V18578 n0_6054_11250 n2_6054_11250 0.0
V18579 n0_6054_11433 n2_6054_11433 0.0
V18580 n0_6054_11466 n2_6054_11466 0.0
V18581 n0_6054_11865 n2_6054_11865 0.0
V18582 n0_6054_11898 n2_6054_11898 0.0
V18583 n0_6054_12081 n2_6054_12081 0.0
V18584 n0_6054_12114 n2_6054_12114 0.0
V18585 n0_6054_12128 n2_6054_12128 0.0
V18586 n0_6054_12297 n2_6054_12297 0.0
V18587 n0_6054_12330 n2_6054_12330 0.0
V18588 n0_6054_12513 n2_6054_12513 0.0
V18589 n0_6054_12546 n2_6054_12546 0.0
V18590 n0_6054_12729 n2_6054_12729 0.0
V18591 n0_6054_12762 n2_6054_12762 0.0
V18592 n0_6054_12945 n2_6054_12945 0.0
V18593 n0_6054_12978 n2_6054_12978 0.0
V18594 n0_6054_13161 n2_6054_13161 0.0
V18595 n0_6054_13194 n2_6054_13194 0.0
V18596 n0_6054_13377 n2_6054_13377 0.0
V18597 n0_6054_13410 n2_6054_13410 0.0
V18598 n0_6054_13424 n2_6054_13424 0.0
V18599 n0_6054_13593 n2_6054_13593 0.0
V18600 n0_6054_13626 n2_6054_13626 0.0
V18601 n0_6054_13809 n2_6054_13809 0.0
V18602 n0_6054_13842 n2_6054_13842 0.0
V18603 n0_6054_14241 n2_6054_14241 0.0
V18604 n0_6054_14274 n2_6054_14274 0.0
V18605 n0_6054_14457 n2_6054_14457 0.0
V18606 n0_6054_14490 n2_6054_14490 0.0
V18607 n0_6054_14536 n2_6054_14536 0.0
V18608 n0_6054_14673 n2_6054_14673 0.0
V18609 n0_6054_14706 n2_6054_14706 0.0
V18610 n0_6054_14889 n2_6054_14889 0.0
V18611 n0_6054_14922 n2_6054_14922 0.0
V18612 n0_6054_15105 n2_6054_15105 0.0
V18613 n0_6054_15138 n2_6054_15138 0.0
V18614 n0_6054_15321 n2_6054_15321 0.0
V18615 n0_6054_15354 n2_6054_15354 0.0
V18616 n0_6054_15537 n2_6054_15537 0.0
V18617 n0_6054_15570 n2_6054_15570 0.0
V18618 n0_6054_15584 n2_6054_15584 0.0
V18619 n0_6054_15753 n2_6054_15753 0.0
V18620 n0_6054_15786 n2_6054_15786 0.0
V18621 n0_6054_15800 n2_6054_15800 0.0
V18622 n0_6054_15969 n2_6054_15969 0.0
V18623 n0_6054_16002 n2_6054_16002 0.0
V18624 n0_6054_16016 n2_6054_16016 0.0
V18625 n0_6054_16185 n2_6054_16185 0.0
V18626 n0_6054_16218 n2_6054_16218 0.0
V18627 n0_6054_16401 n2_6054_16401 0.0
V18628 n0_6054_16434 n2_6054_16434 0.0
V18629 n0_6054_16617 n2_6054_16617 0.0
V18630 n0_6054_16650 n2_6054_16650 0.0
V18631 n0_6054_16833 n2_6054_16833 0.0
V18632 n0_6054_16866 n2_6054_16866 0.0
V18633 n0_6054_17049 n2_6054_17049 0.0
V18634 n0_6054_17082 n2_6054_17082 0.0
V18635 n0_6054_17096 n2_6054_17096 0.0
V18636 n0_6054_17119 n2_6054_17119 0.0
V18637 n0_6054_17265 n2_6054_17265 0.0
V18638 n0_6054_17298 n2_6054_17298 0.0
V18639 n0_6054_17312 n2_6054_17312 0.0
V18640 n0_6054_17335 n2_6054_17335 0.0
V18641 n0_6054_17481 n2_6054_17481 0.0
V18642 n0_6054_17514 n2_6054_17514 0.0
V18643 n0_6054_17528 n2_6054_17528 0.0
V18644 n0_6054_17697 n2_6054_17697 0.0
V18645 n0_6054_17730 n2_6054_17730 0.0
V18646 n0_6054_17913 n2_6054_17913 0.0
V18647 n0_6054_17946 n2_6054_17946 0.0
V18648 n0_6054_18129 n2_6054_18129 0.0
V18649 n0_6054_18162 n2_6054_18162 0.0
V18650 n0_6054_18345 n2_6054_18345 0.0
V18651 n0_6054_18378 n2_6054_18378 0.0
V18652 n0_6054_18392 n2_6054_18392 0.0
V18653 n0_6054_18561 n2_6054_18561 0.0
V18654 n0_6054_18594 n2_6054_18594 0.0
V18655 n0_6054_18608 n2_6054_18608 0.0
V18656 n0_6054_18777 n2_6054_18777 0.0
V18657 n0_6054_18810 n2_6054_18810 0.0
V18658 n0_6054_18824 n2_6054_18824 0.0
V18659 n0_6054_18993 n2_6054_18993 0.0
V18660 n0_6054_19026 n2_6054_19026 0.0
V18661 n0_6054_19040 n2_6054_19040 0.0
V18662 n0_6054_19209 n2_6054_19209 0.0
V18663 n0_6054_19242 n2_6054_19242 0.0
V18664 n0_6054_19425 n2_6054_19425 0.0
V18665 n0_6054_19458 n2_6054_19458 0.0
V18666 n0_6054_19472 n2_6054_19472 0.0
V18667 n0_6054_19641 n2_6054_19641 0.0
V18668 n0_6054_19674 n2_6054_19674 0.0
V18669 n0_6054_19857 n2_6054_19857 0.0
V18670 n0_6054_19890 n2_6054_19890 0.0
V18671 n0_6054_20073 n2_6054_20073 0.0
V18672 n0_6054_20106 n2_6054_20106 0.0
V18673 n0_6054_20289 n2_6054_20289 0.0
V18674 n0_6054_20322 n2_6054_20322 0.0
V18675 n0_6054_20505 n2_6054_20505 0.0
V18676 n0_6054_20538 n2_6054_20538 0.0
V18677 n0_6054_20721 n2_6054_20721 0.0
V18678 n0_6054_20754 n2_6054_20754 0.0
V18679 n0_6054_20937 n2_6054_20937 0.0
V18680 n0_6054_20970 n2_6054_20970 0.0
V18681 n0_6146_201 n2_6146_201 0.0
V18682 n0_6146_234 n2_6146_234 0.0
V18683 n0_6146_356 n2_6146_356 0.0
V18684 n0_6146_417 n2_6146_417 0.0
V18685 n0_6146_450 n2_6146_450 0.0
V18686 n0_6146_633 n2_6146_633 0.0
V18687 n0_6146_666 n2_6146_666 0.0
V18688 n0_6146_788 n2_6146_788 0.0
V18689 n0_6146_849 n2_6146_849 0.0
V18690 n0_6146_882 n2_6146_882 0.0
V18691 n0_6146_1065 n2_6146_1065 0.0
V18692 n0_6146_1098 n2_6146_1098 0.0
V18693 n0_6146_1281 n2_6146_1281 0.0
V18694 n0_6146_1314 n2_6146_1314 0.0
V18695 n0_6146_1497 n2_6146_1497 0.0
V18696 n0_6146_1530 n2_6146_1530 0.0
V18697 n0_6146_1713 n2_6146_1713 0.0
V18698 n0_6146_1746 n2_6146_1746 0.0
V18699 n0_6146_1760 n2_6146_1760 0.0
V18700 n0_6146_1929 n2_6146_1929 0.0
V18701 n0_6146_1962 n2_6146_1962 0.0
V18702 n0_6146_2145 n2_6146_2145 0.0
V18703 n0_6146_2178 n2_6146_2178 0.0
V18704 n0_6146_2361 n2_6146_2361 0.0
V18705 n0_6146_2394 n2_6146_2394 0.0
V18706 n0_6146_2408 n2_6146_2408 0.0
V18707 n0_6146_2577 n2_6146_2577 0.0
V18708 n0_6146_2610 n2_6146_2610 0.0
V18709 n0_6146_2793 n2_6146_2793 0.0
V18710 n0_6146_2826 n2_6146_2826 0.0
V18711 n0_6146_2840 n2_6146_2840 0.0
V18712 n0_6146_3009 n2_6146_3009 0.0
V18713 n0_6146_3042 n2_6146_3042 0.0
V18714 n0_6146_3056 n2_6146_3056 0.0
V18715 n0_6146_3225 n2_6146_3225 0.0
V18716 n0_6146_3258 n2_6146_3258 0.0
V18717 n0_6146_3441 n2_6146_3441 0.0
V18718 n0_6146_3474 n2_6146_3474 0.0
V18719 n0_6146_3488 n2_6146_3488 0.0
V18720 n0_6146_3657 n2_6146_3657 0.0
V18721 n0_6146_3690 n2_6146_3690 0.0
V18722 n0_6146_3873 n2_6146_3873 0.0
V18723 n0_6146_3906 n2_6146_3906 0.0
V18724 n0_6146_4089 n2_6146_4089 0.0
V18725 n0_6146_4122 n2_6146_4122 0.0
V18726 n0_6146_4136 n2_6146_4136 0.0
V18727 n0_6146_4305 n2_6146_4305 0.0
V18728 n0_6146_4338 n2_6146_4338 0.0
V18729 n0_6146_4352 n2_6146_4352 0.0
V18730 n0_6146_4375 n2_6146_4375 0.0
V18731 n0_6146_4521 n2_6146_4521 0.0
V18732 n0_6146_4554 n2_6146_4554 0.0
V18733 n0_6146_4568 n2_6146_4568 0.0
V18734 n0_6146_4737 n2_6146_4737 0.0
V18735 n0_6146_4770 n2_6146_4770 0.0
V18736 n0_6146_4953 n2_6146_4953 0.0
V18737 n0_6146_5169 n2_6146_5169 0.0
V18738 n0_6146_5202 n2_6146_5202 0.0
V18739 n0_6146_5216 n2_6146_5216 0.0
V18740 n0_6146_5385 n2_6146_5385 0.0
V18741 n0_6146_5418 n2_6146_5418 0.0
V18742 n0_6146_5432 n2_6146_5432 0.0
V18743 n0_6146_5455 n2_6146_5455 0.0
V18744 n0_6146_5601 n2_6146_5601 0.0
V18745 n0_6146_5634 n2_6146_5634 0.0
V18746 n0_6146_5817 n2_6146_5817 0.0
V18747 n0_6146_5850 n2_6146_5850 0.0
V18748 n0_6146_6033 n2_6146_6033 0.0
V18749 n0_6146_6066 n2_6146_6066 0.0
V18750 n0_6146_15138 n2_6146_15138 0.0
V18751 n0_6146_15321 n2_6146_15321 0.0
V18752 n0_6146_15354 n2_6146_15354 0.0
V18753 n0_6146_15537 n2_6146_15537 0.0
V18754 n0_6146_15570 n2_6146_15570 0.0
V18755 n0_6146_15584 n2_6146_15584 0.0
V18756 n0_6146_15753 n2_6146_15753 0.0
V18757 n0_6146_15786 n2_6146_15786 0.0
V18758 n0_6146_15800 n2_6146_15800 0.0
V18759 n0_6146_15969 n2_6146_15969 0.0
V18760 n0_6146_16002 n2_6146_16002 0.0
V18761 n0_6146_16016 n2_6146_16016 0.0
V18762 n0_6146_16185 n2_6146_16185 0.0
V18763 n0_6146_16401 n2_6146_16401 0.0
V18764 n0_6146_16434 n2_6146_16434 0.0
V18765 n0_6146_16617 n2_6146_16617 0.0
V18766 n0_6146_16650 n2_6146_16650 0.0
V18767 n0_6146_16833 n2_6146_16833 0.0
V18768 n0_6146_16866 n2_6146_16866 0.0
V18769 n0_6146_17049 n2_6146_17049 0.0
V18770 n0_6146_17082 n2_6146_17082 0.0
V18771 n0_6146_17096 n2_6146_17096 0.0
V18772 n0_6146_17119 n2_6146_17119 0.0
V18773 n0_6146_17265 n2_6146_17265 0.0
V18774 n0_6146_17298 n2_6146_17298 0.0
V18775 n0_6146_17312 n2_6146_17312 0.0
V18776 n0_6146_17481 n2_6146_17481 0.0
V18777 n0_6146_17514 n2_6146_17514 0.0
V18778 n0_6146_17528 n2_6146_17528 0.0
V18779 n0_6146_17697 n2_6146_17697 0.0
V18780 n0_6146_17730 n2_6146_17730 0.0
V18781 n0_6146_17913 n2_6146_17913 0.0
V18782 n0_6146_17946 n2_6146_17946 0.0
V18783 n0_6146_18129 n2_6146_18129 0.0
V18784 n0_6146_18162 n2_6146_18162 0.0
V18785 n0_6146_18345 n2_6146_18345 0.0
V18786 n0_6146_18378 n2_6146_18378 0.0
V18787 n0_6146_18392 n2_6146_18392 0.0
V18788 n0_6146_18561 n2_6146_18561 0.0
V18789 n0_6146_18594 n2_6146_18594 0.0
V18790 n0_6146_18608 n2_6146_18608 0.0
V18791 n0_6146_18777 n2_6146_18777 0.0
V18792 n0_6146_18810 n2_6146_18810 0.0
V18793 n0_6146_18824 n2_6146_18824 0.0
V18794 n0_6146_18993 n2_6146_18993 0.0
V18795 n0_6146_19026 n2_6146_19026 0.0
V18796 n0_6146_19040 n2_6146_19040 0.0
V18797 n0_6146_19209 n2_6146_19209 0.0
V18798 n0_6146_19242 n2_6146_19242 0.0
V18799 n0_6146_19425 n2_6146_19425 0.0
V18800 n0_6146_19458 n2_6146_19458 0.0
V18801 n0_6146_19472 n2_6146_19472 0.0
V18802 n0_6146_19641 n2_6146_19641 0.0
V18803 n0_6146_19674 n2_6146_19674 0.0
V18804 n0_6146_19857 n2_6146_19857 0.0
V18805 n0_6146_19890 n2_6146_19890 0.0
V18806 n0_6146_20073 n2_6146_20073 0.0
V18807 n0_6146_20106 n2_6146_20106 0.0
V18808 n0_6146_20289 n2_6146_20289 0.0
V18809 n0_6146_20322 n2_6146_20322 0.0
V18810 n0_6146_20505 n2_6146_20505 0.0
V18811 n0_6146_20538 n2_6146_20538 0.0
V18812 n0_6146_20754 n2_6146_20754 0.0
V18813 n0_6146_20937 n2_6146_20937 0.0
V18814 n0_6146_20970 n2_6146_20970 0.0
V18815 n0_6991_7329 n2_6991_7329 0.0
V18816 n0_6991_7362 n2_6991_7362 0.0
V18817 n0_6991_7545 n2_6991_7545 0.0
V18818 n0_6991_7578 n2_6991_7578 0.0
V18819 n0_6991_7761 n2_6991_7761 0.0
V18820 n0_6991_7794 n2_6991_7794 0.0
V18821 n0_6991_7808 n2_6991_7808 0.0
V18822 n0_6991_7977 n2_6991_7977 0.0
V18823 n0_6991_8010 n2_6991_8010 0.0
V18824 n0_6991_8193 n2_6991_8193 0.0
V18825 n0_6991_8226 n2_6991_8226 0.0
V18826 n0_6991_8409 n2_6991_8409 0.0
V18827 n0_6991_8442 n2_6991_8442 0.0
V18828 n0_6991_8625 n2_6991_8625 0.0
V18829 n0_6991_8658 n2_6991_8658 0.0
V18830 n0_6991_8841 n2_6991_8841 0.0
V18831 n0_6991_8874 n2_6991_8874 0.0
V18832 n0_6991_8888 n2_6991_8888 0.0
V18833 n0_6991_9057 n2_6991_9057 0.0
V18834 n0_6991_9090 n2_6991_9090 0.0
V18835 n0_6991_9273 n2_6991_9273 0.0
V18836 n0_6991_9306 n2_6991_9306 0.0
V18837 n0_6991_9489 n2_6991_9489 0.0
V18838 n0_6991_9522 n2_6991_9522 0.0
V18839 n0_6991_9705 n2_6991_9705 0.0
V18840 n0_6991_9738 n2_6991_9738 0.0
V18841 n0_6991_9921 n2_6991_9921 0.0
V18842 n0_6991_9954 n2_6991_9954 0.0
V18843 n0_6991_9968 n2_6991_9968 0.0
V18844 n0_6991_10137 n2_6991_10137 0.0
V18845 n0_6991_10170 n2_6991_10170 0.0
V18846 n0_6991_10353 n2_6991_10353 0.0
V18847 n0_6991_10386 n2_6991_10386 0.0
V18848 n0_6991_10569 n2_6991_10569 0.0
V18849 n0_6991_10785 n2_6991_10785 0.0
V18850 n0_6991_10818 n2_6991_10818 0.0
V18851 n0_6991_11001 n2_6991_11001 0.0
V18852 n0_6991_11034 n2_6991_11034 0.0
V18853 n0_6991_11048 n2_6991_11048 0.0
V18854 n0_6991_11217 n2_6991_11217 0.0
V18855 n0_6991_11250 n2_6991_11250 0.0
V18856 n0_6991_11433 n2_6991_11433 0.0
V18857 n0_6991_11466 n2_6991_11466 0.0
V18858 n0_6991_11649 n2_6991_11649 0.0
V18859 n0_6991_11682 n2_6991_11682 0.0
V18860 n0_6991_11865 n2_6991_11865 0.0
V18861 n0_6991_11898 n2_6991_11898 0.0
V18862 n0_6991_12081 n2_6991_12081 0.0
V18863 n0_6991_12114 n2_6991_12114 0.0
V18864 n0_6991_12128 n2_6991_12128 0.0
V18865 n0_6991_12297 n2_6991_12297 0.0
V18866 n0_6991_12330 n2_6991_12330 0.0
V18867 n0_6991_12513 n2_6991_12513 0.0
V18868 n0_6991_12546 n2_6991_12546 0.0
V18869 n0_6991_12729 n2_6991_12729 0.0
V18870 n0_6991_12762 n2_6991_12762 0.0
V18871 n0_6991_12945 n2_6991_12945 0.0
V18872 n0_6991_12978 n2_6991_12978 0.0
V18873 n0_6991_13161 n2_6991_13161 0.0
V18874 n0_6991_13194 n2_6991_13194 0.0
V18875 n0_6991_13377 n2_6991_13377 0.0
V18876 n0_6991_13410 n2_6991_13410 0.0
V18877 n0_6991_13424 n2_6991_13424 0.0
V18878 n0_6991_13593 n2_6991_13593 0.0
V18879 n0_6991_13626 n2_6991_13626 0.0
V18880 n0_6991_13809 n2_6991_13809 0.0
V18881 n0_6991_13842 n2_6991_13842 0.0
V18882 n0_7130_8409 n2_7130_8409 0.0
V18883 n0_7130_10569 n2_7130_10569 0.0
V18884 n0_7130_10602 n2_7130_10602 0.0
V18885 n0_7179_7329 n2_7179_7329 0.0
V18886 n0_7179_7362 n2_7179_7362 0.0
V18887 n0_7179_7545 n2_7179_7545 0.0
V18888 n0_7179_7578 n2_7179_7578 0.0
V18889 n0_7179_7761 n2_7179_7761 0.0
V18890 n0_7179_7794 n2_7179_7794 0.0
V18891 n0_7179_7808 n2_7179_7808 0.0
V18892 n0_7179_7977 n2_7179_7977 0.0
V18893 n0_7179_8010 n2_7179_8010 0.0
V18894 n0_7179_8193 n2_7179_8193 0.0
V18895 n0_7179_8226 n2_7179_8226 0.0
V18896 n0_7179_8409 n2_7179_8409 0.0
V18897 n0_7179_8442 n2_7179_8442 0.0
V18898 n0_7179_8625 n2_7179_8625 0.0
V18899 n0_7179_8658 n2_7179_8658 0.0
V18900 n0_7179_8841 n2_7179_8841 0.0
V18901 n0_7179_8874 n2_7179_8874 0.0
V18902 n0_7179_8888 n2_7179_8888 0.0
V18903 n0_7179_9057 n2_7179_9057 0.0
V18904 n0_7179_9090 n2_7179_9090 0.0
V18905 n0_7179_9273 n2_7179_9273 0.0
V18906 n0_7179_9306 n2_7179_9306 0.0
V18907 n0_7179_9705 n2_7179_9705 0.0
V18908 n0_7179_9738 n2_7179_9738 0.0
V18909 n0_7179_9921 n2_7179_9921 0.0
V18910 n0_7179_9954 n2_7179_9954 0.0
V18911 n0_7179_9968 n2_7179_9968 0.0
V18912 n0_7179_10137 n2_7179_10137 0.0
V18913 n0_7179_10170 n2_7179_10170 0.0
V18914 n0_7179_10353 n2_7179_10353 0.0
V18915 n0_7179_10386 n2_7179_10386 0.0
V18916 n0_7179_10569 n2_7179_10569 0.0
V18917 n0_7179_10602 n2_7179_10602 0.0
V18918 n0_7179_10785 n2_7179_10785 0.0
V18919 n0_7179_10818 n2_7179_10818 0.0
V18920 n0_7179_11001 n2_7179_11001 0.0
V18921 n0_7179_11034 n2_7179_11034 0.0
V18922 n0_7179_11048 n2_7179_11048 0.0
V18923 n0_7179_11217 n2_7179_11217 0.0
V18924 n0_7179_11250 n2_7179_11250 0.0
V18925 n0_7179_11433 n2_7179_11433 0.0
V18926 n0_7179_11466 n2_7179_11466 0.0
V18927 n0_7179_11865 n2_7179_11865 0.0
V18928 n0_7179_11898 n2_7179_11898 0.0
V18929 n0_7179_12081 n2_7179_12081 0.0
V18930 n0_7179_12114 n2_7179_12114 0.0
V18931 n0_7179_12128 n2_7179_12128 0.0
V18932 n0_7179_12297 n2_7179_12297 0.0
V18933 n0_7179_12330 n2_7179_12330 0.0
V18934 n0_7179_12513 n2_7179_12513 0.0
V18935 n0_7179_12546 n2_7179_12546 0.0
V18936 n0_7179_12729 n2_7179_12729 0.0
V18937 n0_7179_12762 n2_7179_12762 0.0
V18938 n0_7179_12945 n2_7179_12945 0.0
V18939 n0_7179_12978 n2_7179_12978 0.0
V18940 n0_7179_13161 n2_7179_13161 0.0
V18941 n0_7179_13194 n2_7179_13194 0.0
V18942 n0_7179_13377 n2_7179_13377 0.0
V18943 n0_7179_13410 n2_7179_13410 0.0
V18944 n0_7179_13424 n2_7179_13424 0.0
V18945 n0_7179_13593 n2_7179_13593 0.0
V18946 n0_7179_13626 n2_7179_13626 0.0
V18947 n0_7179_13809 n2_7179_13809 0.0
V18948 n0_7179_13842 n2_7179_13842 0.0
V18949 n0_8116_201 n2_8116_201 0.0
V18950 n0_8116_234 n2_8116_234 0.0
V18951 n0_8116_417 n2_8116_417 0.0
V18952 n0_8116_450 n2_8116_450 0.0
V18953 n0_8116_633 n2_8116_633 0.0
V18954 n0_8116_666 n2_8116_666 0.0
V18955 n0_8116_849 n2_8116_849 0.0
V18956 n0_8116_882 n2_8116_882 0.0
V18957 n0_8116_1065 n2_8116_1065 0.0
V18958 n0_8116_1098 n2_8116_1098 0.0
V18959 n0_8116_1281 n2_8116_1281 0.0
V18960 n0_8116_1314 n2_8116_1314 0.0
V18961 n0_8116_1497 n2_8116_1497 0.0
V18962 n0_8116_1530 n2_8116_1530 0.0
V18963 n0_8116_1713 n2_8116_1713 0.0
V18964 n0_8116_1746 n2_8116_1746 0.0
V18965 n0_8116_1760 n2_8116_1760 0.0
V18966 n0_8116_1783 n2_8116_1783 0.0
V18967 n0_8116_1929 n2_8116_1929 0.0
V18968 n0_8116_1962 n2_8116_1962 0.0
V18969 n0_8116_2145 n2_8116_2145 0.0
V18970 n0_8116_2178 n2_8116_2178 0.0
V18971 n0_8116_2361 n2_8116_2361 0.0
V18972 n0_8116_2394 n2_8116_2394 0.0
V18973 n0_8116_2408 n2_8116_2408 0.0
V18974 n0_8116_2577 n2_8116_2577 0.0
V18975 n0_8116_2610 n2_8116_2610 0.0
V18976 n0_8116_2793 n2_8116_2793 0.0
V18977 n0_8116_2826 n2_8116_2826 0.0
V18978 n0_8116_2840 n2_8116_2840 0.0
V18979 n0_8116_2863 n2_8116_2863 0.0
V18980 n0_8116_3009 n2_8116_3009 0.0
V18981 n0_8116_3042 n2_8116_3042 0.0
V18982 n0_8116_3225 n2_8116_3225 0.0
V18983 n0_8116_3258 n2_8116_3258 0.0
V18984 n0_8116_3441 n2_8116_3441 0.0
V18985 n0_8116_3474 n2_8116_3474 0.0
V18986 n0_8116_3488 n2_8116_3488 0.0
V18987 n0_8116_3657 n2_8116_3657 0.0
V18988 n0_8116_3690 n2_8116_3690 0.0
V18989 n0_8116_3873 n2_8116_3873 0.0
V18990 n0_8116_3906 n2_8116_3906 0.0
V18991 n0_8116_4089 n2_8116_4089 0.0
V18992 n0_8116_4122 n2_8116_4122 0.0
V18993 n0_8116_4136 n2_8116_4136 0.0
V18994 n0_8116_4305 n2_8116_4305 0.0
V18995 n0_8116_4338 n2_8116_4338 0.0
V18996 n0_8116_4521 n2_8116_4521 0.0
V18997 n0_8116_4554 n2_8116_4554 0.0
V18998 n0_8116_4568 n2_8116_4568 0.0
V18999 n0_8116_4737 n2_8116_4737 0.0
V19000 n0_8116_4770 n2_8116_4770 0.0
V19001 n0_8116_4953 n2_8116_4953 0.0
V19002 n0_8116_5169 n2_8116_5169 0.0
V19003 n0_8116_5202 n2_8116_5202 0.0
V19004 n0_8116_5216 n2_8116_5216 0.0
V19005 n0_8116_5239 n2_8116_5239 0.0
V19006 n0_8116_5385 n2_8116_5385 0.0
V19007 n0_8116_5418 n2_8116_5418 0.0
V19008 n0_8116_5432 n2_8116_5432 0.0
V19009 n0_8116_5455 n2_8116_5455 0.0
V19010 n0_8116_5601 n2_8116_5601 0.0
V19011 n0_8116_5634 n2_8116_5634 0.0
V19012 n0_8116_5817 n2_8116_5817 0.0
V19013 n0_8116_5850 n2_8116_5850 0.0
V19014 n0_8116_6033 n2_8116_6033 0.0
V19015 n0_8116_6066 n2_8116_6066 0.0
V19016 n0_8116_6249 n2_8116_6249 0.0
V19017 n0_8116_6282 n2_8116_6282 0.0
V19018 n0_8116_6465 n2_8116_6465 0.0
V19019 n0_8116_6498 n2_8116_6498 0.0
V19020 n0_8116_6512 n2_8116_6512 0.0
V19021 n0_8116_6535 n2_8116_6535 0.0
V19022 n0_8116_6681 n2_8116_6681 0.0
V19023 n0_8116_6714 n2_8116_6714 0.0
V19024 n0_8116_6897 n2_8116_6897 0.0
V19025 n0_8116_6930 n2_8116_6930 0.0
V19026 n0_8116_6944 n2_8116_6944 0.0
V19027 n0_8116_7113 n2_8116_7113 0.0
V19028 n0_8116_7146 n2_8116_7146 0.0
V19029 n0_8116_7160 n2_8116_7160 0.0
V19030 n0_8116_7329 n2_8116_7329 0.0
V19031 n0_8116_7362 n2_8116_7362 0.0
V19032 n0_8116_7376 n2_8116_7376 0.0
V19033 n0_8116_7545 n2_8116_7545 0.0
V19034 n0_8116_7578 n2_8116_7578 0.0
V19035 n0_8116_7761 n2_8116_7761 0.0
V19036 n0_8116_7794 n2_8116_7794 0.0
V19037 n0_8116_7808 n2_8116_7808 0.0
V19038 n0_8116_7977 n2_8116_7977 0.0
V19039 n0_8116_8010 n2_8116_8010 0.0
V19040 n0_8116_8193 n2_8116_8193 0.0
V19041 n0_8116_8226 n2_8116_8226 0.0
V19042 n0_8116_8409 n2_8116_8409 0.0
V19043 n0_8116_8442 n2_8116_8442 0.0
V19044 n0_8116_8625 n2_8116_8625 0.0
V19045 n0_8116_8658 n2_8116_8658 0.0
V19046 n0_8116_8841 n2_8116_8841 0.0
V19047 n0_8116_8874 n2_8116_8874 0.0
V19048 n0_8116_8888 n2_8116_8888 0.0
V19049 n0_8116_9057 n2_8116_9057 0.0
V19050 n0_8116_9090 n2_8116_9090 0.0
V19051 n0_8116_9273 n2_8116_9273 0.0
V19052 n0_8116_9306 n2_8116_9306 0.0
V19053 n0_8116_9489 n2_8116_9489 0.0
V19054 n0_8116_9522 n2_8116_9522 0.0
V19055 n0_8116_9705 n2_8116_9705 0.0
V19056 n0_8116_9738 n2_8116_9738 0.0
V19057 n0_8116_9921 n2_8116_9921 0.0
V19058 n0_8116_9954 n2_8116_9954 0.0
V19059 n0_8116_9968 n2_8116_9968 0.0
V19060 n0_8116_10137 n2_8116_10137 0.0
V19061 n0_8116_10170 n2_8116_10170 0.0
V19062 n0_8116_10353 n2_8116_10353 0.0
V19063 n0_8116_10386 n2_8116_10386 0.0
V19064 n0_8116_10569 n2_8116_10569 0.0
V19065 n0_8116_10785 n2_8116_10785 0.0
V19066 n0_8116_10818 n2_8116_10818 0.0
V19067 n0_8116_11001 n2_8116_11001 0.0
V19068 n0_8116_11034 n2_8116_11034 0.0
V19069 n0_8116_11048 n2_8116_11048 0.0
V19070 n0_8116_11217 n2_8116_11217 0.0
V19071 n0_8116_11250 n2_8116_11250 0.0
V19072 n0_8116_11433 n2_8116_11433 0.0
V19073 n0_8116_11466 n2_8116_11466 0.0
V19074 n0_8116_11649 n2_8116_11649 0.0
V19075 n0_8116_11682 n2_8116_11682 0.0
V19076 n0_8116_11865 n2_8116_11865 0.0
V19077 n0_8116_11898 n2_8116_11898 0.0
V19078 n0_8116_12081 n2_8116_12081 0.0
V19079 n0_8116_12114 n2_8116_12114 0.0
V19080 n0_8116_12128 n2_8116_12128 0.0
V19081 n0_8116_12297 n2_8116_12297 0.0
V19082 n0_8116_12330 n2_8116_12330 0.0
V19083 n0_8116_12513 n2_8116_12513 0.0
V19084 n0_8116_12546 n2_8116_12546 0.0
V19085 n0_8116_12729 n2_8116_12729 0.0
V19086 n0_8116_12762 n2_8116_12762 0.0
V19087 n0_8116_12945 n2_8116_12945 0.0
V19088 n0_8116_12978 n2_8116_12978 0.0
V19089 n0_8116_13161 n2_8116_13161 0.0
V19090 n0_8116_13194 n2_8116_13194 0.0
V19091 n0_8116_13377 n2_8116_13377 0.0
V19092 n0_8116_13410 n2_8116_13410 0.0
V19093 n0_8116_13424 n2_8116_13424 0.0
V19094 n0_8116_13593 n2_8116_13593 0.0
V19095 n0_8116_13626 n2_8116_13626 0.0
V19096 n0_8116_13640 n2_8116_13640 0.0
V19097 n0_8116_13809 n2_8116_13809 0.0
V19098 n0_8116_13842 n2_8116_13842 0.0
V19099 n0_8116_13856 n2_8116_13856 0.0
V19100 n0_8116_14025 n2_8116_14025 0.0
V19101 n0_8116_14058 n2_8116_14058 0.0
V19102 n0_8116_14072 n2_8116_14072 0.0
V19103 n0_8116_14241 n2_8116_14241 0.0
V19104 n0_8116_14274 n2_8116_14274 0.0
V19105 n0_8116_14396 n2_8116_14396 0.0
V19106 n0_8116_14457 n2_8116_14457 0.0
V19107 n0_8116_14490 n2_8116_14490 0.0
V19108 n0_8116_14504 n2_8116_14504 0.0
V19109 n0_8116_14673 n2_8116_14673 0.0
V19110 n0_8116_14706 n2_8116_14706 0.0
V19111 n0_8116_14889 n2_8116_14889 0.0
V19112 n0_8116_14922 n2_8116_14922 0.0
V19113 n0_8116_15138 n2_8116_15138 0.0
V19114 n0_8116_15321 n2_8116_15321 0.0
V19115 n0_8116_15354 n2_8116_15354 0.0
V19116 n0_8116_15537 n2_8116_15537 0.0
V19117 n0_8116_15570 n2_8116_15570 0.0
V19118 n0_8116_15584 n2_8116_15584 0.0
V19119 n0_8116_15753 n2_8116_15753 0.0
V19120 n0_8116_15786 n2_8116_15786 0.0
V19121 n0_8116_15800 n2_8116_15800 0.0
V19122 n0_8116_15969 n2_8116_15969 0.0
V19123 n0_8116_16002 n2_8116_16002 0.0
V19124 n0_8116_16016 n2_8116_16016 0.0
V19125 n0_8116_16185 n2_8116_16185 0.0
V19126 n0_8116_16401 n2_8116_16401 0.0
V19127 n0_8116_16434 n2_8116_16434 0.0
V19128 n0_8116_16617 n2_8116_16617 0.0
V19129 n0_8116_16650 n2_8116_16650 0.0
V19130 n0_8116_16833 n2_8116_16833 0.0
V19131 n0_8116_16866 n2_8116_16866 0.0
V19132 n0_8116_17049 n2_8116_17049 0.0
V19133 n0_8116_17082 n2_8116_17082 0.0
V19134 n0_8116_17096 n2_8116_17096 0.0
V19135 n0_8116_17119 n2_8116_17119 0.0
V19136 n0_8116_17265 n2_8116_17265 0.0
V19137 n0_8116_17298 n2_8116_17298 0.0
V19138 n0_8116_17312 n2_8116_17312 0.0
V19139 n0_8116_17481 n2_8116_17481 0.0
V19140 n0_8116_17514 n2_8116_17514 0.0
V19141 n0_8116_17697 n2_8116_17697 0.0
V19142 n0_8116_17730 n2_8116_17730 0.0
V19143 n0_8116_17913 n2_8116_17913 0.0
V19144 n0_8116_17946 n2_8116_17946 0.0
V19145 n0_8116_18129 n2_8116_18129 0.0
V19146 n0_8116_18162 n2_8116_18162 0.0
V19147 n0_8116_18345 n2_8116_18345 0.0
V19148 n0_8116_18378 n2_8116_18378 0.0
V19149 n0_8116_18392 n2_8116_18392 0.0
V19150 n0_8116_18421 n2_8116_18421 0.0
V19151 n0_8116_18561 n2_8116_18561 0.0
V19152 n0_8116_18594 n2_8116_18594 0.0
V19153 n0_8116_18608 n2_8116_18608 0.0
V19154 n0_8116_18777 n2_8116_18777 0.0
V19155 n0_8116_18810 n2_8116_18810 0.0
V19156 n0_8116_18993 n2_8116_18993 0.0
V19157 n0_8116_19026 n2_8116_19026 0.0
V19158 n0_8116_19209 n2_8116_19209 0.0
V19159 n0_8116_19242 n2_8116_19242 0.0
V19160 n0_8116_19256 n2_8116_19256 0.0
V19161 n0_8116_19279 n2_8116_19279 0.0
V19162 n0_8116_19425 n2_8116_19425 0.0
V19163 n0_8116_19458 n2_8116_19458 0.0
V19164 n0_8116_19641 n2_8116_19641 0.0
V19165 n0_8116_19674 n2_8116_19674 0.0
V19166 n0_8116_19857 n2_8116_19857 0.0
V19167 n0_8116_19890 n2_8116_19890 0.0
V19168 n0_8116_20073 n2_8116_20073 0.0
V19169 n0_8116_20106 n2_8116_20106 0.0
V19170 n0_8116_20289 n2_8116_20289 0.0
V19171 n0_8116_20322 n2_8116_20322 0.0
V19172 n0_8116_20505 n2_8116_20505 0.0
V19173 n0_8116_20538 n2_8116_20538 0.0
V19174 n0_8116_20754 n2_8116_20754 0.0
V19175 n0_8116_20937 n2_8116_20937 0.0
V19176 n0_8116_20970 n2_8116_20970 0.0
V19177 n0_8208_201 n2_8208_201 0.0
V19178 n0_8208_234 n2_8208_234 0.0
V19179 n0_8208_417 n2_8208_417 0.0
V19180 n0_8208_450 n2_8208_450 0.0
V19181 n0_8208_633 n2_8208_633 0.0
V19182 n0_8208_666 n2_8208_666 0.0
V19183 n0_8208_849 n2_8208_849 0.0
V19184 n0_8208_882 n2_8208_882 0.0
V19185 n0_8208_1065 n2_8208_1065 0.0
V19186 n0_8208_1098 n2_8208_1098 0.0
V19187 n0_8208_1281 n2_8208_1281 0.0
V19188 n0_8208_1314 n2_8208_1314 0.0
V19189 n0_8208_1497 n2_8208_1497 0.0
V19190 n0_8208_1530 n2_8208_1530 0.0
V19191 n0_8208_1713 n2_8208_1713 0.0
V19192 n0_8208_1746 n2_8208_1746 0.0
V19193 n0_8208_1760 n2_8208_1760 0.0
V19194 n0_8208_1783 n2_8208_1783 0.0
V19195 n0_8208_1929 n2_8208_1929 0.0
V19196 n0_8208_1962 n2_8208_1962 0.0
V19197 n0_8208_2145 n2_8208_2145 0.0
V19198 n0_8208_2178 n2_8208_2178 0.0
V19199 n0_8208_2361 n2_8208_2361 0.0
V19200 n0_8208_2394 n2_8208_2394 0.0
V19201 n0_8208_2408 n2_8208_2408 0.0
V19202 n0_8208_2577 n2_8208_2577 0.0
V19203 n0_8208_2610 n2_8208_2610 0.0
V19204 n0_8208_2793 n2_8208_2793 0.0
V19205 n0_8208_2826 n2_8208_2826 0.0
V19206 n0_8208_2840 n2_8208_2840 0.0
V19207 n0_8208_2863 n2_8208_2863 0.0
V19208 n0_8208_3009 n2_8208_3009 0.0
V19209 n0_8208_3042 n2_8208_3042 0.0
V19210 n0_8208_3225 n2_8208_3225 0.0
V19211 n0_8208_3258 n2_8208_3258 0.0
V19212 n0_8208_3441 n2_8208_3441 0.0
V19213 n0_8208_3474 n2_8208_3474 0.0
V19214 n0_8208_3488 n2_8208_3488 0.0
V19215 n0_8208_3657 n2_8208_3657 0.0
V19216 n0_8208_3690 n2_8208_3690 0.0
V19217 n0_8208_3873 n2_8208_3873 0.0
V19218 n0_8208_3906 n2_8208_3906 0.0
V19219 n0_8208_4089 n2_8208_4089 0.0
V19220 n0_8208_4122 n2_8208_4122 0.0
V19221 n0_8208_4136 n2_8208_4136 0.0
V19222 n0_8208_4305 n2_8208_4305 0.0
V19223 n0_8208_4338 n2_8208_4338 0.0
V19224 n0_8208_4521 n2_8208_4521 0.0
V19225 n0_8208_4554 n2_8208_4554 0.0
V19226 n0_8208_4568 n2_8208_4568 0.0
V19227 n0_8208_4737 n2_8208_4737 0.0
V19228 n0_8208_4770 n2_8208_4770 0.0
V19229 n0_8208_4953 n2_8208_4953 0.0
V19230 n0_8208_4986 n2_8208_4986 0.0
V19231 n0_8208_5169 n2_8208_5169 0.0
V19232 n0_8208_5202 n2_8208_5202 0.0
V19233 n0_8208_5216 n2_8208_5216 0.0
V19234 n0_8208_5239 n2_8208_5239 0.0
V19235 n0_8208_5385 n2_8208_5385 0.0
V19236 n0_8208_5418 n2_8208_5418 0.0
V19237 n0_8208_5432 n2_8208_5432 0.0
V19238 n0_8208_5455 n2_8208_5455 0.0
V19239 n0_8208_5601 n2_8208_5601 0.0
V19240 n0_8208_5634 n2_8208_5634 0.0
V19241 n0_8208_5817 n2_8208_5817 0.0
V19242 n0_8208_5850 n2_8208_5850 0.0
V19243 n0_8208_6033 n2_8208_6033 0.0
V19244 n0_8208_6066 n2_8208_6066 0.0
V19245 n0_8208_6249 n2_8208_6249 0.0
V19246 n0_8208_6282 n2_8208_6282 0.0
V19247 n0_8208_6465 n2_8208_6465 0.0
V19248 n0_8208_6498 n2_8208_6498 0.0
V19249 n0_8208_6512 n2_8208_6512 0.0
V19250 n0_8208_6535 n2_8208_6535 0.0
V19251 n0_8208_6681 n2_8208_6681 0.0
V19252 n0_8208_6714 n2_8208_6714 0.0
V19253 n0_8208_6897 n2_8208_6897 0.0
V19254 n0_8208_6930 n2_8208_6930 0.0
V19255 n0_8208_6944 n2_8208_6944 0.0
V19256 n0_8208_7113 n2_8208_7113 0.0
V19257 n0_8208_7146 n2_8208_7146 0.0
V19258 n0_8208_7160 n2_8208_7160 0.0
V19259 n0_8208_7329 n2_8208_7329 0.0
V19260 n0_8208_7362 n2_8208_7362 0.0
V19261 n0_8208_7376 n2_8208_7376 0.0
V19262 n0_8208_7545 n2_8208_7545 0.0
V19263 n0_8208_7578 n2_8208_7578 0.0
V19264 n0_8208_7761 n2_8208_7761 0.0
V19265 n0_8208_7794 n2_8208_7794 0.0
V19266 n0_8208_7808 n2_8208_7808 0.0
V19267 n0_8208_7977 n2_8208_7977 0.0
V19268 n0_8208_8010 n2_8208_8010 0.0
V19269 n0_8208_8193 n2_8208_8193 0.0
V19270 n0_8208_8226 n2_8208_8226 0.0
V19271 n0_8208_8409 n2_8208_8409 0.0
V19272 n0_8208_8442 n2_8208_8442 0.0
V19273 n0_8208_12762 n2_8208_12762 0.0
V19274 n0_8208_12945 n2_8208_12945 0.0
V19275 n0_8208_12978 n2_8208_12978 0.0
V19276 n0_8208_13161 n2_8208_13161 0.0
V19277 n0_8208_13194 n2_8208_13194 0.0
V19278 n0_8208_13377 n2_8208_13377 0.0
V19279 n0_8208_13410 n2_8208_13410 0.0
V19280 n0_8208_13424 n2_8208_13424 0.0
V19281 n0_8208_13593 n2_8208_13593 0.0
V19282 n0_8208_13626 n2_8208_13626 0.0
V19283 n0_8208_13640 n2_8208_13640 0.0
V19284 n0_8208_13809 n2_8208_13809 0.0
V19285 n0_8208_13842 n2_8208_13842 0.0
V19286 n0_8208_13856 n2_8208_13856 0.0
V19287 n0_8208_14025 n2_8208_14025 0.0
V19288 n0_8208_14058 n2_8208_14058 0.0
V19289 n0_8208_14072 n2_8208_14072 0.0
V19290 n0_8208_14241 n2_8208_14241 0.0
V19291 n0_8208_14274 n2_8208_14274 0.0
V19292 n0_8208_14396 n2_8208_14396 0.0
V19293 n0_8208_14457 n2_8208_14457 0.0
V19294 n0_8208_14490 n2_8208_14490 0.0
V19295 n0_8208_14504 n2_8208_14504 0.0
V19296 n0_8208_14673 n2_8208_14673 0.0
V19297 n0_8208_14706 n2_8208_14706 0.0
V19298 n0_8208_14889 n2_8208_14889 0.0
V19299 n0_8208_14922 n2_8208_14922 0.0
V19300 n0_8208_15105 n2_8208_15105 0.0
V19301 n0_8208_15138 n2_8208_15138 0.0
V19302 n0_8208_15321 n2_8208_15321 0.0
V19303 n0_8208_15354 n2_8208_15354 0.0
V19304 n0_8208_15537 n2_8208_15537 0.0
V19305 n0_8208_15570 n2_8208_15570 0.0
V19306 n0_8208_15584 n2_8208_15584 0.0
V19307 n0_8208_15753 n2_8208_15753 0.0
V19308 n0_8208_15786 n2_8208_15786 0.0
V19309 n0_8208_15800 n2_8208_15800 0.0
V19310 n0_8208_15969 n2_8208_15969 0.0
V19311 n0_8208_16002 n2_8208_16002 0.0
V19312 n0_8208_16016 n2_8208_16016 0.0
V19313 n0_8208_16185 n2_8208_16185 0.0
V19314 n0_8208_16218 n2_8208_16218 0.0
V19315 n0_8208_16401 n2_8208_16401 0.0
V19316 n0_8208_16434 n2_8208_16434 0.0
V19317 n0_8208_16617 n2_8208_16617 0.0
V19318 n0_8208_16650 n2_8208_16650 0.0
V19319 n0_8208_16833 n2_8208_16833 0.0
V19320 n0_8208_16866 n2_8208_16866 0.0
V19321 n0_8208_17049 n2_8208_17049 0.0
V19322 n0_8208_17082 n2_8208_17082 0.0
V19323 n0_8208_17096 n2_8208_17096 0.0
V19324 n0_8208_17119 n2_8208_17119 0.0
V19325 n0_8208_17265 n2_8208_17265 0.0
V19326 n0_8208_17298 n2_8208_17298 0.0
V19327 n0_8208_17312 n2_8208_17312 0.0
V19328 n0_8208_17481 n2_8208_17481 0.0
V19329 n0_8208_17514 n2_8208_17514 0.0
V19330 n0_8208_17697 n2_8208_17697 0.0
V19331 n0_8208_17730 n2_8208_17730 0.0
V19332 n0_8208_17913 n2_8208_17913 0.0
V19333 n0_8208_17946 n2_8208_17946 0.0
V19334 n0_8208_18129 n2_8208_18129 0.0
V19335 n0_8208_18162 n2_8208_18162 0.0
V19336 n0_8208_18345 n2_8208_18345 0.0
V19337 n0_8208_18378 n2_8208_18378 0.0
V19338 n0_8208_18392 n2_8208_18392 0.0
V19339 n0_8208_18421 n2_8208_18421 0.0
V19340 n0_8208_18561 n2_8208_18561 0.0
V19341 n0_8208_18594 n2_8208_18594 0.0
V19342 n0_8208_18608 n2_8208_18608 0.0
V19343 n0_8208_18777 n2_8208_18777 0.0
V19344 n0_8208_18810 n2_8208_18810 0.0
V19345 n0_8208_18993 n2_8208_18993 0.0
V19346 n0_8208_19026 n2_8208_19026 0.0
V19347 n0_8208_19209 n2_8208_19209 0.0
V19348 n0_8208_19242 n2_8208_19242 0.0
V19349 n0_8208_19256 n2_8208_19256 0.0
V19350 n0_8208_19279 n2_8208_19279 0.0
V19351 n0_8208_19425 n2_8208_19425 0.0
V19352 n0_8208_19458 n2_8208_19458 0.0
V19353 n0_8208_19641 n2_8208_19641 0.0
V19354 n0_8208_19674 n2_8208_19674 0.0
V19355 n0_8208_19857 n2_8208_19857 0.0
V19356 n0_8208_19890 n2_8208_19890 0.0
V19357 n0_8208_20073 n2_8208_20073 0.0
V19358 n0_8208_20106 n2_8208_20106 0.0
V19359 n0_8208_20289 n2_8208_20289 0.0
V19360 n0_8208_20322 n2_8208_20322 0.0
V19361 n0_8208_20505 n2_8208_20505 0.0
V19362 n0_8208_20538 n2_8208_20538 0.0
V19363 n0_8208_20721 n2_8208_20721 0.0
V19364 n0_8208_20754 n2_8208_20754 0.0
V19365 n0_8208_20937 n2_8208_20937 0.0
V19366 n0_8208_20970 n2_8208_20970 0.0
V19367 n0_8255_417 n2_8255_417 0.0
V19368 n0_8255_450 n2_8255_450 0.0
V19369 n0_8255_1530 n2_8255_1530 0.0
V19370 n0_8255_2793 n2_8255_2793 0.0
V19371 n0_8255_3873 n2_8255_3873 0.0
V19372 n0_8255_3906 n2_8255_3906 0.0
V19373 n0_8255_4953 n2_8255_4953 0.0
V19374 n0_8255_4986 n2_8255_4986 0.0
V19375 n0_8255_6033 n2_8255_6033 0.0
V19376 n0_8255_6066 n2_8255_6066 0.0
V19377 n0_8255_7146 n2_8255_7146 0.0
V19378 n0_8255_7160 n2_8255_7160 0.0
V19379 n0_8255_8409 n2_8255_8409 0.0
V19380 n0_8255_10569 n2_8255_10569 0.0
V19381 n0_8255_10602 n2_8255_10602 0.0
V19382 n0_8255_14025 n2_8255_14025 0.0
V19383 n0_8255_15105 n2_8255_15105 0.0
V19384 n0_8255_15138 n2_8255_15138 0.0
V19385 n0_8255_16185 n2_8255_16185 0.0
V19386 n0_8255_16218 n2_8255_16218 0.0
V19387 n0_8255_17298 n2_8255_17298 0.0
V19388 n0_8255_17312 n2_8255_17312 0.0
V19389 n0_8255_18392 n2_8255_18392 0.0
V19390 n0_8255_18421 n2_8255_18421 0.0
V19391 n0_8255_19641 n2_8255_19641 0.0
V19392 n0_8255_19674 n2_8255_19674 0.0
V19393 n0_8255_20721 n2_8255_20721 0.0
V19394 n0_8255_20754 n2_8255_20754 0.0
V19395 n0_8304_201 n2_8304_201 0.0
V19396 n0_8304_234 n2_8304_234 0.0
V19397 n0_8304_417 n2_8304_417 0.0
V19398 n0_8304_450 n2_8304_450 0.0
V19399 n0_8304_633 n2_8304_633 0.0
V19400 n0_8304_666 n2_8304_666 0.0
V19401 n0_8304_849 n2_8304_849 0.0
V19402 n0_8304_882 n2_8304_882 0.0
V19403 n0_8304_1065 n2_8304_1065 0.0
V19404 n0_8304_1098 n2_8304_1098 0.0
V19405 n0_8304_1281 n2_8304_1281 0.0
V19406 n0_8304_1314 n2_8304_1314 0.0
V19407 n0_8304_1497 n2_8304_1497 0.0
V19408 n0_8304_1530 n2_8304_1530 0.0
V19409 n0_8304_1713 n2_8304_1713 0.0
V19410 n0_8304_1746 n2_8304_1746 0.0
V19411 n0_8304_1760 n2_8304_1760 0.0
V19412 n0_8304_1783 n2_8304_1783 0.0
V19413 n0_8304_1929 n2_8304_1929 0.0
V19414 n0_8304_1962 n2_8304_1962 0.0
V19415 n0_8304_2145 n2_8304_2145 0.0
V19416 n0_8304_2178 n2_8304_2178 0.0
V19417 n0_8304_2361 n2_8304_2361 0.0
V19418 n0_8304_2394 n2_8304_2394 0.0
V19419 n0_8304_2408 n2_8304_2408 0.0
V19420 n0_8304_2577 n2_8304_2577 0.0
V19421 n0_8304_2610 n2_8304_2610 0.0
V19422 n0_8304_2793 n2_8304_2793 0.0
V19423 n0_8304_2826 n2_8304_2826 0.0
V19424 n0_8304_2840 n2_8304_2840 0.0
V19425 n0_8304_2863 n2_8304_2863 0.0
V19426 n0_8304_3009 n2_8304_3009 0.0
V19427 n0_8304_3042 n2_8304_3042 0.0
V19428 n0_8304_3225 n2_8304_3225 0.0
V19429 n0_8304_3258 n2_8304_3258 0.0
V19430 n0_8304_3441 n2_8304_3441 0.0
V19431 n0_8304_3474 n2_8304_3474 0.0
V19432 n0_8304_3488 n2_8304_3488 0.0
V19433 n0_8304_3657 n2_8304_3657 0.0
V19434 n0_8304_3690 n2_8304_3690 0.0
V19435 n0_8304_3873 n2_8304_3873 0.0
V19436 n0_8304_3906 n2_8304_3906 0.0
V19437 n0_8304_4089 n2_8304_4089 0.0
V19438 n0_8304_4122 n2_8304_4122 0.0
V19439 n0_8304_4136 n2_8304_4136 0.0
V19440 n0_8304_4305 n2_8304_4305 0.0
V19441 n0_8304_4338 n2_8304_4338 0.0
V19442 n0_8304_4521 n2_8304_4521 0.0
V19443 n0_8304_4554 n2_8304_4554 0.0
V19444 n0_8304_4568 n2_8304_4568 0.0
V19445 n0_8304_4737 n2_8304_4737 0.0
V19446 n0_8304_4770 n2_8304_4770 0.0
V19447 n0_8304_4953 n2_8304_4953 0.0
V19448 n0_8304_4986 n2_8304_4986 0.0
V19449 n0_8304_5169 n2_8304_5169 0.0
V19450 n0_8304_5202 n2_8304_5202 0.0
V19451 n0_8304_5216 n2_8304_5216 0.0
V19452 n0_8304_5239 n2_8304_5239 0.0
V19453 n0_8304_5385 n2_8304_5385 0.0
V19454 n0_8304_5418 n2_8304_5418 0.0
V19455 n0_8304_5432 n2_8304_5432 0.0
V19456 n0_8304_5455 n2_8304_5455 0.0
V19457 n0_8304_5601 n2_8304_5601 0.0
V19458 n0_8304_5634 n2_8304_5634 0.0
V19459 n0_8304_5817 n2_8304_5817 0.0
V19460 n0_8304_5850 n2_8304_5850 0.0
V19461 n0_8304_6033 n2_8304_6033 0.0
V19462 n0_8304_6066 n2_8304_6066 0.0
V19463 n0_8304_6249 n2_8304_6249 0.0
V19464 n0_8304_6282 n2_8304_6282 0.0
V19465 n0_8304_6465 n2_8304_6465 0.0
V19466 n0_8304_6498 n2_8304_6498 0.0
V19467 n0_8304_6512 n2_8304_6512 0.0
V19468 n0_8304_6535 n2_8304_6535 0.0
V19469 n0_8304_6681 n2_8304_6681 0.0
V19470 n0_8304_6714 n2_8304_6714 0.0
V19471 n0_8304_6897 n2_8304_6897 0.0
V19472 n0_8304_6930 n2_8304_6930 0.0
V19473 n0_8304_6944 n2_8304_6944 0.0
V19474 n0_8304_7113 n2_8304_7113 0.0
V19475 n0_8304_7146 n2_8304_7146 0.0
V19476 n0_8304_7160 n2_8304_7160 0.0
V19477 n0_8304_7329 n2_8304_7329 0.0
V19478 n0_8304_7362 n2_8304_7362 0.0
V19479 n0_8304_7376 n2_8304_7376 0.0
V19480 n0_8304_7545 n2_8304_7545 0.0
V19481 n0_8304_7578 n2_8304_7578 0.0
V19482 n0_8304_7761 n2_8304_7761 0.0
V19483 n0_8304_7794 n2_8304_7794 0.0
V19484 n0_8304_7808 n2_8304_7808 0.0
V19485 n0_8304_7977 n2_8304_7977 0.0
V19486 n0_8304_8010 n2_8304_8010 0.0
V19487 n0_8304_8193 n2_8304_8193 0.0
V19488 n0_8304_8226 n2_8304_8226 0.0
V19489 n0_8304_8409 n2_8304_8409 0.0
V19490 n0_8304_8442 n2_8304_8442 0.0
V19491 n0_8304_8625 n2_8304_8625 0.0
V19492 n0_8304_8658 n2_8304_8658 0.0
V19493 n0_8304_8841 n2_8304_8841 0.0
V19494 n0_8304_8874 n2_8304_8874 0.0
V19495 n0_8304_8888 n2_8304_8888 0.0
V19496 n0_8304_8909 n2_8304_8909 0.0
V19497 n0_8304_9057 n2_8304_9057 0.0
V19498 n0_8304_9090 n2_8304_9090 0.0
V19499 n0_8304_9273 n2_8304_9273 0.0
V19500 n0_8304_9306 n2_8304_9306 0.0
V19501 n0_8304_9705 n2_8304_9705 0.0
V19502 n0_8304_9738 n2_8304_9738 0.0
V19503 n0_8304_9921 n2_8304_9921 0.0
V19504 n0_8304_9954 n2_8304_9954 0.0
V19505 n0_8304_9968 n2_8304_9968 0.0
V19506 n0_8304_10034 n2_8304_10034 0.0
V19507 n0_8304_10137 n2_8304_10137 0.0
V19508 n0_8304_10170 n2_8304_10170 0.0
V19509 n0_8304_10353 n2_8304_10353 0.0
V19510 n0_8304_10386 n2_8304_10386 0.0
V19511 n0_8304_10569 n2_8304_10569 0.0
V19512 n0_8304_10602 n2_8304_10602 0.0
V19513 n0_8304_10785 n2_8304_10785 0.0
V19514 n0_8304_10818 n2_8304_10818 0.0
V19515 n0_8304_11001 n2_8304_11001 0.0
V19516 n0_8304_11034 n2_8304_11034 0.0
V19517 n0_8304_11048 n2_8304_11048 0.0
V19518 n0_8304_11160 n2_8304_11160 0.0
V19519 n0_8304_11217 n2_8304_11217 0.0
V19520 n0_8304_11250 n2_8304_11250 0.0
V19521 n0_8304_11433 n2_8304_11433 0.0
V19522 n0_8304_11466 n2_8304_11466 0.0
V19523 n0_8304_11865 n2_8304_11865 0.0
V19524 n0_8304_11898 n2_8304_11898 0.0
V19525 n0_8304_12081 n2_8304_12081 0.0
V19526 n0_8304_12114 n2_8304_12114 0.0
V19527 n0_8304_12128 n2_8304_12128 0.0
V19528 n0_8304_12285 n2_8304_12285 0.0
V19529 n0_8304_12297 n2_8304_12297 0.0
V19530 n0_8304_12330 n2_8304_12330 0.0
V19531 n0_8304_12513 n2_8304_12513 0.0
V19532 n0_8304_12546 n2_8304_12546 0.0
V19533 n0_8304_12729 n2_8304_12729 0.0
V19534 n0_8304_12762 n2_8304_12762 0.0
V19535 n0_8304_12945 n2_8304_12945 0.0
V19536 n0_8304_12978 n2_8304_12978 0.0
V19537 n0_8304_13161 n2_8304_13161 0.0
V19538 n0_8304_13194 n2_8304_13194 0.0
V19539 n0_8304_13377 n2_8304_13377 0.0
V19540 n0_8304_13410 n2_8304_13410 0.0
V19541 n0_8304_13424 n2_8304_13424 0.0
V19542 n0_8304_13593 n2_8304_13593 0.0
V19543 n0_8304_13626 n2_8304_13626 0.0
V19544 n0_8304_13640 n2_8304_13640 0.0
V19545 n0_8304_13809 n2_8304_13809 0.0
V19546 n0_8304_13842 n2_8304_13842 0.0
V19547 n0_8304_13856 n2_8304_13856 0.0
V19548 n0_8304_14025 n2_8304_14025 0.0
V19549 n0_8304_14058 n2_8304_14058 0.0
V19550 n0_8304_14072 n2_8304_14072 0.0
V19551 n0_8304_14241 n2_8304_14241 0.0
V19552 n0_8304_14274 n2_8304_14274 0.0
V19553 n0_8304_14396 n2_8304_14396 0.0
V19554 n0_8304_14457 n2_8304_14457 0.0
V19555 n0_8304_14490 n2_8304_14490 0.0
V19556 n0_8304_14504 n2_8304_14504 0.0
V19557 n0_8304_14673 n2_8304_14673 0.0
V19558 n0_8304_14706 n2_8304_14706 0.0
V19559 n0_8304_14889 n2_8304_14889 0.0
V19560 n0_8304_14922 n2_8304_14922 0.0
V19561 n0_8304_15105 n2_8304_15105 0.0
V19562 n0_8304_15138 n2_8304_15138 0.0
V19563 n0_8304_15321 n2_8304_15321 0.0
V19564 n0_8304_15354 n2_8304_15354 0.0
V19565 n0_8304_15537 n2_8304_15537 0.0
V19566 n0_8304_15570 n2_8304_15570 0.0
V19567 n0_8304_15584 n2_8304_15584 0.0
V19568 n0_8304_15753 n2_8304_15753 0.0
V19569 n0_8304_15786 n2_8304_15786 0.0
V19570 n0_8304_15800 n2_8304_15800 0.0
V19571 n0_8304_15969 n2_8304_15969 0.0
V19572 n0_8304_16002 n2_8304_16002 0.0
V19573 n0_8304_16016 n2_8304_16016 0.0
V19574 n0_8304_16185 n2_8304_16185 0.0
V19575 n0_8304_16218 n2_8304_16218 0.0
V19576 n0_8304_16401 n2_8304_16401 0.0
V19577 n0_8304_16434 n2_8304_16434 0.0
V19578 n0_8304_16617 n2_8304_16617 0.0
V19579 n0_8304_16650 n2_8304_16650 0.0
V19580 n0_8304_16833 n2_8304_16833 0.0
V19581 n0_8304_16866 n2_8304_16866 0.0
V19582 n0_8304_17049 n2_8304_17049 0.0
V19583 n0_8304_17082 n2_8304_17082 0.0
V19584 n0_8304_17096 n2_8304_17096 0.0
V19585 n0_8304_17119 n2_8304_17119 0.0
V19586 n0_8304_17265 n2_8304_17265 0.0
V19587 n0_8304_17298 n2_8304_17298 0.0
V19588 n0_8304_17312 n2_8304_17312 0.0
V19589 n0_8304_17481 n2_8304_17481 0.0
V19590 n0_8304_17514 n2_8304_17514 0.0
V19591 n0_8304_17697 n2_8304_17697 0.0
V19592 n0_8304_17730 n2_8304_17730 0.0
V19593 n0_8304_17913 n2_8304_17913 0.0
V19594 n0_8304_17946 n2_8304_17946 0.0
V19595 n0_8304_18129 n2_8304_18129 0.0
V19596 n0_8304_18162 n2_8304_18162 0.0
V19597 n0_8304_18345 n2_8304_18345 0.0
V19598 n0_8304_18378 n2_8304_18378 0.0
V19599 n0_8304_18392 n2_8304_18392 0.0
V19600 n0_8304_18421 n2_8304_18421 0.0
V19601 n0_8304_18561 n2_8304_18561 0.0
V19602 n0_8304_18594 n2_8304_18594 0.0
V19603 n0_8304_18608 n2_8304_18608 0.0
V19604 n0_8304_18777 n2_8304_18777 0.0
V19605 n0_8304_18810 n2_8304_18810 0.0
V19606 n0_8304_18993 n2_8304_18993 0.0
V19607 n0_8304_19026 n2_8304_19026 0.0
V19608 n0_8304_19209 n2_8304_19209 0.0
V19609 n0_8304_19242 n2_8304_19242 0.0
V19610 n0_8304_19256 n2_8304_19256 0.0
V19611 n0_8304_19279 n2_8304_19279 0.0
V19612 n0_8304_19425 n2_8304_19425 0.0
V19613 n0_8304_19458 n2_8304_19458 0.0
V19614 n0_8304_19641 n2_8304_19641 0.0
V19615 n0_8304_19674 n2_8304_19674 0.0
V19616 n0_8304_19857 n2_8304_19857 0.0
V19617 n0_8304_19890 n2_8304_19890 0.0
V19618 n0_8304_20073 n2_8304_20073 0.0
V19619 n0_8304_20106 n2_8304_20106 0.0
V19620 n0_8304_20289 n2_8304_20289 0.0
V19621 n0_8304_20322 n2_8304_20322 0.0
V19622 n0_8304_20505 n2_8304_20505 0.0
V19623 n0_8304_20538 n2_8304_20538 0.0
V19624 n0_8304_20721 n2_8304_20721 0.0
V19625 n0_8304_20754 n2_8304_20754 0.0
V19626 n0_8304_20937 n2_8304_20937 0.0
V19627 n0_8304_20970 n2_8304_20970 0.0
V19628 n0_8396_201 n2_8396_201 0.0
V19629 n0_8396_234 n2_8396_234 0.0
V19630 n0_8396_417 n2_8396_417 0.0
V19631 n0_8396_450 n2_8396_450 0.0
V19632 n0_8396_633 n2_8396_633 0.0
V19633 n0_8396_666 n2_8396_666 0.0
V19634 n0_8396_849 n2_8396_849 0.0
V19635 n0_8396_882 n2_8396_882 0.0
V19636 n0_8396_1065 n2_8396_1065 0.0
V19637 n0_8396_1098 n2_8396_1098 0.0
V19638 n0_8396_1281 n2_8396_1281 0.0
V19639 n0_8396_1314 n2_8396_1314 0.0
V19640 n0_8396_1497 n2_8396_1497 0.0
V19641 n0_8396_1530 n2_8396_1530 0.0
V19642 n0_8396_1713 n2_8396_1713 0.0
V19643 n0_8396_1746 n2_8396_1746 0.0
V19644 n0_8396_1760 n2_8396_1760 0.0
V19645 n0_8396_1783 n2_8396_1783 0.0
V19646 n0_8396_1929 n2_8396_1929 0.0
V19647 n0_8396_1962 n2_8396_1962 0.0
V19648 n0_8396_2145 n2_8396_2145 0.0
V19649 n0_8396_2178 n2_8396_2178 0.0
V19650 n0_8396_2361 n2_8396_2361 0.0
V19651 n0_8396_2394 n2_8396_2394 0.0
V19652 n0_8396_2408 n2_8396_2408 0.0
V19653 n0_8396_2577 n2_8396_2577 0.0
V19654 n0_8396_2610 n2_8396_2610 0.0
V19655 n0_8396_2793 n2_8396_2793 0.0
V19656 n0_8396_2826 n2_8396_2826 0.0
V19657 n0_8396_2840 n2_8396_2840 0.0
V19658 n0_8396_2863 n2_8396_2863 0.0
V19659 n0_8396_3009 n2_8396_3009 0.0
V19660 n0_8396_3042 n2_8396_3042 0.0
V19661 n0_8396_3225 n2_8396_3225 0.0
V19662 n0_8396_3258 n2_8396_3258 0.0
V19663 n0_8396_3441 n2_8396_3441 0.0
V19664 n0_8396_3474 n2_8396_3474 0.0
V19665 n0_8396_3488 n2_8396_3488 0.0
V19666 n0_8396_3657 n2_8396_3657 0.0
V19667 n0_8396_3690 n2_8396_3690 0.0
V19668 n0_8396_3873 n2_8396_3873 0.0
V19669 n0_8396_3906 n2_8396_3906 0.0
V19670 n0_8396_4089 n2_8396_4089 0.0
V19671 n0_8396_4122 n2_8396_4122 0.0
V19672 n0_8396_4136 n2_8396_4136 0.0
V19673 n0_8396_4305 n2_8396_4305 0.0
V19674 n0_8396_4338 n2_8396_4338 0.0
V19675 n0_8396_4521 n2_8396_4521 0.0
V19676 n0_8396_4554 n2_8396_4554 0.0
V19677 n0_8396_4568 n2_8396_4568 0.0
V19678 n0_8396_4737 n2_8396_4737 0.0
V19679 n0_8396_4770 n2_8396_4770 0.0
V19680 n0_8396_4953 n2_8396_4953 0.0
V19681 n0_8396_5169 n2_8396_5169 0.0
V19682 n0_8396_5202 n2_8396_5202 0.0
V19683 n0_8396_5216 n2_8396_5216 0.0
V19684 n0_8396_5239 n2_8396_5239 0.0
V19685 n0_8396_5385 n2_8396_5385 0.0
V19686 n0_8396_5418 n2_8396_5418 0.0
V19687 n0_8396_5432 n2_8396_5432 0.0
V19688 n0_8396_5455 n2_8396_5455 0.0
V19689 n0_8396_5601 n2_8396_5601 0.0
V19690 n0_8396_5634 n2_8396_5634 0.0
V19691 n0_8396_5817 n2_8396_5817 0.0
V19692 n0_8396_5850 n2_8396_5850 0.0
V19693 n0_8396_6033 n2_8396_6033 0.0
V19694 n0_8396_6066 n2_8396_6066 0.0
V19695 n0_8396_6249 n2_8396_6249 0.0
V19696 n0_8396_6282 n2_8396_6282 0.0
V19697 n0_8396_6465 n2_8396_6465 0.0
V19698 n0_8396_6498 n2_8396_6498 0.0
V19699 n0_8396_6512 n2_8396_6512 0.0
V19700 n0_8396_6535 n2_8396_6535 0.0
V19701 n0_8396_6681 n2_8396_6681 0.0
V19702 n0_8396_6714 n2_8396_6714 0.0
V19703 n0_8396_6897 n2_8396_6897 0.0
V19704 n0_8396_6930 n2_8396_6930 0.0
V19705 n0_8396_6944 n2_8396_6944 0.0
V19706 n0_8396_7113 n2_8396_7113 0.0
V19707 n0_8396_7146 n2_8396_7146 0.0
V19708 n0_8396_7160 n2_8396_7160 0.0
V19709 n0_8396_7329 n2_8396_7329 0.0
V19710 n0_8396_7362 n2_8396_7362 0.0
V19711 n0_8396_7376 n2_8396_7376 0.0
V19712 n0_8396_7545 n2_8396_7545 0.0
V19713 n0_8396_7578 n2_8396_7578 0.0
V19714 n0_8396_7761 n2_8396_7761 0.0
V19715 n0_8396_7794 n2_8396_7794 0.0
V19716 n0_8396_7808 n2_8396_7808 0.0
V19717 n0_8396_7977 n2_8396_7977 0.0
V19718 n0_8396_8010 n2_8396_8010 0.0
V19719 n0_8396_8193 n2_8396_8193 0.0
V19720 n0_8396_8226 n2_8396_8226 0.0
V19721 n0_8396_12945 n2_8396_12945 0.0
V19722 n0_8396_12978 n2_8396_12978 0.0
V19723 n0_8396_13161 n2_8396_13161 0.0
V19724 n0_8396_13194 n2_8396_13194 0.0
V19725 n0_8396_13377 n2_8396_13377 0.0
V19726 n0_8396_13410 n2_8396_13410 0.0
V19727 n0_8396_13424 n2_8396_13424 0.0
V19728 n0_8396_13593 n2_8396_13593 0.0
V19729 n0_8396_13626 n2_8396_13626 0.0
V19730 n0_8396_13640 n2_8396_13640 0.0
V19731 n0_8396_13809 n2_8396_13809 0.0
V19732 n0_8396_13842 n2_8396_13842 0.0
V19733 n0_8396_13856 n2_8396_13856 0.0
V19734 n0_8396_14025 n2_8396_14025 0.0
V19735 n0_8396_14058 n2_8396_14058 0.0
V19736 n0_8396_14072 n2_8396_14072 0.0
V19737 n0_8396_14241 n2_8396_14241 0.0
V19738 n0_8396_14274 n2_8396_14274 0.0
V19739 n0_8396_14396 n2_8396_14396 0.0
V19740 n0_8396_14457 n2_8396_14457 0.0
V19741 n0_8396_14490 n2_8396_14490 0.0
V19742 n0_8396_14504 n2_8396_14504 0.0
V19743 n0_8396_14673 n2_8396_14673 0.0
V19744 n0_8396_14706 n2_8396_14706 0.0
V19745 n0_8396_14889 n2_8396_14889 0.0
V19746 n0_8396_14922 n2_8396_14922 0.0
V19747 n0_8396_15138 n2_8396_15138 0.0
V19748 n0_8396_15321 n2_8396_15321 0.0
V19749 n0_8396_15354 n2_8396_15354 0.0
V19750 n0_8396_15537 n2_8396_15537 0.0
V19751 n0_8396_15570 n2_8396_15570 0.0
V19752 n0_8396_15584 n2_8396_15584 0.0
V19753 n0_8396_15753 n2_8396_15753 0.0
V19754 n0_8396_15786 n2_8396_15786 0.0
V19755 n0_8396_15800 n2_8396_15800 0.0
V19756 n0_8396_15969 n2_8396_15969 0.0
V19757 n0_8396_16002 n2_8396_16002 0.0
V19758 n0_8396_16016 n2_8396_16016 0.0
V19759 n0_8396_16185 n2_8396_16185 0.0
V19760 n0_8396_16401 n2_8396_16401 0.0
V19761 n0_8396_16434 n2_8396_16434 0.0
V19762 n0_8396_16617 n2_8396_16617 0.0
V19763 n0_8396_16650 n2_8396_16650 0.0
V19764 n0_8396_16833 n2_8396_16833 0.0
V19765 n0_8396_16866 n2_8396_16866 0.0
V19766 n0_8396_17049 n2_8396_17049 0.0
V19767 n0_8396_17082 n2_8396_17082 0.0
V19768 n0_8396_17096 n2_8396_17096 0.0
V19769 n0_8396_17119 n2_8396_17119 0.0
V19770 n0_8396_17265 n2_8396_17265 0.0
V19771 n0_8396_17298 n2_8396_17298 0.0
V19772 n0_8396_17312 n2_8396_17312 0.0
V19773 n0_8396_17481 n2_8396_17481 0.0
V19774 n0_8396_17514 n2_8396_17514 0.0
V19775 n0_8396_17697 n2_8396_17697 0.0
V19776 n0_8396_17730 n2_8396_17730 0.0
V19777 n0_8396_17913 n2_8396_17913 0.0
V19778 n0_8396_17946 n2_8396_17946 0.0
V19779 n0_8396_18129 n2_8396_18129 0.0
V19780 n0_8396_18162 n2_8396_18162 0.0
V19781 n0_8396_18345 n2_8396_18345 0.0
V19782 n0_8396_18378 n2_8396_18378 0.0
V19783 n0_8396_18392 n2_8396_18392 0.0
V19784 n0_8396_18421 n2_8396_18421 0.0
V19785 n0_8396_18561 n2_8396_18561 0.0
V19786 n0_8396_18594 n2_8396_18594 0.0
V19787 n0_8396_18608 n2_8396_18608 0.0
V19788 n0_8396_18777 n2_8396_18777 0.0
V19789 n0_8396_18810 n2_8396_18810 0.0
V19790 n0_8396_18993 n2_8396_18993 0.0
V19791 n0_8396_19026 n2_8396_19026 0.0
V19792 n0_8396_19209 n2_8396_19209 0.0
V19793 n0_8396_19242 n2_8396_19242 0.0
V19794 n0_8396_19256 n2_8396_19256 0.0
V19795 n0_8396_19279 n2_8396_19279 0.0
V19796 n0_8396_19425 n2_8396_19425 0.0
V19797 n0_8396_19458 n2_8396_19458 0.0
V19798 n0_8396_19641 n2_8396_19641 0.0
V19799 n0_8396_19674 n2_8396_19674 0.0
V19800 n0_8396_19857 n2_8396_19857 0.0
V19801 n0_8396_19890 n2_8396_19890 0.0
V19802 n0_8396_20073 n2_8396_20073 0.0
V19803 n0_8396_20106 n2_8396_20106 0.0
V19804 n0_8396_20289 n2_8396_20289 0.0
V19805 n0_8396_20322 n2_8396_20322 0.0
V19806 n0_8396_20505 n2_8396_20505 0.0
V19807 n0_8396_20538 n2_8396_20538 0.0
V19808 n0_8396_20754 n2_8396_20754 0.0
V19809 n0_8396_20937 n2_8396_20937 0.0
V19810 n0_8396_20970 n2_8396_20970 0.0
V19811 n0_9241_9489 n2_9241_9489 0.0
V19812 n0_9241_9522 n2_9241_9522 0.0
V19813 n0_9241_9705 n2_9241_9705 0.0
V19814 n0_9241_9738 n2_9241_9738 0.0
V19815 n0_9241_9921 n2_9241_9921 0.0
V19816 n0_9241_9954 n2_9241_9954 0.0
V19817 n0_9241_10034 n2_9241_10034 0.0
V19818 n0_9241_10137 n2_9241_10137 0.0
V19819 n0_9241_10170 n2_9241_10170 0.0
V19820 n0_9241_10353 n2_9241_10353 0.0
V19821 n0_9241_10386 n2_9241_10386 0.0
V19822 n0_9241_10569 n2_9241_10569 0.0
V19823 n0_9241_10785 n2_9241_10785 0.0
V19824 n0_9241_10818 n2_9241_10818 0.0
V19825 n0_9241_11001 n2_9241_11001 0.0
V19826 n0_9241_11034 n2_9241_11034 0.0
V19827 n0_9241_11160 n2_9241_11160 0.0
V19828 n0_9241_11217 n2_9241_11217 0.0
V19829 n0_9241_11250 n2_9241_11250 0.0
V19830 n0_9241_11433 n2_9241_11433 0.0
V19831 n0_9241_11466 n2_9241_11466 0.0
V19832 n0_9241_11649 n2_9241_11649 0.0
V19833 n0_9241_11682 n2_9241_11682 0.0
V19834 n0_9380_10569 n2_9380_10569 0.0
V19835 n0_9380_10602 n2_9380_10602 0.0
V19836 n0_9429_9705 n2_9429_9705 0.0
V19837 n0_9429_9738 n2_9429_9738 0.0
V19838 n0_9429_9921 n2_9429_9921 0.0
V19839 n0_9429_9954 n2_9429_9954 0.0
V19840 n0_9429_10137 n2_9429_10137 0.0
V19841 n0_9429_10170 n2_9429_10170 0.0
V19842 n0_9429_10353 n2_9429_10353 0.0
V19843 n0_9429_10386 n2_9429_10386 0.0
V19844 n0_9429_10569 n2_9429_10569 0.0
V19845 n0_9429_10602 n2_9429_10602 0.0
V19846 n0_9429_10785 n2_9429_10785 0.0
V19847 n0_9429_10818 n2_9429_10818 0.0
V19848 n0_9429_11001 n2_9429_11001 0.0
V19849 n0_9429_11034 n2_9429_11034 0.0
V19850 n0_9429_11217 n2_9429_11217 0.0
V19851 n0_9429_11250 n2_9429_11250 0.0
V19852 n0_9429_11433 n2_9429_11433 0.0
V19853 n0_9429_11466 n2_9429_11466 0.0
V19854 n0_10366_201 n2_10366_201 0.0
V19855 n0_10366_234 n2_10366_234 0.0
V19856 n0_10366_417 n2_10366_417 0.0
V19857 n0_10366_450 n2_10366_450 0.0
V19858 n0_10366_633 n2_10366_633 0.0
V19859 n0_10366_666 n2_10366_666 0.0
V19860 n0_10366_849 n2_10366_849 0.0
V19861 n0_10366_882 n2_10366_882 0.0
V19862 n0_10366_1065 n2_10366_1065 0.0
V19863 n0_10366_1098 n2_10366_1098 0.0
V19864 n0_10366_1281 n2_10366_1281 0.0
V19865 n0_10366_1314 n2_10366_1314 0.0
V19866 n0_10366_1497 n2_10366_1497 0.0
V19867 n0_10366_1530 n2_10366_1530 0.0
V19868 n0_10366_1713 n2_10366_1713 0.0
V19869 n0_10366_1746 n2_10366_1746 0.0
V19870 n0_10366_1760 n2_10366_1760 0.0
V19871 n0_10366_1783 n2_10366_1783 0.0
V19872 n0_10366_1929 n2_10366_1929 0.0
V19873 n0_10366_1962 n2_10366_1962 0.0
V19874 n0_10366_2145 n2_10366_2145 0.0
V19875 n0_10366_2178 n2_10366_2178 0.0
V19876 n0_10366_2361 n2_10366_2361 0.0
V19877 n0_10366_2394 n2_10366_2394 0.0
V19878 n0_10366_2408 n2_10366_2408 0.0
V19879 n0_10366_2577 n2_10366_2577 0.0
V19880 n0_10366_2610 n2_10366_2610 0.0
V19881 n0_10366_2647 n2_10366_2647 0.0
V19882 n0_10366_2793 n2_10366_2793 0.0
V19883 n0_10366_2826 n2_10366_2826 0.0
V19884 n0_10366_2840 n2_10366_2840 0.0
V19885 n0_10366_2863 n2_10366_2863 0.0
V19886 n0_10366_3009 n2_10366_3009 0.0
V19887 n0_10366_3042 n2_10366_3042 0.0
V19888 n0_10366_3225 n2_10366_3225 0.0
V19889 n0_10366_3258 n2_10366_3258 0.0
V19890 n0_10366_3441 n2_10366_3441 0.0
V19891 n0_10366_3474 n2_10366_3474 0.0
V19892 n0_10366_3488 n2_10366_3488 0.0
V19893 n0_10366_3511 n2_10366_3511 0.0
V19894 n0_10366_3657 n2_10366_3657 0.0
V19895 n0_10366_3690 n2_10366_3690 0.0
V19896 n0_10366_3873 n2_10366_3873 0.0
V19897 n0_10366_3906 n2_10366_3906 0.0
V19898 n0_10366_4089 n2_10366_4089 0.0
V19899 n0_10366_4122 n2_10366_4122 0.0
V19900 n0_10366_4136 n2_10366_4136 0.0
V19901 n0_10366_4159 n2_10366_4159 0.0
V19902 n0_10366_4305 n2_10366_4305 0.0
V19903 n0_10366_4338 n2_10366_4338 0.0
V19904 n0_10366_4521 n2_10366_4521 0.0
V19905 n0_10366_4554 n2_10366_4554 0.0
V19906 n0_10366_4568 n2_10366_4568 0.0
V19907 n0_10366_4591 n2_10366_4591 0.0
V19908 n0_10366_4737 n2_10366_4737 0.0
V19909 n0_10366_4770 n2_10366_4770 0.0
V19910 n0_10366_4953 n2_10366_4953 0.0
V19911 n0_10366_5169 n2_10366_5169 0.0
V19912 n0_10366_5202 n2_10366_5202 0.0
V19913 n0_10366_5239 n2_10366_5239 0.0
V19914 n0_10366_5385 n2_10366_5385 0.0
V19915 n0_10366_5418 n2_10366_5418 0.0
V19916 n0_10366_5432 n2_10366_5432 0.0
V19917 n0_10366_5455 n2_10366_5455 0.0
V19918 n0_10366_5601 n2_10366_5601 0.0
V19919 n0_10366_5634 n2_10366_5634 0.0
V19920 n0_10366_5817 n2_10366_5817 0.0
V19921 n0_10366_5850 n2_10366_5850 0.0
V19922 n0_10366_6033 n2_10366_6033 0.0
V19923 n0_10366_6066 n2_10366_6066 0.0
V19924 n0_10366_6249 n2_10366_6249 0.0
V19925 n0_10366_6282 n2_10366_6282 0.0
V19926 n0_10366_6465 n2_10366_6465 0.0
V19927 n0_10366_6498 n2_10366_6498 0.0
V19928 n0_10366_6512 n2_10366_6512 0.0
V19929 n0_10366_6535 n2_10366_6535 0.0
V19930 n0_10366_6681 n2_10366_6681 0.0
V19931 n0_10366_6714 n2_10366_6714 0.0
V19932 n0_10366_6751 n2_10366_6751 0.0
V19933 n0_10366_6897 n2_10366_6897 0.0
V19934 n0_10366_6930 n2_10366_6930 0.0
V19935 n0_10366_6944 n2_10366_6944 0.0
V19936 n0_10366_6967 n2_10366_6967 0.0
V19937 n0_10366_7113 n2_10366_7113 0.0
V19938 n0_10366_7146 n2_10366_7146 0.0
V19939 n0_10366_7160 n2_10366_7160 0.0
V19940 n0_10366_7178 n2_10366_7178 0.0
V19941 n0_10366_7329 n2_10366_7329 0.0
V19942 n0_10366_7362 n2_10366_7362 0.0
V19943 n0_10366_7376 n2_10366_7376 0.0
V19944 n0_10366_7399 n2_10366_7399 0.0
V19945 n0_10366_7545 n2_10366_7545 0.0
V19946 n0_10366_7578 n2_10366_7578 0.0
V19947 n0_10366_7761 n2_10366_7761 0.0
V19948 n0_10366_7794 n2_10366_7794 0.0
V19949 n0_10366_7977 n2_10366_7977 0.0
V19950 n0_10366_8010 n2_10366_8010 0.0
V19951 n0_10366_8193 n2_10366_8193 0.0
V19952 n0_10366_8226 n2_10366_8226 0.0
V19953 n0_10366_8409 n2_10366_8409 0.0
V19954 n0_10366_8442 n2_10366_8442 0.0
V19955 n0_10366_8613 n2_10366_8613 0.0
V19956 n0_10366_8625 n2_10366_8625 0.0
V19957 n0_10366_8658 n2_10366_8658 0.0
V19958 n0_10366_8841 n2_10366_8841 0.0
V19959 n0_10366_8874 n2_10366_8874 0.0
V19960 n0_10366_9057 n2_10366_9057 0.0
V19961 n0_10366_9090 n2_10366_9090 0.0
V19962 n0_10366_9190 n2_10366_9190 0.0
V19963 n0_10366_9273 n2_10366_9273 0.0
V19964 n0_10366_9306 n2_10366_9306 0.0
V19965 n0_10366_9489 n2_10366_9489 0.0
V19966 n0_10366_9522 n2_10366_9522 0.0
V19967 n0_10366_9705 n2_10366_9705 0.0
V19968 n0_10366_9738 n2_10366_9738 0.0
V19969 n0_10366_9921 n2_10366_9921 0.0
V19970 n0_10366_9954 n2_10366_9954 0.0
V19971 n0_10366_10137 n2_10366_10137 0.0
V19972 n0_10366_10170 n2_10366_10170 0.0
V19973 n0_10366_10353 n2_10366_10353 0.0
V19974 n0_10366_10386 n2_10366_10386 0.0
V19975 n0_10366_10557 n2_10366_10557 0.0
V19976 n0_10366_10569 n2_10366_10569 0.0
V19977 n0_10366_10785 n2_10366_10785 0.0
V19978 n0_10366_10818 n2_10366_10818 0.0
V19979 n0_10366_11001 n2_10366_11001 0.0
V19980 n0_10366_11034 n2_10366_11034 0.0
V19981 n0_10366_11217 n2_10366_11217 0.0
V19982 n0_10366_11250 n2_10366_11250 0.0
V19983 n0_10366_11433 n2_10366_11433 0.0
V19984 n0_10366_11466 n2_10366_11466 0.0
V19985 n0_10366_11649 n2_10366_11649 0.0
V19986 n0_10366_11682 n2_10366_11682 0.0
V19987 n0_10366_11865 n2_10366_11865 0.0
V19988 n0_10366_11898 n2_10366_11898 0.0
V19989 n0_10366_12004 n2_10366_12004 0.0
V19990 n0_10366_12081 n2_10366_12081 0.0
V19991 n0_10366_12114 n2_10366_12114 0.0
V19992 n0_10366_12297 n2_10366_12297 0.0
V19993 n0_10366_12330 n2_10366_12330 0.0
V19994 n0_10366_12513 n2_10366_12513 0.0
V19995 n0_10366_12546 n2_10366_12546 0.0
V19996 n0_10366_12566 n2_10366_12566 0.0
V19997 n0_10366_12729 n2_10366_12729 0.0
V19998 n0_10366_12762 n2_10366_12762 0.0
V19999 n0_10366_12945 n2_10366_12945 0.0
V20000 n0_10366_12978 n2_10366_12978 0.0
V20001 n0_10366_13161 n2_10366_13161 0.0
V20002 n0_10366_13194 n2_10366_13194 0.0
V20003 n0_10366_13377 n2_10366_13377 0.0
V20004 n0_10366_13410 n2_10366_13410 0.0
V20005 n0_10366_13593 n2_10366_13593 0.0
V20006 n0_10366_13626 n2_10366_13626 0.0
V20007 n0_10366_13640 n2_10366_13640 0.0
V20008 n0_10366_13663 n2_10366_13663 0.0
V20009 n0_10366_13809 n2_10366_13809 0.0
V20010 n0_10366_13842 n2_10366_13842 0.0
V20011 n0_10366_13856 n2_10366_13856 0.0
V20012 n0_10366_13879 n2_10366_13879 0.0
V20013 n0_10366_14025 n2_10366_14025 0.0
V20014 n0_10366_14058 n2_10366_14058 0.0
V20015 n0_10366_14072 n2_10366_14072 0.0
V20016 n0_10366_14079 n2_10366_14079 0.0
V20017 n0_10366_14241 n2_10366_14241 0.0
V20018 n0_10366_14274 n2_10366_14274 0.0
V20019 n0_10366_14457 n2_10366_14457 0.0
V20020 n0_10366_14490 n2_10366_14490 0.0
V20021 n0_10366_14504 n2_10366_14504 0.0
V20022 n0_10366_14673 n2_10366_14673 0.0
V20023 n0_10366_14706 n2_10366_14706 0.0
V20024 n0_10366_14889 n2_10366_14889 0.0
V20025 n0_10366_14922 n2_10366_14922 0.0
V20026 n0_10366_15138 n2_10366_15138 0.0
V20027 n0_10366_15321 n2_10366_15321 0.0
V20028 n0_10366_15354 n2_10366_15354 0.0
V20029 n0_10366_15537 n2_10366_15537 0.0
V20030 n0_10366_15570 n2_10366_15570 0.0
V20031 n0_10366_15584 n2_10366_15584 0.0
V20032 n0_10366_15753 n2_10366_15753 0.0
V20033 n0_10366_15786 n2_10366_15786 0.0
V20034 n0_10366_15800 n2_10366_15800 0.0
V20035 n0_10366_15823 n2_10366_15823 0.0
V20036 n0_10366_15969 n2_10366_15969 0.0
V20037 n0_10366_16002 n2_10366_16002 0.0
V20038 n0_10366_16016 n2_10366_16016 0.0
V20039 n0_10366_16185 n2_10366_16185 0.0
V20040 n0_10366_16401 n2_10366_16401 0.0
V20041 n0_10366_16434 n2_10366_16434 0.0
V20042 n0_10366_16617 n2_10366_16617 0.0
V20043 n0_10366_16650 n2_10366_16650 0.0
V20044 n0_10366_16833 n2_10366_16833 0.0
V20045 n0_10366_16866 n2_10366_16866 0.0
V20046 n0_10366_17049 n2_10366_17049 0.0
V20047 n0_10366_17082 n2_10366_17082 0.0
V20048 n0_10366_17096 n2_10366_17096 0.0
V20049 n0_10366_17103 n2_10366_17103 0.0
V20050 n0_10366_17119 n2_10366_17119 0.0
V20051 n0_10366_17265 n2_10366_17265 0.0
V20052 n0_10366_17298 n2_10366_17298 0.0
V20053 n0_10366_17312 n2_10366_17312 0.0
V20054 n0_10366_17481 n2_10366_17481 0.0
V20055 n0_10366_17514 n2_10366_17514 0.0
V20056 n0_10366_17697 n2_10366_17697 0.0
V20057 n0_10366_17730 n2_10366_17730 0.0
V20058 n0_10366_17913 n2_10366_17913 0.0
V20059 n0_10366_17946 n2_10366_17946 0.0
V20060 n0_10366_18129 n2_10366_18129 0.0
V20061 n0_10366_18162 n2_10366_18162 0.0
V20062 n0_10366_18345 n2_10366_18345 0.0
V20063 n0_10366_18378 n2_10366_18378 0.0
V20064 n0_10366_18392 n2_10366_18392 0.0
V20065 n0_10366_18561 n2_10366_18561 0.0
V20066 n0_10366_18594 n2_10366_18594 0.0
V20067 n0_10366_18608 n2_10366_18608 0.0
V20068 n0_10366_18777 n2_10366_18777 0.0
V20069 n0_10366_18810 n2_10366_18810 0.0
V20070 n0_10366_18993 n2_10366_18993 0.0
V20071 n0_10366_19026 n2_10366_19026 0.0
V20072 n0_10366_19209 n2_10366_19209 0.0
V20073 n0_10366_19242 n2_10366_19242 0.0
V20074 n0_10366_19256 n2_10366_19256 0.0
V20075 n0_10366_19425 n2_10366_19425 0.0
V20076 n0_10366_19458 n2_10366_19458 0.0
V20077 n0_10366_19641 n2_10366_19641 0.0
V20078 n0_10366_19674 n2_10366_19674 0.0
V20079 n0_10366_19857 n2_10366_19857 0.0
V20080 n0_10366_19890 n2_10366_19890 0.0
V20081 n0_10366_20073 n2_10366_20073 0.0
V20082 n0_10366_20106 n2_10366_20106 0.0
V20083 n0_10366_20289 n2_10366_20289 0.0
V20084 n0_10366_20322 n2_10366_20322 0.0
V20085 n0_10366_20505 n2_10366_20505 0.0
V20086 n0_10366_20538 n2_10366_20538 0.0
V20087 n0_10366_20754 n2_10366_20754 0.0
V20088 n0_10366_20937 n2_10366_20937 0.0
V20089 n0_10366_20970 n2_10366_20970 0.0
V20090 n0_10458_201 n2_10458_201 0.0
V20091 n0_10458_234 n2_10458_234 0.0
V20092 n0_10458_417 n2_10458_417 0.0
V20093 n0_10458_450 n2_10458_450 0.0
V20094 n0_10458_633 n2_10458_633 0.0
V20095 n0_10458_666 n2_10458_666 0.0
V20096 n0_10458_849 n2_10458_849 0.0
V20097 n0_10458_882 n2_10458_882 0.0
V20098 n0_10458_1065 n2_10458_1065 0.0
V20099 n0_10458_1098 n2_10458_1098 0.0
V20100 n0_10458_1281 n2_10458_1281 0.0
V20101 n0_10458_1314 n2_10458_1314 0.0
V20102 n0_10458_1497 n2_10458_1497 0.0
V20103 n0_10458_1530 n2_10458_1530 0.0
V20104 n0_10458_1713 n2_10458_1713 0.0
V20105 n0_10458_1746 n2_10458_1746 0.0
V20106 n0_10458_1760 n2_10458_1760 0.0
V20107 n0_10458_1783 n2_10458_1783 0.0
V20108 n0_10458_1929 n2_10458_1929 0.0
V20109 n0_10458_1962 n2_10458_1962 0.0
V20110 n0_10458_2145 n2_10458_2145 0.0
V20111 n0_10458_2178 n2_10458_2178 0.0
V20112 n0_10458_2361 n2_10458_2361 0.0
V20113 n0_10458_2394 n2_10458_2394 0.0
V20114 n0_10458_2408 n2_10458_2408 0.0
V20115 n0_10458_2577 n2_10458_2577 0.0
V20116 n0_10458_2610 n2_10458_2610 0.0
V20117 n0_10458_2647 n2_10458_2647 0.0
V20118 n0_10458_2793 n2_10458_2793 0.0
V20119 n0_10458_2826 n2_10458_2826 0.0
V20120 n0_10458_2840 n2_10458_2840 0.0
V20121 n0_10458_2863 n2_10458_2863 0.0
V20122 n0_10458_3009 n2_10458_3009 0.0
V20123 n0_10458_3042 n2_10458_3042 0.0
V20124 n0_10458_3225 n2_10458_3225 0.0
V20125 n0_10458_3258 n2_10458_3258 0.0
V20126 n0_10458_3441 n2_10458_3441 0.0
V20127 n0_10458_3474 n2_10458_3474 0.0
V20128 n0_10458_3488 n2_10458_3488 0.0
V20129 n0_10458_3511 n2_10458_3511 0.0
V20130 n0_10458_3657 n2_10458_3657 0.0
V20131 n0_10458_3690 n2_10458_3690 0.0
V20132 n0_10458_3873 n2_10458_3873 0.0
V20133 n0_10458_3906 n2_10458_3906 0.0
V20134 n0_10458_4089 n2_10458_4089 0.0
V20135 n0_10458_4122 n2_10458_4122 0.0
V20136 n0_10458_4136 n2_10458_4136 0.0
V20137 n0_10458_4159 n2_10458_4159 0.0
V20138 n0_10458_4305 n2_10458_4305 0.0
V20139 n0_10458_4338 n2_10458_4338 0.0
V20140 n0_10458_4521 n2_10458_4521 0.0
V20141 n0_10458_4554 n2_10458_4554 0.0
V20142 n0_10458_4568 n2_10458_4568 0.0
V20143 n0_10458_4591 n2_10458_4591 0.0
V20144 n0_10458_4737 n2_10458_4737 0.0
V20145 n0_10458_4770 n2_10458_4770 0.0
V20146 n0_10458_4953 n2_10458_4953 0.0
V20147 n0_10458_4986 n2_10458_4986 0.0
V20148 n0_10458_5169 n2_10458_5169 0.0
V20149 n0_10458_5202 n2_10458_5202 0.0
V20150 n0_10458_5239 n2_10458_5239 0.0
V20151 n0_10458_5385 n2_10458_5385 0.0
V20152 n0_10458_5418 n2_10458_5418 0.0
V20153 n0_10458_5432 n2_10458_5432 0.0
V20154 n0_10458_5455 n2_10458_5455 0.0
V20155 n0_10458_5601 n2_10458_5601 0.0
V20156 n0_10458_5634 n2_10458_5634 0.0
V20157 n0_10458_5817 n2_10458_5817 0.0
V20158 n0_10458_5850 n2_10458_5850 0.0
V20159 n0_10458_6033 n2_10458_6033 0.0
V20160 n0_10458_6066 n2_10458_6066 0.0
V20161 n0_10458_6249 n2_10458_6249 0.0
V20162 n0_10458_6282 n2_10458_6282 0.0
V20163 n0_10458_6465 n2_10458_6465 0.0
V20164 n0_10458_6498 n2_10458_6498 0.0
V20165 n0_10458_6512 n2_10458_6512 0.0
V20166 n0_10458_6535 n2_10458_6535 0.0
V20167 n0_10458_6681 n2_10458_6681 0.0
V20168 n0_10458_6714 n2_10458_6714 0.0
V20169 n0_10458_6751 n2_10458_6751 0.0
V20170 n0_10458_6897 n2_10458_6897 0.0
V20171 n0_10458_6930 n2_10458_6930 0.0
V20172 n0_10458_6944 n2_10458_6944 0.0
V20173 n0_10458_6967 n2_10458_6967 0.0
V20174 n0_10458_7113 n2_10458_7113 0.0
V20175 n0_10458_7146 n2_10458_7146 0.0
V20176 n0_10458_7160 n2_10458_7160 0.0
V20177 n0_10458_7178 n2_10458_7178 0.0
V20178 n0_10458_7329 n2_10458_7329 0.0
V20179 n0_10458_7362 n2_10458_7362 0.0
V20180 n0_10458_7376 n2_10458_7376 0.0
V20181 n0_10458_7399 n2_10458_7399 0.0
V20182 n0_10458_7545 n2_10458_7545 0.0
V20183 n0_10458_7578 n2_10458_7578 0.0
V20184 n0_10458_7761 n2_10458_7761 0.0
V20185 n0_10458_7794 n2_10458_7794 0.0
V20186 n0_10458_7977 n2_10458_7977 0.0
V20187 n0_10458_8010 n2_10458_8010 0.0
V20188 n0_10458_8193 n2_10458_8193 0.0
V20189 n0_10458_8226 n2_10458_8226 0.0
V20190 n0_10458_8409 n2_10458_8409 0.0
V20191 n0_10458_8442 n2_10458_8442 0.0
V20192 n0_10458_8625 n2_10458_8625 0.0
V20193 n0_10458_8658 n2_10458_8658 0.0
V20194 n0_10458_8841 n2_10458_8841 0.0
V20195 n0_10458_8874 n2_10458_8874 0.0
V20196 n0_10458_9057 n2_10458_9057 0.0
V20197 n0_10458_9090 n2_10458_9090 0.0
V20198 n0_10458_9273 n2_10458_9273 0.0
V20199 n0_10458_9306 n2_10458_9306 0.0
V20200 n0_10458_9489 n2_10458_9489 0.0
V20201 n0_10458_9522 n2_10458_9522 0.0
V20202 n0_10458_9705 n2_10458_9705 0.0
V20203 n0_10458_9738 n2_10458_9738 0.0
V20204 n0_10458_9921 n2_10458_9921 0.0
V20205 n0_10458_9954 n2_10458_9954 0.0
V20206 n0_10458_10137 n2_10458_10137 0.0
V20207 n0_10458_10170 n2_10458_10170 0.0
V20208 n0_10458_10353 n2_10458_10353 0.0
V20209 n0_10458_10386 n2_10458_10386 0.0
V20210 n0_10458_10569 n2_10458_10569 0.0
V20211 n0_10458_10602 n2_10458_10602 0.0
V20212 n0_10458_10785 n2_10458_10785 0.0
V20213 n0_10458_10818 n2_10458_10818 0.0
V20214 n0_10458_11001 n2_10458_11001 0.0
V20215 n0_10458_11034 n2_10458_11034 0.0
V20216 n0_10458_11217 n2_10458_11217 0.0
V20217 n0_10458_11250 n2_10458_11250 0.0
V20218 n0_10458_11433 n2_10458_11433 0.0
V20219 n0_10458_11466 n2_10458_11466 0.0
V20220 n0_10458_11649 n2_10458_11649 0.0
V20221 n0_10458_11682 n2_10458_11682 0.0
V20222 n0_10458_11865 n2_10458_11865 0.0
V20223 n0_10458_11898 n2_10458_11898 0.0
V20224 n0_10458_12081 n2_10458_12081 0.0
V20225 n0_10458_12114 n2_10458_12114 0.0
V20226 n0_10458_12297 n2_10458_12297 0.0
V20227 n0_10458_12330 n2_10458_12330 0.0
V20228 n0_10458_12513 n2_10458_12513 0.0
V20229 n0_10458_12546 n2_10458_12546 0.0
V20230 n0_10458_12729 n2_10458_12729 0.0
V20231 n0_10458_12762 n2_10458_12762 0.0
V20232 n0_10458_12945 n2_10458_12945 0.0
V20233 n0_10458_12978 n2_10458_12978 0.0
V20234 n0_10458_13161 n2_10458_13161 0.0
V20235 n0_10458_13194 n2_10458_13194 0.0
V20236 n0_10458_13377 n2_10458_13377 0.0
V20237 n0_10458_13410 n2_10458_13410 0.0
V20238 n0_10458_13593 n2_10458_13593 0.0
V20239 n0_10458_13626 n2_10458_13626 0.0
V20240 n0_10458_13640 n2_10458_13640 0.0
V20241 n0_10458_13663 n2_10458_13663 0.0
V20242 n0_10458_13809 n2_10458_13809 0.0
V20243 n0_10458_13842 n2_10458_13842 0.0
V20244 n0_10458_13856 n2_10458_13856 0.0
V20245 n0_10458_13879 n2_10458_13879 0.0
V20246 n0_10458_14025 n2_10458_14025 0.0
V20247 n0_10458_14058 n2_10458_14058 0.0
V20248 n0_10458_14072 n2_10458_14072 0.0
V20249 n0_10458_14079 n2_10458_14079 0.0
V20250 n0_10458_14241 n2_10458_14241 0.0
V20251 n0_10458_14274 n2_10458_14274 0.0
V20252 n0_10458_14457 n2_10458_14457 0.0
V20253 n0_10458_14490 n2_10458_14490 0.0
V20254 n0_10458_14504 n2_10458_14504 0.0
V20255 n0_10458_14673 n2_10458_14673 0.0
V20256 n0_10458_14706 n2_10458_14706 0.0
V20257 n0_10458_14889 n2_10458_14889 0.0
V20258 n0_10458_14922 n2_10458_14922 0.0
V20259 n0_10458_15105 n2_10458_15105 0.0
V20260 n0_10458_15138 n2_10458_15138 0.0
V20261 n0_10458_15321 n2_10458_15321 0.0
V20262 n0_10458_15354 n2_10458_15354 0.0
V20263 n0_10458_15537 n2_10458_15537 0.0
V20264 n0_10458_15570 n2_10458_15570 0.0
V20265 n0_10458_15584 n2_10458_15584 0.0
V20266 n0_10458_15753 n2_10458_15753 0.0
V20267 n0_10458_15786 n2_10458_15786 0.0
V20268 n0_10458_15800 n2_10458_15800 0.0
V20269 n0_10458_15823 n2_10458_15823 0.0
V20270 n0_10458_15969 n2_10458_15969 0.0
V20271 n0_10458_16002 n2_10458_16002 0.0
V20272 n0_10458_16016 n2_10458_16016 0.0
V20273 n0_10458_16185 n2_10458_16185 0.0
V20274 n0_10458_16218 n2_10458_16218 0.0
V20275 n0_10458_16401 n2_10458_16401 0.0
V20276 n0_10458_16434 n2_10458_16434 0.0
V20277 n0_10458_16617 n2_10458_16617 0.0
V20278 n0_10458_16650 n2_10458_16650 0.0
V20279 n0_10458_16833 n2_10458_16833 0.0
V20280 n0_10458_16866 n2_10458_16866 0.0
V20281 n0_10458_17049 n2_10458_17049 0.0
V20282 n0_10458_17082 n2_10458_17082 0.0
V20283 n0_10458_17096 n2_10458_17096 0.0
V20284 n0_10458_17103 n2_10458_17103 0.0
V20285 n0_10458_17119 n2_10458_17119 0.0
V20286 n0_10458_17265 n2_10458_17265 0.0
V20287 n0_10458_17298 n2_10458_17298 0.0
V20288 n0_10458_17312 n2_10458_17312 0.0
V20289 n0_10458_17481 n2_10458_17481 0.0
V20290 n0_10458_17514 n2_10458_17514 0.0
V20291 n0_10458_17697 n2_10458_17697 0.0
V20292 n0_10458_17730 n2_10458_17730 0.0
V20293 n0_10458_17913 n2_10458_17913 0.0
V20294 n0_10458_17946 n2_10458_17946 0.0
V20295 n0_10458_18129 n2_10458_18129 0.0
V20296 n0_10458_18162 n2_10458_18162 0.0
V20297 n0_10458_18345 n2_10458_18345 0.0
V20298 n0_10458_18378 n2_10458_18378 0.0
V20299 n0_10458_18392 n2_10458_18392 0.0
V20300 n0_10458_18561 n2_10458_18561 0.0
V20301 n0_10458_18594 n2_10458_18594 0.0
V20302 n0_10458_18608 n2_10458_18608 0.0
V20303 n0_10458_18777 n2_10458_18777 0.0
V20304 n0_10458_18810 n2_10458_18810 0.0
V20305 n0_10458_18993 n2_10458_18993 0.0
V20306 n0_10458_19026 n2_10458_19026 0.0
V20307 n0_10458_19209 n2_10458_19209 0.0
V20308 n0_10458_19242 n2_10458_19242 0.0
V20309 n0_10458_19256 n2_10458_19256 0.0
V20310 n0_10458_19425 n2_10458_19425 0.0
V20311 n0_10458_19458 n2_10458_19458 0.0
V20312 n0_10458_19641 n2_10458_19641 0.0
V20313 n0_10458_19674 n2_10458_19674 0.0
V20314 n0_10458_19857 n2_10458_19857 0.0
V20315 n0_10458_19890 n2_10458_19890 0.0
V20316 n0_10458_20073 n2_10458_20073 0.0
V20317 n0_10458_20106 n2_10458_20106 0.0
V20318 n0_10458_20289 n2_10458_20289 0.0
V20319 n0_10458_20322 n2_10458_20322 0.0
V20320 n0_10458_20505 n2_10458_20505 0.0
V20321 n0_10458_20538 n2_10458_20538 0.0
V20322 n0_10458_20721 n2_10458_20721 0.0
V20323 n0_10458_20754 n2_10458_20754 0.0
V20324 n0_10458_20937 n2_10458_20937 0.0
V20325 n0_10458_20970 n2_10458_20970 0.0
V20326 n0_10505_417 n2_10505_417 0.0
V20327 n0_10505_450 n2_10505_450 0.0
V20328 n0_10505_1530 n2_10505_1530 0.0
V20329 n0_10505_2647 n2_10505_2647 0.0
V20330 n0_10505_2793 n2_10505_2793 0.0
V20331 n0_10505_3873 n2_10505_3873 0.0
V20332 n0_10505_3906 n2_10505_3906 0.0
V20333 n0_10505_4953 n2_10505_4953 0.0
V20334 n0_10505_4986 n2_10505_4986 0.0
V20335 n0_10505_6033 n2_10505_6033 0.0
V20336 n0_10505_6066 n2_10505_6066 0.0
V20337 n0_10505_7146 n2_10505_7146 0.0
V20338 n0_10505_7160 n2_10505_7160 0.0
V20339 n0_10505_7178 n2_10505_7178 0.0
V20340 n0_10505_8409 n2_10505_8409 0.0
V20341 n0_10505_9489 n2_10505_9489 0.0
V20342 n0_10505_9522 n2_10505_9522 0.0
V20343 n0_10505_10569 n2_10505_10569 0.0
V20344 n0_10505_10602 n2_10505_10602 0.0
V20345 n0_10505_11649 n2_10505_11649 0.0
V20346 n0_10505_11682 n2_10505_11682 0.0
V20347 n0_10505_14025 n2_10505_14025 0.0
V20348 n0_10505_15105 n2_10505_15105 0.0
V20349 n0_10505_15138 n2_10505_15138 0.0
V20350 n0_10505_16185 n2_10505_16185 0.0
V20351 n0_10505_16218 n2_10505_16218 0.0
V20352 n0_10505_17298 n2_10505_17298 0.0
V20353 n0_10505_17312 n2_10505_17312 0.0
V20354 n0_10505_18392 n2_10505_18392 0.0
V20355 n0_10505_19641 n2_10505_19641 0.0
V20356 n0_10505_19674 n2_10505_19674 0.0
V20357 n0_10505_20721 n2_10505_20721 0.0
V20358 n0_10505_20754 n2_10505_20754 0.0
V20359 n0_10554_201 n2_10554_201 0.0
V20360 n0_10554_234 n2_10554_234 0.0
V20361 n0_10554_417 n2_10554_417 0.0
V20362 n0_10554_450 n2_10554_450 0.0
V20363 n0_10554_633 n2_10554_633 0.0
V20364 n0_10554_666 n2_10554_666 0.0
V20365 n0_10554_849 n2_10554_849 0.0
V20366 n0_10554_882 n2_10554_882 0.0
V20367 n0_10554_1065 n2_10554_1065 0.0
V20368 n0_10554_1098 n2_10554_1098 0.0
V20369 n0_10554_1281 n2_10554_1281 0.0
V20370 n0_10554_1314 n2_10554_1314 0.0
V20371 n0_10554_1497 n2_10554_1497 0.0
V20372 n0_10554_1530 n2_10554_1530 0.0
V20373 n0_10554_1713 n2_10554_1713 0.0
V20374 n0_10554_1746 n2_10554_1746 0.0
V20375 n0_10554_1760 n2_10554_1760 0.0
V20376 n0_10554_1783 n2_10554_1783 0.0
V20377 n0_10554_1929 n2_10554_1929 0.0
V20378 n0_10554_1962 n2_10554_1962 0.0
V20379 n0_10554_2145 n2_10554_2145 0.0
V20380 n0_10554_2178 n2_10554_2178 0.0
V20381 n0_10554_2361 n2_10554_2361 0.0
V20382 n0_10554_2394 n2_10554_2394 0.0
V20383 n0_10554_2408 n2_10554_2408 0.0
V20384 n0_10554_2577 n2_10554_2577 0.0
V20385 n0_10554_2610 n2_10554_2610 0.0
V20386 n0_10554_2647 n2_10554_2647 0.0
V20387 n0_10554_2793 n2_10554_2793 0.0
V20388 n0_10554_2826 n2_10554_2826 0.0
V20389 n0_10554_2840 n2_10554_2840 0.0
V20390 n0_10554_2863 n2_10554_2863 0.0
V20391 n0_10554_3009 n2_10554_3009 0.0
V20392 n0_10554_3042 n2_10554_3042 0.0
V20393 n0_10554_3225 n2_10554_3225 0.0
V20394 n0_10554_3258 n2_10554_3258 0.0
V20395 n0_10554_3441 n2_10554_3441 0.0
V20396 n0_10554_3474 n2_10554_3474 0.0
V20397 n0_10554_3488 n2_10554_3488 0.0
V20398 n0_10554_3511 n2_10554_3511 0.0
V20399 n0_10554_3657 n2_10554_3657 0.0
V20400 n0_10554_3690 n2_10554_3690 0.0
V20401 n0_10554_3873 n2_10554_3873 0.0
V20402 n0_10554_3906 n2_10554_3906 0.0
V20403 n0_10554_4089 n2_10554_4089 0.0
V20404 n0_10554_4122 n2_10554_4122 0.0
V20405 n0_10554_4136 n2_10554_4136 0.0
V20406 n0_10554_4159 n2_10554_4159 0.0
V20407 n0_10554_4305 n2_10554_4305 0.0
V20408 n0_10554_4338 n2_10554_4338 0.0
V20409 n0_10554_4521 n2_10554_4521 0.0
V20410 n0_10554_4554 n2_10554_4554 0.0
V20411 n0_10554_4568 n2_10554_4568 0.0
V20412 n0_10554_4591 n2_10554_4591 0.0
V20413 n0_10554_4737 n2_10554_4737 0.0
V20414 n0_10554_4770 n2_10554_4770 0.0
V20415 n0_10554_4953 n2_10554_4953 0.0
V20416 n0_10554_4986 n2_10554_4986 0.0
V20417 n0_10554_5169 n2_10554_5169 0.0
V20418 n0_10554_5202 n2_10554_5202 0.0
V20419 n0_10554_5239 n2_10554_5239 0.0
V20420 n0_10554_5385 n2_10554_5385 0.0
V20421 n0_10554_5418 n2_10554_5418 0.0
V20422 n0_10554_5432 n2_10554_5432 0.0
V20423 n0_10554_5455 n2_10554_5455 0.0
V20424 n0_10554_5601 n2_10554_5601 0.0
V20425 n0_10554_5634 n2_10554_5634 0.0
V20426 n0_10554_5817 n2_10554_5817 0.0
V20427 n0_10554_5850 n2_10554_5850 0.0
V20428 n0_10554_6033 n2_10554_6033 0.0
V20429 n0_10554_6066 n2_10554_6066 0.0
V20430 n0_10554_6249 n2_10554_6249 0.0
V20431 n0_10554_6282 n2_10554_6282 0.0
V20432 n0_10554_6465 n2_10554_6465 0.0
V20433 n0_10554_6498 n2_10554_6498 0.0
V20434 n0_10554_6512 n2_10554_6512 0.0
V20435 n0_10554_6535 n2_10554_6535 0.0
V20436 n0_10554_6681 n2_10554_6681 0.0
V20437 n0_10554_6714 n2_10554_6714 0.0
V20438 n0_10554_6751 n2_10554_6751 0.0
V20439 n0_10554_6897 n2_10554_6897 0.0
V20440 n0_10554_6930 n2_10554_6930 0.0
V20441 n0_10554_6944 n2_10554_6944 0.0
V20442 n0_10554_6967 n2_10554_6967 0.0
V20443 n0_10554_7113 n2_10554_7113 0.0
V20444 n0_10554_7146 n2_10554_7146 0.0
V20445 n0_10554_7160 n2_10554_7160 0.0
V20446 n0_10554_7178 n2_10554_7178 0.0
V20447 n0_10554_7329 n2_10554_7329 0.0
V20448 n0_10554_7362 n2_10554_7362 0.0
V20449 n0_10554_7376 n2_10554_7376 0.0
V20450 n0_10554_7399 n2_10554_7399 0.0
V20451 n0_10554_7545 n2_10554_7545 0.0
V20452 n0_10554_7578 n2_10554_7578 0.0
V20453 n0_10554_7761 n2_10554_7761 0.0
V20454 n0_10554_7794 n2_10554_7794 0.0
V20455 n0_10554_7977 n2_10554_7977 0.0
V20456 n0_10554_8010 n2_10554_8010 0.0
V20457 n0_10554_8193 n2_10554_8193 0.0
V20458 n0_10554_8226 n2_10554_8226 0.0
V20459 n0_10554_8409 n2_10554_8409 0.0
V20460 n0_10554_8442 n2_10554_8442 0.0
V20461 n0_10554_8625 n2_10554_8625 0.0
V20462 n0_10554_8658 n2_10554_8658 0.0
V20463 n0_10554_8841 n2_10554_8841 0.0
V20464 n0_10554_8874 n2_10554_8874 0.0
V20465 n0_10554_9057 n2_10554_9057 0.0
V20466 n0_10554_9090 n2_10554_9090 0.0
V20467 n0_10554_9273 n2_10554_9273 0.0
V20468 n0_10554_9306 n2_10554_9306 0.0
V20469 n0_10554_9489 n2_10554_9489 0.0
V20470 n0_10554_9522 n2_10554_9522 0.0
V20471 n0_10554_9705 n2_10554_9705 0.0
V20472 n0_10554_9738 n2_10554_9738 0.0
V20473 n0_10554_9921 n2_10554_9921 0.0
V20474 n0_10554_9954 n2_10554_9954 0.0
V20475 n0_10554_10137 n2_10554_10137 0.0
V20476 n0_10554_10170 n2_10554_10170 0.0
V20477 n0_10554_10353 n2_10554_10353 0.0
V20478 n0_10554_10386 n2_10554_10386 0.0
V20479 n0_10554_10569 n2_10554_10569 0.0
V20480 n0_10554_10602 n2_10554_10602 0.0
V20481 n0_10554_10785 n2_10554_10785 0.0
V20482 n0_10554_10818 n2_10554_10818 0.0
V20483 n0_10554_11001 n2_10554_11001 0.0
V20484 n0_10554_11034 n2_10554_11034 0.0
V20485 n0_10554_11217 n2_10554_11217 0.0
V20486 n0_10554_11250 n2_10554_11250 0.0
V20487 n0_10554_11433 n2_10554_11433 0.0
V20488 n0_10554_11466 n2_10554_11466 0.0
V20489 n0_10554_11649 n2_10554_11649 0.0
V20490 n0_10554_11682 n2_10554_11682 0.0
V20491 n0_10554_11865 n2_10554_11865 0.0
V20492 n0_10554_11898 n2_10554_11898 0.0
V20493 n0_10554_12081 n2_10554_12081 0.0
V20494 n0_10554_12114 n2_10554_12114 0.0
V20495 n0_10554_12297 n2_10554_12297 0.0
V20496 n0_10554_12330 n2_10554_12330 0.0
V20497 n0_10554_12513 n2_10554_12513 0.0
V20498 n0_10554_12546 n2_10554_12546 0.0
V20499 n0_10554_12729 n2_10554_12729 0.0
V20500 n0_10554_12762 n2_10554_12762 0.0
V20501 n0_10554_12945 n2_10554_12945 0.0
V20502 n0_10554_12978 n2_10554_12978 0.0
V20503 n0_10554_13161 n2_10554_13161 0.0
V20504 n0_10554_13194 n2_10554_13194 0.0
V20505 n0_10554_13377 n2_10554_13377 0.0
V20506 n0_10554_13410 n2_10554_13410 0.0
V20507 n0_10554_13593 n2_10554_13593 0.0
V20508 n0_10554_13626 n2_10554_13626 0.0
V20509 n0_10554_13640 n2_10554_13640 0.0
V20510 n0_10554_13663 n2_10554_13663 0.0
V20511 n0_10554_13809 n2_10554_13809 0.0
V20512 n0_10554_13842 n2_10554_13842 0.0
V20513 n0_10554_13856 n2_10554_13856 0.0
V20514 n0_10554_13879 n2_10554_13879 0.0
V20515 n0_10554_14025 n2_10554_14025 0.0
V20516 n0_10554_14058 n2_10554_14058 0.0
V20517 n0_10554_14072 n2_10554_14072 0.0
V20518 n0_10554_14079 n2_10554_14079 0.0
V20519 n0_10554_14241 n2_10554_14241 0.0
V20520 n0_10554_14274 n2_10554_14274 0.0
V20521 n0_10554_14457 n2_10554_14457 0.0
V20522 n0_10554_14490 n2_10554_14490 0.0
V20523 n0_10554_14504 n2_10554_14504 0.0
V20524 n0_10554_14673 n2_10554_14673 0.0
V20525 n0_10554_14706 n2_10554_14706 0.0
V20526 n0_10554_14889 n2_10554_14889 0.0
V20527 n0_10554_14922 n2_10554_14922 0.0
V20528 n0_10554_15105 n2_10554_15105 0.0
V20529 n0_10554_15138 n2_10554_15138 0.0
V20530 n0_10554_15321 n2_10554_15321 0.0
V20531 n0_10554_15354 n2_10554_15354 0.0
V20532 n0_10554_15537 n2_10554_15537 0.0
V20533 n0_10554_15570 n2_10554_15570 0.0
V20534 n0_10554_15584 n2_10554_15584 0.0
V20535 n0_10554_15753 n2_10554_15753 0.0
V20536 n0_10554_15786 n2_10554_15786 0.0
V20537 n0_10554_15800 n2_10554_15800 0.0
V20538 n0_10554_15823 n2_10554_15823 0.0
V20539 n0_10554_15969 n2_10554_15969 0.0
V20540 n0_10554_16002 n2_10554_16002 0.0
V20541 n0_10554_16016 n2_10554_16016 0.0
V20542 n0_10554_16185 n2_10554_16185 0.0
V20543 n0_10554_16218 n2_10554_16218 0.0
V20544 n0_10554_16401 n2_10554_16401 0.0
V20545 n0_10554_16434 n2_10554_16434 0.0
V20546 n0_10554_16617 n2_10554_16617 0.0
V20547 n0_10554_16650 n2_10554_16650 0.0
V20548 n0_10554_16833 n2_10554_16833 0.0
V20549 n0_10554_16866 n2_10554_16866 0.0
V20550 n0_10554_17049 n2_10554_17049 0.0
V20551 n0_10554_17082 n2_10554_17082 0.0
V20552 n0_10554_17096 n2_10554_17096 0.0
V20553 n0_10554_17103 n2_10554_17103 0.0
V20554 n0_10554_17119 n2_10554_17119 0.0
V20555 n0_10554_17265 n2_10554_17265 0.0
V20556 n0_10554_17298 n2_10554_17298 0.0
V20557 n0_10554_17312 n2_10554_17312 0.0
V20558 n0_10554_17481 n2_10554_17481 0.0
V20559 n0_10554_17514 n2_10554_17514 0.0
V20560 n0_10554_17697 n2_10554_17697 0.0
V20561 n0_10554_17730 n2_10554_17730 0.0
V20562 n0_10554_17913 n2_10554_17913 0.0
V20563 n0_10554_17946 n2_10554_17946 0.0
V20564 n0_10554_18129 n2_10554_18129 0.0
V20565 n0_10554_18162 n2_10554_18162 0.0
V20566 n0_10554_18345 n2_10554_18345 0.0
V20567 n0_10554_18378 n2_10554_18378 0.0
V20568 n0_10554_18392 n2_10554_18392 0.0
V20569 n0_10554_18561 n2_10554_18561 0.0
V20570 n0_10554_18594 n2_10554_18594 0.0
V20571 n0_10554_18608 n2_10554_18608 0.0
V20572 n0_10554_18777 n2_10554_18777 0.0
V20573 n0_10554_18810 n2_10554_18810 0.0
V20574 n0_10554_18993 n2_10554_18993 0.0
V20575 n0_10554_19026 n2_10554_19026 0.0
V20576 n0_10554_19209 n2_10554_19209 0.0
V20577 n0_10554_19242 n2_10554_19242 0.0
V20578 n0_10554_19256 n2_10554_19256 0.0
V20579 n0_10554_19425 n2_10554_19425 0.0
V20580 n0_10554_19458 n2_10554_19458 0.0
V20581 n0_10554_19641 n2_10554_19641 0.0
V20582 n0_10554_19674 n2_10554_19674 0.0
V20583 n0_10554_19857 n2_10554_19857 0.0
V20584 n0_10554_19890 n2_10554_19890 0.0
V20585 n0_10554_20073 n2_10554_20073 0.0
V20586 n0_10554_20106 n2_10554_20106 0.0
V20587 n0_10554_20289 n2_10554_20289 0.0
V20588 n0_10554_20322 n2_10554_20322 0.0
V20589 n0_10554_20505 n2_10554_20505 0.0
V20590 n0_10554_20538 n2_10554_20538 0.0
V20591 n0_10554_20721 n2_10554_20721 0.0
V20592 n0_10554_20754 n2_10554_20754 0.0
V20593 n0_10554_20937 n2_10554_20937 0.0
V20594 n0_10554_20970 n2_10554_20970 0.0
V20595 n0_10646_201 n2_10646_201 0.0
V20596 n0_10646_234 n2_10646_234 0.0
V20597 n0_10646_417 n2_10646_417 0.0
V20598 n0_10646_450 n2_10646_450 0.0
V20599 n0_10646_633 n2_10646_633 0.0
V20600 n0_10646_666 n2_10646_666 0.0
V20601 n0_10646_849 n2_10646_849 0.0
V20602 n0_10646_882 n2_10646_882 0.0
V20603 n0_10646_1065 n2_10646_1065 0.0
V20604 n0_10646_1098 n2_10646_1098 0.0
V20605 n0_10646_1281 n2_10646_1281 0.0
V20606 n0_10646_1314 n2_10646_1314 0.0
V20607 n0_10646_1497 n2_10646_1497 0.0
V20608 n0_10646_1530 n2_10646_1530 0.0
V20609 n0_10646_1713 n2_10646_1713 0.0
V20610 n0_10646_1746 n2_10646_1746 0.0
V20611 n0_10646_1760 n2_10646_1760 0.0
V20612 n0_10646_1783 n2_10646_1783 0.0
V20613 n0_10646_1929 n2_10646_1929 0.0
V20614 n0_10646_1962 n2_10646_1962 0.0
V20615 n0_10646_2145 n2_10646_2145 0.0
V20616 n0_10646_2178 n2_10646_2178 0.0
V20617 n0_10646_2361 n2_10646_2361 0.0
V20618 n0_10646_2394 n2_10646_2394 0.0
V20619 n0_10646_2408 n2_10646_2408 0.0
V20620 n0_10646_2577 n2_10646_2577 0.0
V20621 n0_10646_2610 n2_10646_2610 0.0
V20622 n0_10646_2647 n2_10646_2647 0.0
V20623 n0_10646_2793 n2_10646_2793 0.0
V20624 n0_10646_2826 n2_10646_2826 0.0
V20625 n0_10646_2840 n2_10646_2840 0.0
V20626 n0_10646_2863 n2_10646_2863 0.0
V20627 n0_10646_3009 n2_10646_3009 0.0
V20628 n0_10646_3042 n2_10646_3042 0.0
V20629 n0_10646_3225 n2_10646_3225 0.0
V20630 n0_10646_3258 n2_10646_3258 0.0
V20631 n0_10646_3441 n2_10646_3441 0.0
V20632 n0_10646_3474 n2_10646_3474 0.0
V20633 n0_10646_3488 n2_10646_3488 0.0
V20634 n0_10646_3511 n2_10646_3511 0.0
V20635 n0_10646_3657 n2_10646_3657 0.0
V20636 n0_10646_3690 n2_10646_3690 0.0
V20637 n0_10646_3873 n2_10646_3873 0.0
V20638 n0_10646_3906 n2_10646_3906 0.0
V20639 n0_10646_4089 n2_10646_4089 0.0
V20640 n0_10646_4122 n2_10646_4122 0.0
V20641 n0_10646_4136 n2_10646_4136 0.0
V20642 n0_10646_4159 n2_10646_4159 0.0
V20643 n0_10646_4305 n2_10646_4305 0.0
V20644 n0_10646_4338 n2_10646_4338 0.0
V20645 n0_10646_4521 n2_10646_4521 0.0
V20646 n0_10646_4554 n2_10646_4554 0.0
V20647 n0_10646_4568 n2_10646_4568 0.0
V20648 n0_10646_4591 n2_10646_4591 0.0
V20649 n0_10646_4737 n2_10646_4737 0.0
V20650 n0_10646_4770 n2_10646_4770 0.0
V20651 n0_10646_4953 n2_10646_4953 0.0
V20652 n0_10646_5169 n2_10646_5169 0.0
V20653 n0_10646_5202 n2_10646_5202 0.0
V20654 n0_10646_5239 n2_10646_5239 0.0
V20655 n0_10646_5385 n2_10646_5385 0.0
V20656 n0_10646_5418 n2_10646_5418 0.0
V20657 n0_10646_5432 n2_10646_5432 0.0
V20658 n0_10646_5455 n2_10646_5455 0.0
V20659 n0_10646_5601 n2_10646_5601 0.0
V20660 n0_10646_5634 n2_10646_5634 0.0
V20661 n0_10646_5817 n2_10646_5817 0.0
V20662 n0_10646_5850 n2_10646_5850 0.0
V20663 n0_10646_6033 n2_10646_6033 0.0
V20664 n0_10646_6066 n2_10646_6066 0.0
V20665 n0_10646_6249 n2_10646_6249 0.0
V20666 n0_10646_6282 n2_10646_6282 0.0
V20667 n0_10646_6465 n2_10646_6465 0.0
V20668 n0_10646_6498 n2_10646_6498 0.0
V20669 n0_10646_6512 n2_10646_6512 0.0
V20670 n0_10646_6535 n2_10646_6535 0.0
V20671 n0_10646_6681 n2_10646_6681 0.0
V20672 n0_10646_6714 n2_10646_6714 0.0
V20673 n0_10646_6751 n2_10646_6751 0.0
V20674 n0_10646_6897 n2_10646_6897 0.0
V20675 n0_10646_6930 n2_10646_6930 0.0
V20676 n0_10646_6944 n2_10646_6944 0.0
V20677 n0_10646_6967 n2_10646_6967 0.0
V20678 n0_10646_7113 n2_10646_7113 0.0
V20679 n0_10646_7146 n2_10646_7146 0.0
V20680 n0_10646_7160 n2_10646_7160 0.0
V20681 n0_10646_7178 n2_10646_7178 0.0
V20682 n0_10646_7329 n2_10646_7329 0.0
V20683 n0_10646_7362 n2_10646_7362 0.0
V20684 n0_10646_7376 n2_10646_7376 0.0
V20685 n0_10646_7399 n2_10646_7399 0.0
V20686 n0_10646_7545 n2_10646_7545 0.0
V20687 n0_10646_7578 n2_10646_7578 0.0
V20688 n0_10646_7761 n2_10646_7761 0.0
V20689 n0_10646_7794 n2_10646_7794 0.0
V20690 n0_10646_7977 n2_10646_7977 0.0
V20691 n0_10646_8010 n2_10646_8010 0.0
V20692 n0_10646_8193 n2_10646_8193 0.0
V20693 n0_10646_8226 n2_10646_8226 0.0
V20694 n0_10646_8409 n2_10646_8409 0.0
V20695 n0_10646_8442 n2_10646_8442 0.0
V20696 n0_10646_8613 n2_10646_8613 0.0
V20697 n0_10646_8625 n2_10646_8625 0.0
V20698 n0_10646_8658 n2_10646_8658 0.0
V20699 n0_10646_8841 n2_10646_8841 0.0
V20700 n0_10646_8874 n2_10646_8874 0.0
V20701 n0_10646_9057 n2_10646_9057 0.0
V20702 n0_10646_9090 n2_10646_9090 0.0
V20703 n0_10646_9190 n2_10646_9190 0.0
V20704 n0_10646_9273 n2_10646_9273 0.0
V20705 n0_10646_9306 n2_10646_9306 0.0
V20706 n0_10646_9489 n2_10646_9489 0.0
V20707 n0_10646_9522 n2_10646_9522 0.0
V20708 n0_10646_9705 n2_10646_9705 0.0
V20709 n0_10646_9738 n2_10646_9738 0.0
V20710 n0_10646_9921 n2_10646_9921 0.0
V20711 n0_10646_9954 n2_10646_9954 0.0
V20712 n0_10646_10137 n2_10646_10137 0.0
V20713 n0_10646_10170 n2_10646_10170 0.0
V20714 n0_10646_10353 n2_10646_10353 0.0
V20715 n0_10646_10386 n2_10646_10386 0.0
V20716 n0_10646_10569 n2_10646_10569 0.0
V20717 n0_10646_10785 n2_10646_10785 0.0
V20718 n0_10646_10818 n2_10646_10818 0.0
V20719 n0_10646_11001 n2_10646_11001 0.0
V20720 n0_10646_11034 n2_10646_11034 0.0
V20721 n0_10646_11217 n2_10646_11217 0.0
V20722 n0_10646_11250 n2_10646_11250 0.0
V20723 n0_10646_11433 n2_10646_11433 0.0
V20724 n0_10646_11466 n2_10646_11466 0.0
V20725 n0_10646_11649 n2_10646_11649 0.0
V20726 n0_10646_11682 n2_10646_11682 0.0
V20727 n0_10646_11865 n2_10646_11865 0.0
V20728 n0_10646_11898 n2_10646_11898 0.0
V20729 n0_10646_12004 n2_10646_12004 0.0
V20730 n0_10646_12081 n2_10646_12081 0.0
V20731 n0_10646_12114 n2_10646_12114 0.0
V20732 n0_10646_12297 n2_10646_12297 0.0
V20733 n0_10646_12330 n2_10646_12330 0.0
V20734 n0_10646_12513 n2_10646_12513 0.0
V20735 n0_10646_12546 n2_10646_12546 0.0
V20736 n0_10646_12566 n2_10646_12566 0.0
V20737 n0_10646_12729 n2_10646_12729 0.0
V20738 n0_10646_12762 n2_10646_12762 0.0
V20739 n0_10646_12945 n2_10646_12945 0.0
V20740 n0_10646_12978 n2_10646_12978 0.0
V20741 n0_10646_13161 n2_10646_13161 0.0
V20742 n0_10646_13194 n2_10646_13194 0.0
V20743 n0_10646_13377 n2_10646_13377 0.0
V20744 n0_10646_13410 n2_10646_13410 0.0
V20745 n0_10646_13593 n2_10646_13593 0.0
V20746 n0_10646_13626 n2_10646_13626 0.0
V20747 n0_10646_13640 n2_10646_13640 0.0
V20748 n0_10646_13663 n2_10646_13663 0.0
V20749 n0_10646_13809 n2_10646_13809 0.0
V20750 n0_10646_13842 n2_10646_13842 0.0
V20751 n0_10646_13856 n2_10646_13856 0.0
V20752 n0_10646_13879 n2_10646_13879 0.0
V20753 n0_10646_14025 n2_10646_14025 0.0
V20754 n0_10646_14058 n2_10646_14058 0.0
V20755 n0_10646_14072 n2_10646_14072 0.0
V20756 n0_10646_14079 n2_10646_14079 0.0
V20757 n0_10646_14241 n2_10646_14241 0.0
V20758 n0_10646_14274 n2_10646_14274 0.0
V20759 n0_10646_14457 n2_10646_14457 0.0
V20760 n0_10646_14490 n2_10646_14490 0.0
V20761 n0_10646_14504 n2_10646_14504 0.0
V20762 n0_10646_14673 n2_10646_14673 0.0
V20763 n0_10646_14706 n2_10646_14706 0.0
V20764 n0_10646_14889 n2_10646_14889 0.0
V20765 n0_10646_14922 n2_10646_14922 0.0
V20766 n0_10646_15138 n2_10646_15138 0.0
V20767 n0_10646_15321 n2_10646_15321 0.0
V20768 n0_10646_15354 n2_10646_15354 0.0
V20769 n0_10646_15537 n2_10646_15537 0.0
V20770 n0_10646_15570 n2_10646_15570 0.0
V20771 n0_10646_15584 n2_10646_15584 0.0
V20772 n0_10646_15753 n2_10646_15753 0.0
V20773 n0_10646_15786 n2_10646_15786 0.0
V20774 n0_10646_15800 n2_10646_15800 0.0
V20775 n0_10646_15823 n2_10646_15823 0.0
V20776 n0_10646_15969 n2_10646_15969 0.0
V20777 n0_10646_16002 n2_10646_16002 0.0
V20778 n0_10646_16016 n2_10646_16016 0.0
V20779 n0_10646_16185 n2_10646_16185 0.0
V20780 n0_10646_16401 n2_10646_16401 0.0
V20781 n0_10646_16434 n2_10646_16434 0.0
V20782 n0_10646_16617 n2_10646_16617 0.0
V20783 n0_10646_16650 n2_10646_16650 0.0
V20784 n0_10646_16833 n2_10646_16833 0.0
V20785 n0_10646_16866 n2_10646_16866 0.0
V20786 n0_10646_17049 n2_10646_17049 0.0
V20787 n0_10646_17082 n2_10646_17082 0.0
V20788 n0_10646_17096 n2_10646_17096 0.0
V20789 n0_10646_17103 n2_10646_17103 0.0
V20790 n0_10646_17119 n2_10646_17119 0.0
V20791 n0_10646_17265 n2_10646_17265 0.0
V20792 n0_10646_17298 n2_10646_17298 0.0
V20793 n0_10646_17312 n2_10646_17312 0.0
V20794 n0_10646_17481 n2_10646_17481 0.0
V20795 n0_10646_17514 n2_10646_17514 0.0
V20796 n0_10646_17697 n2_10646_17697 0.0
V20797 n0_10646_17730 n2_10646_17730 0.0
V20798 n0_10646_17913 n2_10646_17913 0.0
V20799 n0_10646_17946 n2_10646_17946 0.0
V20800 n0_10646_18129 n2_10646_18129 0.0
V20801 n0_10646_18162 n2_10646_18162 0.0
V20802 n0_10646_18345 n2_10646_18345 0.0
V20803 n0_10646_18378 n2_10646_18378 0.0
V20804 n0_10646_18392 n2_10646_18392 0.0
V20805 n0_10646_18561 n2_10646_18561 0.0
V20806 n0_10646_18594 n2_10646_18594 0.0
V20807 n0_10646_18608 n2_10646_18608 0.0
V20808 n0_10646_18777 n2_10646_18777 0.0
V20809 n0_10646_18810 n2_10646_18810 0.0
V20810 n0_10646_18993 n2_10646_18993 0.0
V20811 n0_10646_19026 n2_10646_19026 0.0
V20812 n0_10646_19209 n2_10646_19209 0.0
V20813 n0_10646_19242 n2_10646_19242 0.0
V20814 n0_10646_19256 n2_10646_19256 0.0
V20815 n0_10646_19425 n2_10646_19425 0.0
V20816 n0_10646_19458 n2_10646_19458 0.0
V20817 n0_10646_19641 n2_10646_19641 0.0
V20818 n0_10646_19674 n2_10646_19674 0.0
V20819 n0_10646_19857 n2_10646_19857 0.0
V20820 n0_10646_19890 n2_10646_19890 0.0
V20821 n0_10646_20073 n2_10646_20073 0.0
V20822 n0_10646_20106 n2_10646_20106 0.0
V20823 n0_10646_20289 n2_10646_20289 0.0
V20824 n0_10646_20322 n2_10646_20322 0.0
V20825 n0_10646_20505 n2_10646_20505 0.0
V20826 n0_10646_20538 n2_10646_20538 0.0
V20827 n0_10646_20754 n2_10646_20754 0.0
V20828 n0_10646_20937 n2_10646_20937 0.0
V20829 n0_10646_20970 n2_10646_20970 0.0
V20830 n0_11491_9489 n2_11491_9489 0.0
V20831 n0_11491_9522 n2_11491_9522 0.0
V20832 n0_11491_9705 n2_11491_9705 0.0
V20833 n0_11491_9738 n2_11491_9738 0.0
V20834 n0_11491_9921 n2_11491_9921 0.0
V20835 n0_11491_9954 n2_11491_9954 0.0
V20836 n0_11491_10137 n2_11491_10137 0.0
V20837 n0_11491_10170 n2_11491_10170 0.0
V20838 n0_11491_10353 n2_11491_10353 0.0
V20839 n0_11491_10386 n2_11491_10386 0.0
V20840 n0_11491_10569 n2_11491_10569 0.0
V20841 n0_11491_10785 n2_11491_10785 0.0
V20842 n0_11491_10818 n2_11491_10818 0.0
V20843 n0_11491_11001 n2_11491_11001 0.0
V20844 n0_11491_11034 n2_11491_11034 0.0
V20845 n0_11491_11217 n2_11491_11217 0.0
V20846 n0_11491_11250 n2_11491_11250 0.0
V20847 n0_11491_11433 n2_11491_11433 0.0
V20848 n0_11491_11466 n2_11491_11466 0.0
V20849 n0_11491_11649 n2_11491_11649 0.0
V20850 n0_11491_11682 n2_11491_11682 0.0
V20851 n0_11630_10569 n2_11630_10569 0.0
V20852 n0_11630_10602 n2_11630_10602 0.0
V20853 n0_11679_9705 n2_11679_9705 0.0
V20854 n0_11679_9738 n2_11679_9738 0.0
V20855 n0_11679_9921 n2_11679_9921 0.0
V20856 n0_11679_9954 n2_11679_9954 0.0
V20857 n0_11679_10034 n2_11679_10034 0.0
V20858 n0_11679_10137 n2_11679_10137 0.0
V20859 n0_11679_10170 n2_11679_10170 0.0
V20860 n0_11679_10353 n2_11679_10353 0.0
V20861 n0_11679_10386 n2_11679_10386 0.0
V20862 n0_11679_10569 n2_11679_10569 0.0
V20863 n0_11679_10602 n2_11679_10602 0.0
V20864 n0_11679_10785 n2_11679_10785 0.0
V20865 n0_11679_10818 n2_11679_10818 0.0
V20866 n0_11679_11001 n2_11679_11001 0.0
V20867 n0_11679_11034 n2_11679_11034 0.0
V20868 n0_11679_11160 n2_11679_11160 0.0
V20869 n0_11679_11217 n2_11679_11217 0.0
V20870 n0_11679_11250 n2_11679_11250 0.0
V20871 n0_11679_11433 n2_11679_11433 0.0
V20872 n0_11679_11466 n2_11679_11466 0.0
V20873 n0_12616_201 n2_12616_201 0.0
V20874 n0_12616_234 n2_12616_234 0.0
V20875 n0_12616_417 n2_12616_417 0.0
V20876 n0_12616_450 n2_12616_450 0.0
V20877 n0_12616_633 n2_12616_633 0.0
V20878 n0_12616_666 n2_12616_666 0.0
V20879 n0_12616_849 n2_12616_849 0.0
V20880 n0_12616_882 n2_12616_882 0.0
V20881 n0_12616_1065 n2_12616_1065 0.0
V20882 n0_12616_1098 n2_12616_1098 0.0
V20883 n0_12616_1281 n2_12616_1281 0.0
V20884 n0_12616_1314 n2_12616_1314 0.0
V20885 n0_12616_1497 n2_12616_1497 0.0
V20886 n0_12616_1530 n2_12616_1530 0.0
V20887 n0_12616_1713 n2_12616_1713 0.0
V20888 n0_12616_1746 n2_12616_1746 0.0
V20889 n0_12616_1783 n2_12616_1783 0.0
V20890 n0_12616_1929 n2_12616_1929 0.0
V20891 n0_12616_1962 n2_12616_1962 0.0
V20892 n0_12616_2145 n2_12616_2145 0.0
V20893 n0_12616_2178 n2_12616_2178 0.0
V20894 n0_12616_2361 n2_12616_2361 0.0
V20895 n0_12616_2394 n2_12616_2394 0.0
V20896 n0_12616_2431 n2_12616_2431 0.0
V20897 n0_12616_2577 n2_12616_2577 0.0
V20898 n0_12616_2610 n2_12616_2610 0.0
V20899 n0_12616_2793 n2_12616_2793 0.0
V20900 n0_12616_2826 n2_12616_2826 0.0
V20901 n0_12616_2863 n2_12616_2863 0.0
V20902 n0_12616_3009 n2_12616_3009 0.0
V20903 n0_12616_3042 n2_12616_3042 0.0
V20904 n0_12616_3225 n2_12616_3225 0.0
V20905 n0_12616_3258 n2_12616_3258 0.0
V20906 n0_12616_3441 n2_12616_3441 0.0
V20907 n0_12616_3474 n2_12616_3474 0.0
V20908 n0_12616_3511 n2_12616_3511 0.0
V20909 n0_12616_3657 n2_12616_3657 0.0
V20910 n0_12616_3690 n2_12616_3690 0.0
V20911 n0_12616_3873 n2_12616_3873 0.0
V20912 n0_12616_3906 n2_12616_3906 0.0
V20913 n0_12616_3943 n2_12616_3943 0.0
V20914 n0_12616_4089 n2_12616_4089 0.0
V20915 n0_12616_4122 n2_12616_4122 0.0
V20916 n0_12616_4159 n2_12616_4159 0.0
V20917 n0_12616_4305 n2_12616_4305 0.0
V20918 n0_12616_4338 n2_12616_4338 0.0
V20919 n0_12616_4521 n2_12616_4521 0.0
V20920 n0_12616_4554 n2_12616_4554 0.0
V20921 n0_12616_4591 n2_12616_4591 0.0
V20922 n0_12616_4737 n2_12616_4737 0.0
V20923 n0_12616_4770 n2_12616_4770 0.0
V20924 n0_12616_4953 n2_12616_4953 0.0
V20925 n0_12616_5023 n2_12616_5023 0.0
V20926 n0_12616_5169 n2_12616_5169 0.0
V20927 n0_12616_5202 n2_12616_5202 0.0
V20928 n0_12616_5239 n2_12616_5239 0.0
V20929 n0_12616_5385 n2_12616_5385 0.0
V20930 n0_12616_5418 n2_12616_5418 0.0
V20931 n0_12616_5601 n2_12616_5601 0.0
V20932 n0_12616_5634 n2_12616_5634 0.0
V20933 n0_12616_5671 n2_12616_5671 0.0
V20934 n0_12616_5817 n2_12616_5817 0.0
V20935 n0_12616_5850 n2_12616_5850 0.0
V20936 n0_12616_6033 n2_12616_6033 0.0
V20937 n0_12616_6066 n2_12616_6066 0.0
V20938 n0_12616_6249 n2_12616_6249 0.0
V20939 n0_12616_6282 n2_12616_6282 0.0
V20940 n0_12616_6319 n2_12616_6319 0.0
V20941 n0_12616_6465 n2_12616_6465 0.0
V20942 n0_12616_6498 n2_12616_6498 0.0
V20943 n0_12616_6681 n2_12616_6681 0.0
V20944 n0_12616_6714 n2_12616_6714 0.0
V20945 n0_12616_6751 n2_12616_6751 0.0
V20946 n0_12616_6897 n2_12616_6897 0.0
V20947 n0_12616_6930 n2_12616_6930 0.0
V20948 n0_12616_6967 n2_12616_6967 0.0
V20949 n0_12616_7113 n2_12616_7113 0.0
V20950 n0_12616_7146 n2_12616_7146 0.0
V20951 n0_12616_7178 n2_12616_7178 0.0
V20952 n0_12616_7329 n2_12616_7329 0.0
V20953 n0_12616_7362 n2_12616_7362 0.0
V20954 n0_12616_7399 n2_12616_7399 0.0
V20955 n0_12616_7545 n2_12616_7545 0.0
V20956 n0_12616_7578 n2_12616_7578 0.0
V20957 n0_12616_7761 n2_12616_7761 0.0
V20958 n0_12616_7794 n2_12616_7794 0.0
V20959 n0_12616_7831 n2_12616_7831 0.0
V20960 n0_12616_7977 n2_12616_7977 0.0
V20961 n0_12616_8010 n2_12616_8010 0.0
V20962 n0_12616_8193 n2_12616_8193 0.0
V20963 n0_12616_8226 n2_12616_8226 0.0
V20964 n0_12616_8409 n2_12616_8409 0.0
V20965 n0_12616_8442 n2_12616_8442 0.0
V20966 n0_12616_8625 n2_12616_8625 0.0
V20967 n0_12616_8658 n2_12616_8658 0.0
V20968 n0_12616_8695 n2_12616_8695 0.0
V20969 n0_12616_8841 n2_12616_8841 0.0
V20970 n0_12616_8874 n2_12616_8874 0.0
V20971 n0_12616_8911 n2_12616_8911 0.0
V20972 n0_12616_8948 n2_12616_8948 0.0
V20973 n0_12616_9057 n2_12616_9057 0.0
V20974 n0_12616_9090 n2_12616_9090 0.0
V20975 n0_12616_9273 n2_12616_9273 0.0
V20976 n0_12616_9306 n2_12616_9306 0.0
V20977 n0_12616_9489 n2_12616_9489 0.0
V20978 n0_12616_9522 n2_12616_9522 0.0
V20979 n0_12616_9705 n2_12616_9705 0.0
V20980 n0_12616_9738 n2_12616_9738 0.0
V20981 n0_12616_9775 n2_12616_9775 0.0
V20982 n0_12616_9921 n2_12616_9921 0.0
V20983 n0_12616_9954 n2_12616_9954 0.0
V20984 n0_12616_9991 n2_12616_9991 0.0
V20985 n0_12616_10034 n2_12616_10034 0.0
V20986 n0_12616_10137 n2_12616_10137 0.0
V20987 n0_12616_10170 n2_12616_10170 0.0
V20988 n0_12616_10353 n2_12616_10353 0.0
V20989 n0_12616_10386 n2_12616_10386 0.0
V20990 n0_12616_10569 n2_12616_10569 0.0
V20991 n0_12616_10785 n2_12616_10785 0.0
V20992 n0_12616_10818 n2_12616_10818 0.0
V20993 n0_12616_10832 n2_12616_10832 0.0
V20994 n0_12616_11001 n2_12616_11001 0.0
V20995 n0_12616_11034 n2_12616_11034 0.0
V20996 n0_12616_11048 n2_12616_11048 0.0
V20997 n0_12616_11160 n2_12616_11160 0.0
V20998 n0_12616_11217 n2_12616_11217 0.0
V20999 n0_12616_11250 n2_12616_11250 0.0
V21000 n0_12616_11433 n2_12616_11433 0.0
V21001 n0_12616_11466 n2_12616_11466 0.0
V21002 n0_12616_11649 n2_12616_11649 0.0
V21003 n0_12616_11682 n2_12616_11682 0.0
V21004 n0_12616_11865 n2_12616_11865 0.0
V21005 n0_12616_11898 n2_12616_11898 0.0
V21006 n0_12616_11912 n2_12616_11912 0.0
V21007 n0_12616_12081 n2_12616_12081 0.0
V21008 n0_12616_12114 n2_12616_12114 0.0
V21009 n0_12616_12128 n2_12616_12128 0.0
V21010 n0_12616_12285 n2_12616_12285 0.0
V21011 n0_12616_12297 n2_12616_12297 0.0
V21012 n0_12616_12330 n2_12616_12330 0.0
V21013 n0_12616_12513 n2_12616_12513 0.0
V21014 n0_12616_12546 n2_12616_12546 0.0
V21015 n0_12616_12729 n2_12616_12729 0.0
V21016 n0_12616_12762 n2_12616_12762 0.0
V21017 n0_12616_12945 n2_12616_12945 0.0
V21018 n0_12616_12978 n2_12616_12978 0.0
V21019 n0_12616_13129 n2_12616_13129 0.0
V21020 n0_12616_13161 n2_12616_13161 0.0
V21021 n0_12616_13194 n2_12616_13194 0.0
V21022 n0_12616_13377 n2_12616_13377 0.0
V21023 n0_12616_13410 n2_12616_13410 0.0
V21024 n0_12616_13593 n2_12616_13593 0.0
V21025 n0_12616_13626 n2_12616_13626 0.0
V21026 n0_12616_13663 n2_12616_13663 0.0
V21027 n0_12616_13700 n2_12616_13700 0.0
V21028 n0_12616_13809 n2_12616_13809 0.0
V21029 n0_12616_13842 n2_12616_13842 0.0
V21030 n0_12616_14025 n2_12616_14025 0.0
V21031 n0_12616_14058 n2_12616_14058 0.0
V21032 n0_12616_14079 n2_12616_14079 0.0
V21033 n0_12616_14229 n2_12616_14229 0.0
V21034 n0_12616_14241 n2_12616_14241 0.0
V21035 n0_12616_14274 n2_12616_14274 0.0
V21036 n0_12616_14457 n2_12616_14457 0.0
V21037 n0_12616_14490 n2_12616_14490 0.0
V21038 n0_12616_14673 n2_12616_14673 0.0
V21039 n0_12616_14706 n2_12616_14706 0.0
V21040 n0_12616_14727 n2_12616_14727 0.0
V21041 n0_12616_14816 n2_12616_14816 0.0
V21042 n0_12616_14889 n2_12616_14889 0.0
V21043 n0_12616_14922 n2_12616_14922 0.0
V21044 n0_12616_15138 n2_12616_15138 0.0
V21045 n0_12616_15321 n2_12616_15321 0.0
V21046 n0_12616_15354 n2_12616_15354 0.0
V21047 n0_12616_15368 n2_12616_15368 0.0
V21048 n0_12616_15537 n2_12616_15537 0.0
V21049 n0_12616_15570 n2_12616_15570 0.0
V21050 n0_12616_15753 n2_12616_15753 0.0
V21051 n0_12616_15786 n2_12616_15786 0.0
V21052 n0_12616_15800 n2_12616_15800 0.0
V21053 n0_12616_15807 n2_12616_15807 0.0
V21054 n0_12616_15969 n2_12616_15969 0.0
V21055 n0_12616_16002 n2_12616_16002 0.0
V21056 n0_12616_16185 n2_12616_16185 0.0
V21057 n0_12616_16401 n2_12616_16401 0.0
V21058 n0_12616_16434 n2_12616_16434 0.0
V21059 n0_12616_16448 n2_12616_16448 0.0
V21060 n0_12616_16617 n2_12616_16617 0.0
V21061 n0_12616_16650 n2_12616_16650 0.0
V21062 n0_12616_16833 n2_12616_16833 0.0
V21063 n0_12616_16866 n2_12616_16866 0.0
V21064 n0_12616_17049 n2_12616_17049 0.0
V21065 n0_12616_17082 n2_12616_17082 0.0
V21066 n0_12616_17096 n2_12616_17096 0.0
V21067 n0_12616_17103 n2_12616_17103 0.0
V21068 n0_12616_17265 n2_12616_17265 0.0
V21069 n0_12616_17298 n2_12616_17298 0.0
V21070 n0_12616_17481 n2_12616_17481 0.0
V21071 n0_12616_17514 n2_12616_17514 0.0
V21072 n0_12616_17528 n2_12616_17528 0.0
V21073 n0_12616_17697 n2_12616_17697 0.0
V21074 n0_12616_17730 n2_12616_17730 0.0
V21075 n0_12616_17913 n2_12616_17913 0.0
V21076 n0_12616_17946 n2_12616_17946 0.0
V21077 n0_12616_17983 n2_12616_17983 0.0
V21078 n0_12616_18129 n2_12616_18129 0.0
V21079 n0_12616_18162 n2_12616_18162 0.0
V21080 n0_12616_18176 n2_12616_18176 0.0
V21081 n0_12616_18183 n2_12616_18183 0.0
V21082 n0_12616_18345 n2_12616_18345 0.0
V21083 n0_12616_18378 n2_12616_18378 0.0
V21084 n0_12616_18561 n2_12616_18561 0.0
V21085 n0_12616_18594 n2_12616_18594 0.0
V21086 n0_12616_18608 n2_12616_18608 0.0
V21087 n0_12616_18777 n2_12616_18777 0.0
V21088 n0_12616_18810 n2_12616_18810 0.0
V21089 n0_12616_18993 n2_12616_18993 0.0
V21090 n0_12616_19026 n2_12616_19026 0.0
V21091 n0_12616_19209 n2_12616_19209 0.0
V21092 n0_12616_19242 n2_12616_19242 0.0
V21093 n0_12616_19256 n2_12616_19256 0.0
V21094 n0_12616_19263 n2_12616_19263 0.0
V21095 n0_12616_19425 n2_12616_19425 0.0
V21096 n0_12616_19458 n2_12616_19458 0.0
V21097 n0_12616_19641 n2_12616_19641 0.0
V21098 n0_12616_19674 n2_12616_19674 0.0
V21099 n0_12616_19857 n2_12616_19857 0.0
V21100 n0_12616_19890 n2_12616_19890 0.0
V21101 n0_12616_20073 n2_12616_20073 0.0
V21102 n0_12616_20106 n2_12616_20106 0.0
V21103 n0_12616_20289 n2_12616_20289 0.0
V21104 n0_12616_20322 n2_12616_20322 0.0
V21105 n0_12616_20505 n2_12616_20505 0.0
V21106 n0_12616_20538 n2_12616_20538 0.0
V21107 n0_12616_20754 n2_12616_20754 0.0
V21108 n0_12616_20937 n2_12616_20937 0.0
V21109 n0_12616_20970 n2_12616_20970 0.0
V21110 n0_12708_201 n2_12708_201 0.0
V21111 n0_12708_234 n2_12708_234 0.0
V21112 n0_12708_417 n2_12708_417 0.0
V21113 n0_12708_450 n2_12708_450 0.0
V21114 n0_12708_633 n2_12708_633 0.0
V21115 n0_12708_666 n2_12708_666 0.0
V21116 n0_12708_849 n2_12708_849 0.0
V21117 n0_12708_882 n2_12708_882 0.0
V21118 n0_12708_1065 n2_12708_1065 0.0
V21119 n0_12708_1098 n2_12708_1098 0.0
V21120 n0_12708_1281 n2_12708_1281 0.0
V21121 n0_12708_1314 n2_12708_1314 0.0
V21122 n0_12708_1497 n2_12708_1497 0.0
V21123 n0_12708_1530 n2_12708_1530 0.0
V21124 n0_12708_1713 n2_12708_1713 0.0
V21125 n0_12708_1746 n2_12708_1746 0.0
V21126 n0_12708_1783 n2_12708_1783 0.0
V21127 n0_12708_1929 n2_12708_1929 0.0
V21128 n0_12708_1962 n2_12708_1962 0.0
V21129 n0_12708_2145 n2_12708_2145 0.0
V21130 n0_12708_2178 n2_12708_2178 0.0
V21131 n0_12708_2361 n2_12708_2361 0.0
V21132 n0_12708_2394 n2_12708_2394 0.0
V21133 n0_12708_2431 n2_12708_2431 0.0
V21134 n0_12708_2577 n2_12708_2577 0.0
V21135 n0_12708_2610 n2_12708_2610 0.0
V21136 n0_12708_2793 n2_12708_2793 0.0
V21137 n0_12708_2826 n2_12708_2826 0.0
V21138 n0_12708_2863 n2_12708_2863 0.0
V21139 n0_12708_3009 n2_12708_3009 0.0
V21140 n0_12708_3042 n2_12708_3042 0.0
V21141 n0_12708_3225 n2_12708_3225 0.0
V21142 n0_12708_3258 n2_12708_3258 0.0
V21143 n0_12708_3441 n2_12708_3441 0.0
V21144 n0_12708_3474 n2_12708_3474 0.0
V21145 n0_12708_3511 n2_12708_3511 0.0
V21146 n0_12708_3657 n2_12708_3657 0.0
V21147 n0_12708_3690 n2_12708_3690 0.0
V21148 n0_12708_3873 n2_12708_3873 0.0
V21149 n0_12708_3906 n2_12708_3906 0.0
V21150 n0_12708_3943 n2_12708_3943 0.0
V21151 n0_12708_4089 n2_12708_4089 0.0
V21152 n0_12708_4122 n2_12708_4122 0.0
V21153 n0_12708_4159 n2_12708_4159 0.0
V21154 n0_12708_4305 n2_12708_4305 0.0
V21155 n0_12708_4338 n2_12708_4338 0.0
V21156 n0_12708_4521 n2_12708_4521 0.0
V21157 n0_12708_4554 n2_12708_4554 0.0
V21158 n0_12708_4591 n2_12708_4591 0.0
V21159 n0_12708_4737 n2_12708_4737 0.0
V21160 n0_12708_4770 n2_12708_4770 0.0
V21161 n0_12708_4953 n2_12708_4953 0.0
V21162 n0_12708_4986 n2_12708_4986 0.0
V21163 n0_12708_5023 n2_12708_5023 0.0
V21164 n0_12708_5169 n2_12708_5169 0.0
V21165 n0_12708_5202 n2_12708_5202 0.0
V21166 n0_12708_5239 n2_12708_5239 0.0
V21167 n0_12708_5385 n2_12708_5385 0.0
V21168 n0_12708_5418 n2_12708_5418 0.0
V21169 n0_12708_5601 n2_12708_5601 0.0
V21170 n0_12708_5634 n2_12708_5634 0.0
V21171 n0_12708_5671 n2_12708_5671 0.0
V21172 n0_12708_5817 n2_12708_5817 0.0
V21173 n0_12708_5850 n2_12708_5850 0.0
V21174 n0_12708_6033 n2_12708_6033 0.0
V21175 n0_12708_6066 n2_12708_6066 0.0
V21176 n0_12708_6249 n2_12708_6249 0.0
V21177 n0_12708_6282 n2_12708_6282 0.0
V21178 n0_12708_6319 n2_12708_6319 0.0
V21179 n0_12708_6465 n2_12708_6465 0.0
V21180 n0_12708_6498 n2_12708_6498 0.0
V21181 n0_12708_6681 n2_12708_6681 0.0
V21182 n0_12708_6714 n2_12708_6714 0.0
V21183 n0_12708_6751 n2_12708_6751 0.0
V21184 n0_12708_6897 n2_12708_6897 0.0
V21185 n0_12708_6930 n2_12708_6930 0.0
V21186 n0_12708_6967 n2_12708_6967 0.0
V21187 n0_12708_7113 n2_12708_7113 0.0
V21188 n0_12708_7146 n2_12708_7146 0.0
V21189 n0_12708_7178 n2_12708_7178 0.0
V21190 n0_12708_7329 n2_12708_7329 0.0
V21191 n0_12708_7362 n2_12708_7362 0.0
V21192 n0_12708_7399 n2_12708_7399 0.0
V21193 n0_12708_7545 n2_12708_7545 0.0
V21194 n0_12708_7578 n2_12708_7578 0.0
V21195 n0_12708_7761 n2_12708_7761 0.0
V21196 n0_12708_7794 n2_12708_7794 0.0
V21197 n0_12708_7831 n2_12708_7831 0.0
V21198 n0_12708_7977 n2_12708_7977 0.0
V21199 n0_12708_8010 n2_12708_8010 0.0
V21200 n0_12708_8193 n2_12708_8193 0.0
V21201 n0_12708_8226 n2_12708_8226 0.0
V21202 n0_12708_8409 n2_12708_8409 0.0
V21203 n0_12708_8442 n2_12708_8442 0.0
V21204 n0_12708_12762 n2_12708_12762 0.0
V21205 n0_12708_12945 n2_12708_12945 0.0
V21206 n0_12708_12978 n2_12708_12978 0.0
V21207 n0_12708_13161 n2_12708_13161 0.0
V21208 n0_12708_13194 n2_12708_13194 0.0
V21209 n0_12708_13377 n2_12708_13377 0.0
V21210 n0_12708_13410 n2_12708_13410 0.0
V21211 n0_12708_13593 n2_12708_13593 0.0
V21212 n0_12708_13626 n2_12708_13626 0.0
V21213 n0_12708_13663 n2_12708_13663 0.0
V21214 n0_12708_13809 n2_12708_13809 0.0
V21215 n0_12708_13842 n2_12708_13842 0.0
V21216 n0_12708_14025 n2_12708_14025 0.0
V21217 n0_12708_14058 n2_12708_14058 0.0
V21218 n0_12708_14079 n2_12708_14079 0.0
V21219 n0_12708_14241 n2_12708_14241 0.0
V21220 n0_12708_14274 n2_12708_14274 0.0
V21221 n0_12708_14457 n2_12708_14457 0.0
V21222 n0_12708_14490 n2_12708_14490 0.0
V21223 n0_12708_14673 n2_12708_14673 0.0
V21224 n0_12708_14706 n2_12708_14706 0.0
V21225 n0_12708_14727 n2_12708_14727 0.0
V21226 n0_12708_14889 n2_12708_14889 0.0
V21227 n0_12708_14922 n2_12708_14922 0.0
V21228 n0_12708_15105 n2_12708_15105 0.0
V21229 n0_12708_15138 n2_12708_15138 0.0
V21230 n0_12708_15321 n2_12708_15321 0.0
V21231 n0_12708_15354 n2_12708_15354 0.0
V21232 n0_12708_15368 n2_12708_15368 0.0
V21233 n0_12708_15537 n2_12708_15537 0.0
V21234 n0_12708_15570 n2_12708_15570 0.0
V21235 n0_12708_15753 n2_12708_15753 0.0
V21236 n0_12708_15786 n2_12708_15786 0.0
V21237 n0_12708_15800 n2_12708_15800 0.0
V21238 n0_12708_15807 n2_12708_15807 0.0
V21239 n0_12708_15969 n2_12708_15969 0.0
V21240 n0_12708_16002 n2_12708_16002 0.0
V21241 n0_12708_16185 n2_12708_16185 0.0
V21242 n0_12708_16218 n2_12708_16218 0.0
V21243 n0_12708_16401 n2_12708_16401 0.0
V21244 n0_12708_16434 n2_12708_16434 0.0
V21245 n0_12708_16448 n2_12708_16448 0.0
V21246 n0_12708_16617 n2_12708_16617 0.0
V21247 n0_12708_16650 n2_12708_16650 0.0
V21248 n0_12708_16833 n2_12708_16833 0.0
V21249 n0_12708_16866 n2_12708_16866 0.0
V21250 n0_12708_17049 n2_12708_17049 0.0
V21251 n0_12708_17082 n2_12708_17082 0.0
V21252 n0_12708_17096 n2_12708_17096 0.0
V21253 n0_12708_17103 n2_12708_17103 0.0
V21254 n0_12708_17265 n2_12708_17265 0.0
V21255 n0_12708_17298 n2_12708_17298 0.0
V21256 n0_12708_17481 n2_12708_17481 0.0
V21257 n0_12708_17514 n2_12708_17514 0.0
V21258 n0_12708_17528 n2_12708_17528 0.0
V21259 n0_12708_17697 n2_12708_17697 0.0
V21260 n0_12708_17730 n2_12708_17730 0.0
V21261 n0_12708_17913 n2_12708_17913 0.0
V21262 n0_12708_17946 n2_12708_17946 0.0
V21263 n0_12708_17983 n2_12708_17983 0.0
V21264 n0_12708_18129 n2_12708_18129 0.0
V21265 n0_12708_18162 n2_12708_18162 0.0
V21266 n0_12708_18176 n2_12708_18176 0.0
V21267 n0_12708_18183 n2_12708_18183 0.0
V21268 n0_12708_18345 n2_12708_18345 0.0
V21269 n0_12708_18378 n2_12708_18378 0.0
V21270 n0_12708_18561 n2_12708_18561 0.0
V21271 n0_12708_18594 n2_12708_18594 0.0
V21272 n0_12708_18608 n2_12708_18608 0.0
V21273 n0_12708_18777 n2_12708_18777 0.0
V21274 n0_12708_18810 n2_12708_18810 0.0
V21275 n0_12708_18993 n2_12708_18993 0.0
V21276 n0_12708_19026 n2_12708_19026 0.0
V21277 n0_12708_19209 n2_12708_19209 0.0
V21278 n0_12708_19242 n2_12708_19242 0.0
V21279 n0_12708_19256 n2_12708_19256 0.0
V21280 n0_12708_19263 n2_12708_19263 0.0
V21281 n0_12708_19425 n2_12708_19425 0.0
V21282 n0_12708_19458 n2_12708_19458 0.0
V21283 n0_12708_19641 n2_12708_19641 0.0
V21284 n0_12708_19674 n2_12708_19674 0.0
V21285 n0_12708_19857 n2_12708_19857 0.0
V21286 n0_12708_19890 n2_12708_19890 0.0
V21287 n0_12708_20073 n2_12708_20073 0.0
V21288 n0_12708_20106 n2_12708_20106 0.0
V21289 n0_12708_20289 n2_12708_20289 0.0
V21290 n0_12708_20322 n2_12708_20322 0.0
V21291 n0_12708_20505 n2_12708_20505 0.0
V21292 n0_12708_20538 n2_12708_20538 0.0
V21293 n0_12708_20721 n2_12708_20721 0.0
V21294 n0_12708_20754 n2_12708_20754 0.0
V21295 n0_12708_20937 n2_12708_20937 0.0
V21296 n0_12708_20970 n2_12708_20970 0.0
V21297 n0_12755_417 n2_12755_417 0.0
V21298 n0_12755_450 n2_12755_450 0.0
V21299 n0_12755_1530 n2_12755_1530 0.0
V21300 n0_12755_2793 n2_12755_2793 0.0
V21301 n0_12755_3873 n2_12755_3873 0.0
V21302 n0_12755_3906 n2_12755_3906 0.0
V21303 n0_12755_4953 n2_12755_4953 0.0
V21304 n0_12755_4986 n2_12755_4986 0.0
V21305 n0_12755_5023 n2_12755_5023 0.0
V21306 n0_12755_6033 n2_12755_6033 0.0
V21307 n0_12755_6066 n2_12755_6066 0.0
V21308 n0_12755_7146 n2_12755_7146 0.0
V21309 n0_12755_7178 n2_12755_7178 0.0
V21310 n0_12755_8409 n2_12755_8409 0.0
V21311 n0_12755_10569 n2_12755_10569 0.0
V21312 n0_12755_10602 n2_12755_10602 0.0
V21313 n0_12755_14025 n2_12755_14025 0.0
V21314 n0_12755_15105 n2_12755_15105 0.0
V21315 n0_12755_15138 n2_12755_15138 0.0
V21316 n0_12755_16185 n2_12755_16185 0.0
V21317 n0_12755_16218 n2_12755_16218 0.0
V21318 n0_12755_17298 n2_12755_17298 0.0
V21319 n0_12755_19641 n2_12755_19641 0.0
V21320 n0_12755_19674 n2_12755_19674 0.0
V21321 n0_12755_20721 n2_12755_20721 0.0
V21322 n0_12755_20754 n2_12755_20754 0.0
V21323 n0_12804_201 n2_12804_201 0.0
V21324 n0_12804_234 n2_12804_234 0.0
V21325 n0_12804_417 n2_12804_417 0.0
V21326 n0_12804_450 n2_12804_450 0.0
V21327 n0_12804_633 n2_12804_633 0.0
V21328 n0_12804_666 n2_12804_666 0.0
V21329 n0_12804_849 n2_12804_849 0.0
V21330 n0_12804_882 n2_12804_882 0.0
V21331 n0_12804_1065 n2_12804_1065 0.0
V21332 n0_12804_1098 n2_12804_1098 0.0
V21333 n0_12804_1281 n2_12804_1281 0.0
V21334 n0_12804_1314 n2_12804_1314 0.0
V21335 n0_12804_1497 n2_12804_1497 0.0
V21336 n0_12804_1530 n2_12804_1530 0.0
V21337 n0_12804_1713 n2_12804_1713 0.0
V21338 n0_12804_1746 n2_12804_1746 0.0
V21339 n0_12804_1783 n2_12804_1783 0.0
V21340 n0_12804_1929 n2_12804_1929 0.0
V21341 n0_12804_1962 n2_12804_1962 0.0
V21342 n0_12804_2145 n2_12804_2145 0.0
V21343 n0_12804_2178 n2_12804_2178 0.0
V21344 n0_12804_2361 n2_12804_2361 0.0
V21345 n0_12804_2394 n2_12804_2394 0.0
V21346 n0_12804_2431 n2_12804_2431 0.0
V21347 n0_12804_2577 n2_12804_2577 0.0
V21348 n0_12804_2610 n2_12804_2610 0.0
V21349 n0_12804_2793 n2_12804_2793 0.0
V21350 n0_12804_2826 n2_12804_2826 0.0
V21351 n0_12804_2863 n2_12804_2863 0.0
V21352 n0_12804_3009 n2_12804_3009 0.0
V21353 n0_12804_3042 n2_12804_3042 0.0
V21354 n0_12804_3225 n2_12804_3225 0.0
V21355 n0_12804_3258 n2_12804_3258 0.0
V21356 n0_12804_3441 n2_12804_3441 0.0
V21357 n0_12804_3474 n2_12804_3474 0.0
V21358 n0_12804_3511 n2_12804_3511 0.0
V21359 n0_12804_3657 n2_12804_3657 0.0
V21360 n0_12804_3690 n2_12804_3690 0.0
V21361 n0_12804_3873 n2_12804_3873 0.0
V21362 n0_12804_3906 n2_12804_3906 0.0
V21363 n0_12804_3943 n2_12804_3943 0.0
V21364 n0_12804_4089 n2_12804_4089 0.0
V21365 n0_12804_4122 n2_12804_4122 0.0
V21366 n0_12804_4159 n2_12804_4159 0.0
V21367 n0_12804_4305 n2_12804_4305 0.0
V21368 n0_12804_4338 n2_12804_4338 0.0
V21369 n0_12804_4521 n2_12804_4521 0.0
V21370 n0_12804_4554 n2_12804_4554 0.0
V21371 n0_12804_4591 n2_12804_4591 0.0
V21372 n0_12804_4737 n2_12804_4737 0.0
V21373 n0_12804_4770 n2_12804_4770 0.0
V21374 n0_12804_4953 n2_12804_4953 0.0
V21375 n0_12804_4986 n2_12804_4986 0.0
V21376 n0_12804_5023 n2_12804_5023 0.0
V21377 n0_12804_5169 n2_12804_5169 0.0
V21378 n0_12804_5202 n2_12804_5202 0.0
V21379 n0_12804_5239 n2_12804_5239 0.0
V21380 n0_12804_5385 n2_12804_5385 0.0
V21381 n0_12804_5418 n2_12804_5418 0.0
V21382 n0_12804_5601 n2_12804_5601 0.0
V21383 n0_12804_5634 n2_12804_5634 0.0
V21384 n0_12804_5671 n2_12804_5671 0.0
V21385 n0_12804_5817 n2_12804_5817 0.0
V21386 n0_12804_5850 n2_12804_5850 0.0
V21387 n0_12804_6033 n2_12804_6033 0.0
V21388 n0_12804_6066 n2_12804_6066 0.0
V21389 n0_12804_6249 n2_12804_6249 0.0
V21390 n0_12804_6282 n2_12804_6282 0.0
V21391 n0_12804_6319 n2_12804_6319 0.0
V21392 n0_12804_6465 n2_12804_6465 0.0
V21393 n0_12804_6498 n2_12804_6498 0.0
V21394 n0_12804_6681 n2_12804_6681 0.0
V21395 n0_12804_6714 n2_12804_6714 0.0
V21396 n0_12804_6751 n2_12804_6751 0.0
V21397 n0_12804_6897 n2_12804_6897 0.0
V21398 n0_12804_6930 n2_12804_6930 0.0
V21399 n0_12804_6967 n2_12804_6967 0.0
V21400 n0_12804_7113 n2_12804_7113 0.0
V21401 n0_12804_7146 n2_12804_7146 0.0
V21402 n0_12804_7178 n2_12804_7178 0.0
V21403 n0_12804_7329 n2_12804_7329 0.0
V21404 n0_12804_7362 n2_12804_7362 0.0
V21405 n0_12804_7399 n2_12804_7399 0.0
V21406 n0_12804_7545 n2_12804_7545 0.0
V21407 n0_12804_7578 n2_12804_7578 0.0
V21408 n0_12804_7761 n2_12804_7761 0.0
V21409 n0_12804_7794 n2_12804_7794 0.0
V21410 n0_12804_7831 n2_12804_7831 0.0
V21411 n0_12804_7977 n2_12804_7977 0.0
V21412 n0_12804_8010 n2_12804_8010 0.0
V21413 n0_12804_8193 n2_12804_8193 0.0
V21414 n0_12804_8226 n2_12804_8226 0.0
V21415 n0_12804_8409 n2_12804_8409 0.0
V21416 n0_12804_8442 n2_12804_8442 0.0
V21417 n0_12804_8625 n2_12804_8625 0.0
V21418 n0_12804_8658 n2_12804_8658 0.0
V21419 n0_12804_8695 n2_12804_8695 0.0
V21420 n0_12804_8841 n2_12804_8841 0.0
V21421 n0_12804_8874 n2_12804_8874 0.0
V21422 n0_12804_8911 n2_12804_8911 0.0
V21423 n0_12804_9057 n2_12804_9057 0.0
V21424 n0_12804_9090 n2_12804_9090 0.0
V21425 n0_12804_9273 n2_12804_9273 0.0
V21426 n0_12804_9306 n2_12804_9306 0.0
V21427 n0_12804_9705 n2_12804_9705 0.0
V21428 n0_12804_9738 n2_12804_9738 0.0
V21429 n0_12804_9775 n2_12804_9775 0.0
V21430 n0_12804_9921 n2_12804_9921 0.0
V21431 n0_12804_9954 n2_12804_9954 0.0
V21432 n0_12804_9991 n2_12804_9991 0.0
V21433 n0_12804_10137 n2_12804_10137 0.0
V21434 n0_12804_10170 n2_12804_10170 0.0
V21435 n0_12804_10353 n2_12804_10353 0.0
V21436 n0_12804_10386 n2_12804_10386 0.0
V21437 n0_12804_10569 n2_12804_10569 0.0
V21438 n0_12804_10602 n2_12804_10602 0.0
V21439 n0_12804_10785 n2_12804_10785 0.0
V21440 n0_12804_10818 n2_12804_10818 0.0
V21441 n0_12804_10832 n2_12804_10832 0.0
V21442 n0_12804_11001 n2_12804_11001 0.0
V21443 n0_12804_11034 n2_12804_11034 0.0
V21444 n0_12804_11048 n2_12804_11048 0.0
V21445 n0_12804_11217 n2_12804_11217 0.0
V21446 n0_12804_11250 n2_12804_11250 0.0
V21447 n0_12804_11433 n2_12804_11433 0.0
V21448 n0_12804_11466 n2_12804_11466 0.0
V21449 n0_12804_11865 n2_12804_11865 0.0
V21450 n0_12804_11898 n2_12804_11898 0.0
V21451 n0_12804_11912 n2_12804_11912 0.0
V21452 n0_12804_12081 n2_12804_12081 0.0
V21453 n0_12804_12114 n2_12804_12114 0.0
V21454 n0_12804_12128 n2_12804_12128 0.0
V21455 n0_12804_12297 n2_12804_12297 0.0
V21456 n0_12804_12330 n2_12804_12330 0.0
V21457 n0_12804_12513 n2_12804_12513 0.0
V21458 n0_12804_12546 n2_12804_12546 0.0
V21459 n0_12804_12729 n2_12804_12729 0.0
V21460 n0_12804_12762 n2_12804_12762 0.0
V21461 n0_12804_12945 n2_12804_12945 0.0
V21462 n0_12804_12978 n2_12804_12978 0.0
V21463 n0_12804_13161 n2_12804_13161 0.0
V21464 n0_12804_13194 n2_12804_13194 0.0
V21465 n0_12804_13377 n2_12804_13377 0.0
V21466 n0_12804_13410 n2_12804_13410 0.0
V21467 n0_12804_13593 n2_12804_13593 0.0
V21468 n0_12804_13626 n2_12804_13626 0.0
V21469 n0_12804_13663 n2_12804_13663 0.0
V21470 n0_12804_13809 n2_12804_13809 0.0
V21471 n0_12804_13842 n2_12804_13842 0.0
V21472 n0_12804_14025 n2_12804_14025 0.0
V21473 n0_12804_14058 n2_12804_14058 0.0
V21474 n0_12804_14079 n2_12804_14079 0.0
V21475 n0_12804_14241 n2_12804_14241 0.0
V21476 n0_12804_14274 n2_12804_14274 0.0
V21477 n0_12804_14457 n2_12804_14457 0.0
V21478 n0_12804_14490 n2_12804_14490 0.0
V21479 n0_12804_14673 n2_12804_14673 0.0
V21480 n0_12804_14706 n2_12804_14706 0.0
V21481 n0_12804_14727 n2_12804_14727 0.0
V21482 n0_12804_14889 n2_12804_14889 0.0
V21483 n0_12804_14922 n2_12804_14922 0.0
V21484 n0_12804_15105 n2_12804_15105 0.0
V21485 n0_12804_15138 n2_12804_15138 0.0
V21486 n0_12804_15321 n2_12804_15321 0.0
V21487 n0_12804_15354 n2_12804_15354 0.0
V21488 n0_12804_15368 n2_12804_15368 0.0
V21489 n0_12804_15537 n2_12804_15537 0.0
V21490 n0_12804_15570 n2_12804_15570 0.0
V21491 n0_12804_15753 n2_12804_15753 0.0
V21492 n0_12804_15786 n2_12804_15786 0.0
V21493 n0_12804_15800 n2_12804_15800 0.0
V21494 n0_12804_15807 n2_12804_15807 0.0
V21495 n0_12804_15969 n2_12804_15969 0.0
V21496 n0_12804_16002 n2_12804_16002 0.0
V21497 n0_12804_16185 n2_12804_16185 0.0
V21498 n0_12804_16218 n2_12804_16218 0.0
V21499 n0_12804_16401 n2_12804_16401 0.0
V21500 n0_12804_16434 n2_12804_16434 0.0
V21501 n0_12804_16448 n2_12804_16448 0.0
V21502 n0_12804_16617 n2_12804_16617 0.0
V21503 n0_12804_16650 n2_12804_16650 0.0
V21504 n0_12804_16833 n2_12804_16833 0.0
V21505 n0_12804_16866 n2_12804_16866 0.0
V21506 n0_12804_17049 n2_12804_17049 0.0
V21507 n0_12804_17082 n2_12804_17082 0.0
V21508 n0_12804_17096 n2_12804_17096 0.0
V21509 n0_12804_17103 n2_12804_17103 0.0
V21510 n0_12804_17265 n2_12804_17265 0.0
V21511 n0_12804_17298 n2_12804_17298 0.0
V21512 n0_12804_17481 n2_12804_17481 0.0
V21513 n0_12804_17514 n2_12804_17514 0.0
V21514 n0_12804_17528 n2_12804_17528 0.0
V21515 n0_12804_17697 n2_12804_17697 0.0
V21516 n0_12804_17730 n2_12804_17730 0.0
V21517 n0_12804_17913 n2_12804_17913 0.0
V21518 n0_12804_17946 n2_12804_17946 0.0
V21519 n0_12804_17983 n2_12804_17983 0.0
V21520 n0_12804_18129 n2_12804_18129 0.0
V21521 n0_12804_18162 n2_12804_18162 0.0
V21522 n0_12804_18176 n2_12804_18176 0.0
V21523 n0_12804_18183 n2_12804_18183 0.0
V21524 n0_12804_18345 n2_12804_18345 0.0
V21525 n0_12804_18378 n2_12804_18378 0.0
V21526 n0_12804_18561 n2_12804_18561 0.0
V21527 n0_12804_18594 n2_12804_18594 0.0
V21528 n0_12804_18608 n2_12804_18608 0.0
V21529 n0_12804_18777 n2_12804_18777 0.0
V21530 n0_12804_18810 n2_12804_18810 0.0
V21531 n0_12804_18993 n2_12804_18993 0.0
V21532 n0_12804_19026 n2_12804_19026 0.0
V21533 n0_12804_19209 n2_12804_19209 0.0
V21534 n0_12804_19242 n2_12804_19242 0.0
V21535 n0_12804_19256 n2_12804_19256 0.0
V21536 n0_12804_19263 n2_12804_19263 0.0
V21537 n0_12804_19425 n2_12804_19425 0.0
V21538 n0_12804_19458 n2_12804_19458 0.0
V21539 n0_12804_19641 n2_12804_19641 0.0
V21540 n0_12804_19674 n2_12804_19674 0.0
V21541 n0_12804_19857 n2_12804_19857 0.0
V21542 n0_12804_19890 n2_12804_19890 0.0
V21543 n0_12804_20073 n2_12804_20073 0.0
V21544 n0_12804_20106 n2_12804_20106 0.0
V21545 n0_12804_20289 n2_12804_20289 0.0
V21546 n0_12804_20322 n2_12804_20322 0.0
V21547 n0_12804_20505 n2_12804_20505 0.0
V21548 n0_12804_20538 n2_12804_20538 0.0
V21549 n0_12804_20721 n2_12804_20721 0.0
V21550 n0_12804_20754 n2_12804_20754 0.0
V21551 n0_12804_20937 n2_12804_20937 0.0
V21552 n0_12804_20970 n2_12804_20970 0.0
V21553 n0_12896_201 n2_12896_201 0.0
V21554 n0_12896_234 n2_12896_234 0.0
V21555 n0_12896_417 n2_12896_417 0.0
V21556 n0_12896_450 n2_12896_450 0.0
V21557 n0_12896_633 n2_12896_633 0.0
V21558 n0_12896_666 n2_12896_666 0.0
V21559 n0_12896_849 n2_12896_849 0.0
V21560 n0_12896_882 n2_12896_882 0.0
V21561 n0_12896_1065 n2_12896_1065 0.0
V21562 n0_12896_1098 n2_12896_1098 0.0
V21563 n0_12896_1281 n2_12896_1281 0.0
V21564 n0_12896_1314 n2_12896_1314 0.0
V21565 n0_12896_1497 n2_12896_1497 0.0
V21566 n0_12896_1530 n2_12896_1530 0.0
V21567 n0_12896_1713 n2_12896_1713 0.0
V21568 n0_12896_1746 n2_12896_1746 0.0
V21569 n0_12896_1783 n2_12896_1783 0.0
V21570 n0_12896_1929 n2_12896_1929 0.0
V21571 n0_12896_1962 n2_12896_1962 0.0
V21572 n0_12896_2145 n2_12896_2145 0.0
V21573 n0_12896_2178 n2_12896_2178 0.0
V21574 n0_12896_2361 n2_12896_2361 0.0
V21575 n0_12896_2394 n2_12896_2394 0.0
V21576 n0_12896_2431 n2_12896_2431 0.0
V21577 n0_12896_2577 n2_12896_2577 0.0
V21578 n0_12896_2610 n2_12896_2610 0.0
V21579 n0_12896_2793 n2_12896_2793 0.0
V21580 n0_12896_2826 n2_12896_2826 0.0
V21581 n0_12896_2863 n2_12896_2863 0.0
V21582 n0_12896_3009 n2_12896_3009 0.0
V21583 n0_12896_3042 n2_12896_3042 0.0
V21584 n0_12896_3225 n2_12896_3225 0.0
V21585 n0_12896_3258 n2_12896_3258 0.0
V21586 n0_12896_3441 n2_12896_3441 0.0
V21587 n0_12896_3474 n2_12896_3474 0.0
V21588 n0_12896_3511 n2_12896_3511 0.0
V21589 n0_12896_3657 n2_12896_3657 0.0
V21590 n0_12896_3690 n2_12896_3690 0.0
V21591 n0_12896_3873 n2_12896_3873 0.0
V21592 n0_12896_3906 n2_12896_3906 0.0
V21593 n0_12896_3943 n2_12896_3943 0.0
V21594 n0_12896_4089 n2_12896_4089 0.0
V21595 n0_12896_4122 n2_12896_4122 0.0
V21596 n0_12896_4159 n2_12896_4159 0.0
V21597 n0_12896_4305 n2_12896_4305 0.0
V21598 n0_12896_4338 n2_12896_4338 0.0
V21599 n0_12896_4521 n2_12896_4521 0.0
V21600 n0_12896_4554 n2_12896_4554 0.0
V21601 n0_12896_4591 n2_12896_4591 0.0
V21602 n0_12896_4737 n2_12896_4737 0.0
V21603 n0_12896_4770 n2_12896_4770 0.0
V21604 n0_12896_4953 n2_12896_4953 0.0
V21605 n0_12896_5023 n2_12896_5023 0.0
V21606 n0_12896_5169 n2_12896_5169 0.0
V21607 n0_12896_5202 n2_12896_5202 0.0
V21608 n0_12896_5239 n2_12896_5239 0.0
V21609 n0_12896_5385 n2_12896_5385 0.0
V21610 n0_12896_5418 n2_12896_5418 0.0
V21611 n0_12896_5601 n2_12896_5601 0.0
V21612 n0_12896_5634 n2_12896_5634 0.0
V21613 n0_12896_5671 n2_12896_5671 0.0
V21614 n0_12896_5817 n2_12896_5817 0.0
V21615 n0_12896_5850 n2_12896_5850 0.0
V21616 n0_12896_6033 n2_12896_6033 0.0
V21617 n0_12896_6066 n2_12896_6066 0.0
V21618 n0_12896_6249 n2_12896_6249 0.0
V21619 n0_12896_6282 n2_12896_6282 0.0
V21620 n0_12896_6319 n2_12896_6319 0.0
V21621 n0_12896_6465 n2_12896_6465 0.0
V21622 n0_12896_6498 n2_12896_6498 0.0
V21623 n0_12896_6681 n2_12896_6681 0.0
V21624 n0_12896_6714 n2_12896_6714 0.0
V21625 n0_12896_6751 n2_12896_6751 0.0
V21626 n0_12896_6897 n2_12896_6897 0.0
V21627 n0_12896_6930 n2_12896_6930 0.0
V21628 n0_12896_6967 n2_12896_6967 0.0
V21629 n0_12896_7113 n2_12896_7113 0.0
V21630 n0_12896_7146 n2_12896_7146 0.0
V21631 n0_12896_7178 n2_12896_7178 0.0
V21632 n0_12896_7329 n2_12896_7329 0.0
V21633 n0_12896_7362 n2_12896_7362 0.0
V21634 n0_12896_7399 n2_12896_7399 0.0
V21635 n0_12896_7545 n2_12896_7545 0.0
V21636 n0_12896_7578 n2_12896_7578 0.0
V21637 n0_12896_7761 n2_12896_7761 0.0
V21638 n0_12896_7794 n2_12896_7794 0.0
V21639 n0_12896_7831 n2_12896_7831 0.0
V21640 n0_12896_7977 n2_12896_7977 0.0
V21641 n0_12896_8010 n2_12896_8010 0.0
V21642 n0_12896_8193 n2_12896_8193 0.0
V21643 n0_12896_8226 n2_12896_8226 0.0
V21644 n0_12896_12945 n2_12896_12945 0.0
V21645 n0_12896_12978 n2_12896_12978 0.0
V21646 n0_12896_13161 n2_12896_13161 0.0
V21647 n0_12896_13194 n2_12896_13194 0.0
V21648 n0_12896_13377 n2_12896_13377 0.0
V21649 n0_12896_13410 n2_12896_13410 0.0
V21650 n0_12896_13593 n2_12896_13593 0.0
V21651 n0_12896_13626 n2_12896_13626 0.0
V21652 n0_12896_13663 n2_12896_13663 0.0
V21653 n0_12896_13809 n2_12896_13809 0.0
V21654 n0_12896_13842 n2_12896_13842 0.0
V21655 n0_12896_14025 n2_12896_14025 0.0
V21656 n0_12896_14058 n2_12896_14058 0.0
V21657 n0_12896_14079 n2_12896_14079 0.0
V21658 n0_12896_14241 n2_12896_14241 0.0
V21659 n0_12896_14274 n2_12896_14274 0.0
V21660 n0_12896_14457 n2_12896_14457 0.0
V21661 n0_12896_14490 n2_12896_14490 0.0
V21662 n0_12896_14673 n2_12896_14673 0.0
V21663 n0_12896_14706 n2_12896_14706 0.0
V21664 n0_12896_14727 n2_12896_14727 0.0
V21665 n0_12896_14889 n2_12896_14889 0.0
V21666 n0_12896_14922 n2_12896_14922 0.0
V21667 n0_12896_15138 n2_12896_15138 0.0
V21668 n0_12896_15321 n2_12896_15321 0.0
V21669 n0_12896_15354 n2_12896_15354 0.0
V21670 n0_12896_15368 n2_12896_15368 0.0
V21671 n0_12896_15537 n2_12896_15537 0.0
V21672 n0_12896_15570 n2_12896_15570 0.0
V21673 n0_12896_15753 n2_12896_15753 0.0
V21674 n0_12896_15786 n2_12896_15786 0.0
V21675 n0_12896_15800 n2_12896_15800 0.0
V21676 n0_12896_15807 n2_12896_15807 0.0
V21677 n0_12896_15969 n2_12896_15969 0.0
V21678 n0_12896_16002 n2_12896_16002 0.0
V21679 n0_12896_16185 n2_12896_16185 0.0
V21680 n0_12896_16401 n2_12896_16401 0.0
V21681 n0_12896_16434 n2_12896_16434 0.0
V21682 n0_12896_16448 n2_12896_16448 0.0
V21683 n0_12896_16617 n2_12896_16617 0.0
V21684 n0_12896_16650 n2_12896_16650 0.0
V21685 n0_12896_16833 n2_12896_16833 0.0
V21686 n0_12896_16866 n2_12896_16866 0.0
V21687 n0_12896_17049 n2_12896_17049 0.0
V21688 n0_12896_17082 n2_12896_17082 0.0
V21689 n0_12896_17096 n2_12896_17096 0.0
V21690 n0_12896_17103 n2_12896_17103 0.0
V21691 n0_12896_17265 n2_12896_17265 0.0
V21692 n0_12896_17298 n2_12896_17298 0.0
V21693 n0_12896_17481 n2_12896_17481 0.0
V21694 n0_12896_17514 n2_12896_17514 0.0
V21695 n0_12896_17528 n2_12896_17528 0.0
V21696 n0_12896_17697 n2_12896_17697 0.0
V21697 n0_12896_17730 n2_12896_17730 0.0
V21698 n0_12896_17913 n2_12896_17913 0.0
V21699 n0_12896_17946 n2_12896_17946 0.0
V21700 n0_12896_17983 n2_12896_17983 0.0
V21701 n0_12896_18129 n2_12896_18129 0.0
V21702 n0_12896_18162 n2_12896_18162 0.0
V21703 n0_12896_18176 n2_12896_18176 0.0
V21704 n0_12896_18183 n2_12896_18183 0.0
V21705 n0_12896_18345 n2_12896_18345 0.0
V21706 n0_12896_18378 n2_12896_18378 0.0
V21707 n0_12896_18561 n2_12896_18561 0.0
V21708 n0_12896_18594 n2_12896_18594 0.0
V21709 n0_12896_18608 n2_12896_18608 0.0
V21710 n0_12896_18777 n2_12896_18777 0.0
V21711 n0_12896_18810 n2_12896_18810 0.0
V21712 n0_12896_18993 n2_12896_18993 0.0
V21713 n0_12896_19026 n2_12896_19026 0.0
V21714 n0_12896_19209 n2_12896_19209 0.0
V21715 n0_12896_19242 n2_12896_19242 0.0
V21716 n0_12896_19256 n2_12896_19256 0.0
V21717 n0_12896_19263 n2_12896_19263 0.0
V21718 n0_12896_19425 n2_12896_19425 0.0
V21719 n0_12896_19458 n2_12896_19458 0.0
V21720 n0_12896_19641 n2_12896_19641 0.0
V21721 n0_12896_19674 n2_12896_19674 0.0
V21722 n0_12896_19857 n2_12896_19857 0.0
V21723 n0_12896_19890 n2_12896_19890 0.0
V21724 n0_12896_20073 n2_12896_20073 0.0
V21725 n0_12896_20106 n2_12896_20106 0.0
V21726 n0_12896_20289 n2_12896_20289 0.0
V21727 n0_12896_20322 n2_12896_20322 0.0
V21728 n0_12896_20505 n2_12896_20505 0.0
V21729 n0_12896_20538 n2_12896_20538 0.0
V21730 n0_12896_20754 n2_12896_20754 0.0
V21731 n0_12896_20937 n2_12896_20937 0.0
V21732 n0_12896_20970 n2_12896_20970 0.0
V21733 n0_13741_7329 n2_13741_7329 0.0
V21734 n0_13741_7362 n2_13741_7362 0.0
V21735 n0_13741_7545 n2_13741_7545 0.0
V21736 n0_13741_7578 n2_13741_7578 0.0
V21737 n0_13741_7761 n2_13741_7761 0.0
V21738 n0_13741_7794 n2_13741_7794 0.0
V21739 n0_13741_7831 n2_13741_7831 0.0
V21740 n0_13741_7977 n2_13741_7977 0.0
V21741 n0_13741_8010 n2_13741_8010 0.0
V21742 n0_13741_8193 n2_13741_8193 0.0
V21743 n0_13741_8226 n2_13741_8226 0.0
V21744 n0_13741_8409 n2_13741_8409 0.0
V21745 n0_13741_8442 n2_13741_8442 0.0
V21746 n0_13741_8625 n2_13741_8625 0.0
V21747 n0_13741_8658 n2_13741_8658 0.0
V21748 n0_13741_8695 n2_13741_8695 0.0
V21749 n0_13741_8841 n2_13741_8841 0.0
V21750 n0_13741_8874 n2_13741_8874 0.0
V21751 n0_13741_8911 n2_13741_8911 0.0
V21752 n0_13741_9057 n2_13741_9057 0.0
V21753 n0_13741_9090 n2_13741_9090 0.0
V21754 n0_13741_9273 n2_13741_9273 0.0
V21755 n0_13741_9306 n2_13741_9306 0.0
V21756 n0_13741_9489 n2_13741_9489 0.0
V21757 n0_13741_9522 n2_13741_9522 0.0
V21758 n0_13741_9705 n2_13741_9705 0.0
V21759 n0_13741_9738 n2_13741_9738 0.0
V21760 n0_13741_9775 n2_13741_9775 0.0
V21761 n0_13741_9921 n2_13741_9921 0.0
V21762 n0_13741_9954 n2_13741_9954 0.0
V21763 n0_13741_9991 n2_13741_9991 0.0
V21764 n0_13741_10137 n2_13741_10137 0.0
V21765 n0_13741_10170 n2_13741_10170 0.0
V21766 n0_13741_10353 n2_13741_10353 0.0
V21767 n0_13741_10386 n2_13741_10386 0.0
V21768 n0_13741_10569 n2_13741_10569 0.0
V21769 n0_13741_10785 n2_13741_10785 0.0
V21770 n0_13741_10818 n2_13741_10818 0.0
V21771 n0_13741_10832 n2_13741_10832 0.0
V21772 n0_13741_11001 n2_13741_11001 0.0
V21773 n0_13741_11034 n2_13741_11034 0.0
V21774 n0_13741_11048 n2_13741_11048 0.0
V21775 n0_13741_11217 n2_13741_11217 0.0
V21776 n0_13741_11250 n2_13741_11250 0.0
V21777 n0_13741_11433 n2_13741_11433 0.0
V21778 n0_13741_11466 n2_13741_11466 0.0
V21779 n0_13741_11649 n2_13741_11649 0.0
V21780 n0_13741_11682 n2_13741_11682 0.0
V21781 n0_13741_11865 n2_13741_11865 0.0
V21782 n0_13741_11898 n2_13741_11898 0.0
V21783 n0_13741_11912 n2_13741_11912 0.0
V21784 n0_13741_12081 n2_13741_12081 0.0
V21785 n0_13741_12114 n2_13741_12114 0.0
V21786 n0_13741_12128 n2_13741_12128 0.0
V21787 n0_13741_12297 n2_13741_12297 0.0
V21788 n0_13741_12330 n2_13741_12330 0.0
V21789 n0_13741_12513 n2_13741_12513 0.0
V21790 n0_13741_12546 n2_13741_12546 0.0
V21791 n0_13741_12729 n2_13741_12729 0.0
V21792 n0_13741_12762 n2_13741_12762 0.0
V21793 n0_13741_12776 n2_13741_12776 0.0
V21794 n0_13741_12945 n2_13741_12945 0.0
V21795 n0_13741_12978 n2_13741_12978 0.0
V21796 n0_13741_12992 n2_13741_12992 0.0
V21797 n0_13741_13161 n2_13741_13161 0.0
V21798 n0_13741_13194 n2_13741_13194 0.0
V21799 n0_13741_13377 n2_13741_13377 0.0
V21800 n0_13741_13410 n2_13741_13410 0.0
V21801 n0_13741_13423 n2_13741_13423 0.0
V21802 n0_13741_13593 n2_13741_13593 0.0
V21803 n0_13741_13626 n2_13741_13626 0.0
V21804 n0_13741_13809 n2_13741_13809 0.0
V21805 n0_13741_13842 n2_13741_13842 0.0
V21806 n0_13880_8409 n2_13880_8409 0.0
V21807 n0_13880_10569 n2_13880_10569 0.0
V21808 n0_13880_10602 n2_13880_10602 0.0
V21809 n0_13880_12776 n2_13880_12776 0.0
V21810 n0_13929_7329 n2_13929_7329 0.0
V21811 n0_13929_7362 n2_13929_7362 0.0
V21812 n0_13929_7545 n2_13929_7545 0.0
V21813 n0_13929_7578 n2_13929_7578 0.0
V21814 n0_13929_7761 n2_13929_7761 0.0
V21815 n0_13929_7794 n2_13929_7794 0.0
V21816 n0_13929_7831 n2_13929_7831 0.0
V21817 n0_13929_7977 n2_13929_7977 0.0
V21818 n0_13929_8010 n2_13929_8010 0.0
V21819 n0_13929_8193 n2_13929_8193 0.0
V21820 n0_13929_8226 n2_13929_8226 0.0
V21821 n0_13929_8409 n2_13929_8409 0.0
V21822 n0_13929_8442 n2_13929_8442 0.0
V21823 n0_13929_8625 n2_13929_8625 0.0
V21824 n0_13929_8658 n2_13929_8658 0.0
V21825 n0_13929_8695 n2_13929_8695 0.0
V21826 n0_13929_8841 n2_13929_8841 0.0
V21827 n0_13929_8874 n2_13929_8874 0.0
V21828 n0_13929_8911 n2_13929_8911 0.0
V21829 n0_13929_9057 n2_13929_9057 0.0
V21830 n0_13929_9090 n2_13929_9090 0.0
V21831 n0_13929_9273 n2_13929_9273 0.0
V21832 n0_13929_9306 n2_13929_9306 0.0
V21833 n0_13929_9705 n2_13929_9705 0.0
V21834 n0_13929_9738 n2_13929_9738 0.0
V21835 n0_13929_9775 n2_13929_9775 0.0
V21836 n0_13929_9921 n2_13929_9921 0.0
V21837 n0_13929_9954 n2_13929_9954 0.0
V21838 n0_13929_9991 n2_13929_9991 0.0
V21839 n0_13929_10137 n2_13929_10137 0.0
V21840 n0_13929_10170 n2_13929_10170 0.0
V21841 n0_13929_10353 n2_13929_10353 0.0
V21842 n0_13929_10386 n2_13929_10386 0.0
V21843 n0_13929_10569 n2_13929_10569 0.0
V21844 n0_13929_10602 n2_13929_10602 0.0
V21845 n0_13929_10785 n2_13929_10785 0.0
V21846 n0_13929_10818 n2_13929_10818 0.0
V21847 n0_13929_10832 n2_13929_10832 0.0
V21848 n0_13929_11001 n2_13929_11001 0.0
V21849 n0_13929_11034 n2_13929_11034 0.0
V21850 n0_13929_11048 n2_13929_11048 0.0
V21851 n0_13929_11217 n2_13929_11217 0.0
V21852 n0_13929_11250 n2_13929_11250 0.0
V21853 n0_13929_11433 n2_13929_11433 0.0
V21854 n0_13929_11466 n2_13929_11466 0.0
V21855 n0_13929_11865 n2_13929_11865 0.0
V21856 n0_13929_11898 n2_13929_11898 0.0
V21857 n0_13929_11912 n2_13929_11912 0.0
V21858 n0_13929_12081 n2_13929_12081 0.0
V21859 n0_13929_12114 n2_13929_12114 0.0
V21860 n0_13929_12128 n2_13929_12128 0.0
V21861 n0_13929_12297 n2_13929_12297 0.0
V21862 n0_13929_12330 n2_13929_12330 0.0
V21863 n0_13929_12513 n2_13929_12513 0.0
V21864 n0_13929_12546 n2_13929_12546 0.0
V21865 n0_13929_12729 n2_13929_12729 0.0
V21866 n0_13929_12762 n2_13929_12762 0.0
V21867 n0_13929_12776 n2_13929_12776 0.0
V21868 n0_13929_12945 n2_13929_12945 0.0
V21869 n0_13929_12978 n2_13929_12978 0.0
V21870 n0_13929_12992 n2_13929_12992 0.0
V21871 n0_13929_13161 n2_13929_13161 0.0
V21872 n0_13929_13194 n2_13929_13194 0.0
V21873 n0_13929_13377 n2_13929_13377 0.0
V21874 n0_13929_13410 n2_13929_13410 0.0
V21875 n0_13929_13423 n2_13929_13423 0.0
V21876 n0_13929_13593 n2_13929_13593 0.0
V21877 n0_13929_13626 n2_13929_13626 0.0
V21878 n0_13929_13809 n2_13929_13809 0.0
V21879 n0_13929_13842 n2_13929_13842 0.0
V21880 n0_14866_201 n2_14866_201 0.0
V21881 n0_14866_234 n2_14866_234 0.0
V21882 n0_14866_417 n2_14866_417 0.0
V21883 n0_14866_450 n2_14866_450 0.0
V21884 n0_14866_633 n2_14866_633 0.0
V21885 n0_14866_666 n2_14866_666 0.0
V21886 n0_14866_849 n2_14866_849 0.0
V21887 n0_14866_882 n2_14866_882 0.0
V21888 n0_14866_1065 n2_14866_1065 0.0
V21889 n0_14866_1098 n2_14866_1098 0.0
V21890 n0_14866_1281 n2_14866_1281 0.0
V21891 n0_14866_1314 n2_14866_1314 0.0
V21892 n0_14866_1497 n2_14866_1497 0.0
V21893 n0_14866_1530 n2_14866_1530 0.0
V21894 n0_14866_1713 n2_14866_1713 0.0
V21895 n0_14866_1746 n2_14866_1746 0.0
V21896 n0_14866_1783 n2_14866_1783 0.0
V21897 n0_14866_1929 n2_14866_1929 0.0
V21898 n0_14866_1962 n2_14866_1962 0.0
V21899 n0_14866_2145 n2_14866_2145 0.0
V21900 n0_14866_2178 n2_14866_2178 0.0
V21901 n0_14866_2361 n2_14866_2361 0.0
V21902 n0_14866_2394 n2_14866_2394 0.0
V21903 n0_14866_2431 n2_14866_2431 0.0
V21904 n0_14866_2577 n2_14866_2577 0.0
V21905 n0_14866_2610 n2_14866_2610 0.0
V21906 n0_14866_2793 n2_14866_2793 0.0
V21907 n0_14866_2826 n2_14866_2826 0.0
V21908 n0_14866_2863 n2_14866_2863 0.0
V21909 n0_14866_3009 n2_14866_3009 0.0
V21910 n0_14866_3042 n2_14866_3042 0.0
V21911 n0_14866_3225 n2_14866_3225 0.0
V21912 n0_14866_3258 n2_14866_3258 0.0
V21913 n0_14866_3295 n2_14866_3295 0.0
V21914 n0_14866_3441 n2_14866_3441 0.0
V21915 n0_14866_3474 n2_14866_3474 0.0
V21916 n0_14866_3511 n2_14866_3511 0.0
V21917 n0_14866_3657 n2_14866_3657 0.0
V21918 n0_14866_3690 n2_14866_3690 0.0
V21919 n0_14866_3873 n2_14866_3873 0.0
V21920 n0_14866_3906 n2_14866_3906 0.0
V21921 n0_14866_3943 n2_14866_3943 0.0
V21922 n0_14866_4089 n2_14866_4089 0.0
V21923 n0_14866_4122 n2_14866_4122 0.0
V21924 n0_14866_4159 n2_14866_4159 0.0
V21925 n0_14866_4305 n2_14866_4305 0.0
V21926 n0_14866_4338 n2_14866_4338 0.0
V21927 n0_14866_4375 n2_14866_4375 0.0
V21928 n0_14866_4521 n2_14866_4521 0.0
V21929 n0_14866_4554 n2_14866_4554 0.0
V21930 n0_14866_4591 n2_14866_4591 0.0
V21931 n0_14866_4737 n2_14866_4737 0.0
V21932 n0_14866_4770 n2_14866_4770 0.0
V21933 n0_14866_4807 n2_14866_4807 0.0
V21934 n0_14866_4953 n2_14866_4953 0.0
V21935 n0_14866_5169 n2_14866_5169 0.0
V21936 n0_14866_5202 n2_14866_5202 0.0
V21937 n0_14866_5239 n2_14866_5239 0.0
V21938 n0_14866_5385 n2_14866_5385 0.0
V21939 n0_14866_5418 n2_14866_5418 0.0
V21940 n0_14866_5455 n2_14866_5455 0.0
V21941 n0_14866_5601 n2_14866_5601 0.0
V21942 n0_14866_5634 n2_14866_5634 0.0
V21943 n0_14866_5671 n2_14866_5671 0.0
V21944 n0_14866_5817 n2_14866_5817 0.0
V21945 n0_14866_5850 n2_14866_5850 0.0
V21946 n0_14866_6033 n2_14866_6033 0.0
V21947 n0_14866_6066 n2_14866_6066 0.0
V21948 n0_14866_6249 n2_14866_6249 0.0
V21949 n0_14866_6282 n2_14866_6282 0.0
V21950 n0_14866_6319 n2_14866_6319 0.0
V21951 n0_14866_6465 n2_14866_6465 0.0
V21952 n0_14866_6498 n2_14866_6498 0.0
V21953 n0_14866_6535 n2_14866_6535 0.0
V21954 n0_14866_6681 n2_14866_6681 0.0
V21955 n0_14866_6714 n2_14866_6714 0.0
V21956 n0_14866_6897 n2_14866_6897 0.0
V21957 n0_14866_6930 n2_14866_6930 0.0
V21958 n0_14866_7113 n2_14866_7113 0.0
V21959 n0_14866_7146 n2_14866_7146 0.0
V21960 n0_14866_7329 n2_14866_7329 0.0
V21961 n0_14866_7362 n2_14866_7362 0.0
V21962 n0_14866_7545 n2_14866_7545 0.0
V21963 n0_14866_7578 n2_14866_7578 0.0
V21964 n0_14866_7761 n2_14866_7761 0.0
V21965 n0_14866_7794 n2_14866_7794 0.0
V21966 n0_14866_7831 n2_14866_7831 0.0
V21967 n0_14866_7977 n2_14866_7977 0.0
V21968 n0_14866_8010 n2_14866_8010 0.0
V21969 n0_14866_8193 n2_14866_8193 0.0
V21970 n0_14866_8226 n2_14866_8226 0.0
V21971 n0_14866_8409 n2_14866_8409 0.0
V21972 n0_14866_8442 n2_14866_8442 0.0
V21973 n0_14866_8625 n2_14866_8625 0.0
V21974 n0_14866_8658 n2_14866_8658 0.0
V21975 n0_14866_8841 n2_14866_8841 0.0
V21976 n0_14866_8874 n2_14866_8874 0.0
V21977 n0_14866_8911 n2_14866_8911 0.0
V21978 n0_14866_9057 n2_14866_9057 0.0
V21979 n0_14866_9090 n2_14866_9090 0.0
V21980 n0_14866_9273 n2_14866_9273 0.0
V21981 n0_14866_9306 n2_14866_9306 0.0
V21982 n0_14866_9489 n2_14866_9489 0.0
V21983 n0_14866_9522 n2_14866_9522 0.0
V21984 n0_14866_9705 n2_14866_9705 0.0
V21985 n0_14866_9738 n2_14866_9738 0.0
V21986 n0_14866_9921 n2_14866_9921 0.0
V21987 n0_14866_9954 n2_14866_9954 0.0
V21988 n0_14866_9991 n2_14866_9991 0.0
V21989 n0_14866_10137 n2_14866_10137 0.0
V21990 n0_14866_10170 n2_14866_10170 0.0
V21991 n0_14866_10353 n2_14866_10353 0.0
V21992 n0_14866_10386 n2_14866_10386 0.0
V21993 n0_14866_10569 n2_14866_10569 0.0
V21994 n0_14866_10785 n2_14866_10785 0.0
V21995 n0_14866_10818 n2_14866_10818 0.0
V21996 n0_14866_11001 n2_14866_11001 0.0
V21997 n0_14866_11034 n2_14866_11034 0.0
V21998 n0_14866_11048 n2_14866_11048 0.0
V21999 n0_14866_11217 n2_14866_11217 0.0
V22000 n0_14866_11250 n2_14866_11250 0.0
V22001 n0_14866_11433 n2_14866_11433 0.0
V22002 n0_14866_11466 n2_14866_11466 0.0
V22003 n0_14866_11649 n2_14866_11649 0.0
V22004 n0_14866_11682 n2_14866_11682 0.0
V22005 n0_14866_11865 n2_14866_11865 0.0
V22006 n0_14866_11898 n2_14866_11898 0.0
V22007 n0_14866_12081 n2_14866_12081 0.0
V22008 n0_14866_12114 n2_14866_12114 0.0
V22009 n0_14866_12128 n2_14866_12128 0.0
V22010 n0_14866_12135 n2_14866_12135 0.0
V22011 n0_14866_12297 n2_14866_12297 0.0
V22012 n0_14866_12330 n2_14866_12330 0.0
V22013 n0_14866_12513 n2_14866_12513 0.0
V22014 n0_14866_12546 n2_14866_12546 0.0
V22015 n0_14866_12729 n2_14866_12729 0.0
V22016 n0_14866_12762 n2_14866_12762 0.0
V22017 n0_14866_12776 n2_14866_12776 0.0
V22018 n0_14866_12945 n2_14866_12945 0.0
V22019 n0_14866_12978 n2_14866_12978 0.0
V22020 n0_14866_12992 n2_14866_12992 0.0
V22021 n0_14866_13161 n2_14866_13161 0.0
V22022 n0_14866_13194 n2_14866_13194 0.0
V22023 n0_14866_13377 n2_14866_13377 0.0
V22024 n0_14866_13410 n2_14866_13410 0.0
V22025 n0_14866_13423 n2_14866_13423 0.0
V22026 n0_14866_13593 n2_14866_13593 0.0
V22027 n0_14866_13626 n2_14866_13626 0.0
V22028 n0_14866_13809 n2_14866_13809 0.0
V22029 n0_14866_13842 n2_14866_13842 0.0
V22030 n0_14866_14025 n2_14866_14025 0.0
V22031 n0_14866_14058 n2_14866_14058 0.0
V22032 n0_14866_14241 n2_14866_14241 0.0
V22033 n0_14866_14274 n2_14866_14274 0.0
V22034 n0_14866_14457 n2_14866_14457 0.0
V22035 n0_14866_14490 n2_14866_14490 0.0
V22036 n0_14866_14511 n2_14866_14511 0.0
V22037 n0_14866_14673 n2_14866_14673 0.0
V22038 n0_14866_14706 n2_14866_14706 0.0
V22039 n0_14866_14889 n2_14866_14889 0.0
V22040 n0_14866_14922 n2_14866_14922 0.0
V22041 n0_14866_14943 n2_14866_14943 0.0
V22042 n0_14866_15138 n2_14866_15138 0.0
V22043 n0_14866_15159 n2_14866_15159 0.0
V22044 n0_14866_15321 n2_14866_15321 0.0
V22045 n0_14866_15354 n2_14866_15354 0.0
V22046 n0_14866_15368 n2_14866_15368 0.0
V22047 n0_14866_15537 n2_14866_15537 0.0
V22048 n0_14866_15570 n2_14866_15570 0.0
V22049 n0_14866_15584 n2_14866_15584 0.0
V22050 n0_14866_15753 n2_14866_15753 0.0
V22051 n0_14866_15786 n2_14866_15786 0.0
V22052 n0_14866_15800 n2_14866_15800 0.0
V22053 n0_14866_15969 n2_14866_15969 0.0
V22054 n0_14866_16002 n2_14866_16002 0.0
V22055 n0_14866_16185 n2_14866_16185 0.0
V22056 n0_14866_16401 n2_14866_16401 0.0
V22057 n0_14866_16434 n2_14866_16434 0.0
V22058 n0_14866_16448 n2_14866_16448 0.0
V22059 n0_14866_16617 n2_14866_16617 0.0
V22060 n0_14866_16650 n2_14866_16650 0.0
V22061 n0_14866_16687 n2_14866_16687 0.0
V22062 n0_14866_16833 n2_14866_16833 0.0
V22063 n0_14866_16866 n2_14866_16866 0.0
V22064 n0_14866_17049 n2_14866_17049 0.0
V22065 n0_14866_17082 n2_14866_17082 0.0
V22066 n0_14866_17096 n2_14866_17096 0.0
V22067 n0_14866_17265 n2_14866_17265 0.0
V22068 n0_14866_17298 n2_14866_17298 0.0
V22069 n0_14866_17481 n2_14866_17481 0.0
V22070 n0_14866_17514 n2_14866_17514 0.0
V22071 n0_14866_17528 n2_14866_17528 0.0
V22072 n0_14866_17697 n2_14866_17697 0.0
V22073 n0_14866_17730 n2_14866_17730 0.0
V22074 n0_14866_17913 n2_14866_17913 0.0
V22075 n0_14866_17946 n2_14866_17946 0.0
V22076 n0_14866_17983 n2_14866_17983 0.0
V22077 n0_14866_18129 n2_14866_18129 0.0
V22078 n0_14866_18162 n2_14866_18162 0.0
V22079 n0_14866_18176 n2_14866_18176 0.0
V22080 n0_14866_18345 n2_14866_18345 0.0
V22081 n0_14866_18378 n2_14866_18378 0.0
V22082 n0_14866_18561 n2_14866_18561 0.0
V22083 n0_14866_18594 n2_14866_18594 0.0
V22084 n0_14866_18608 n2_14866_18608 0.0
V22085 n0_14866_18777 n2_14866_18777 0.0
V22086 n0_14866_18810 n2_14866_18810 0.0
V22087 n0_14866_18993 n2_14866_18993 0.0
V22088 n0_14866_19026 n2_14866_19026 0.0
V22089 n0_14866_19209 n2_14866_19209 0.0
V22090 n0_14866_19242 n2_14866_19242 0.0
V22091 n0_14866_19256 n2_14866_19256 0.0
V22092 n0_14866_19263 n2_14866_19263 0.0
V22093 n0_14866_19425 n2_14866_19425 0.0
V22094 n0_14866_19458 n2_14866_19458 0.0
V22095 n0_14866_19641 n2_14866_19641 0.0
V22096 n0_14866_19674 n2_14866_19674 0.0
V22097 n0_14866_19857 n2_14866_19857 0.0
V22098 n0_14866_19890 n2_14866_19890 0.0
V22099 n0_14866_20073 n2_14866_20073 0.0
V22100 n0_14866_20106 n2_14866_20106 0.0
V22101 n0_14866_20289 n2_14866_20289 0.0
V22102 n0_14866_20322 n2_14866_20322 0.0
V22103 n0_14866_20505 n2_14866_20505 0.0
V22104 n0_14866_20538 n2_14866_20538 0.0
V22105 n0_14866_20754 n2_14866_20754 0.0
V22106 n0_14866_20937 n2_14866_20937 0.0
V22107 n0_14866_20970 n2_14866_20970 0.0
V22108 n0_14958_201 n2_14958_201 0.0
V22109 n0_14958_234 n2_14958_234 0.0
V22110 n0_14958_417 n2_14958_417 0.0
V22111 n0_14958_450 n2_14958_450 0.0
V22112 n0_14958_633 n2_14958_633 0.0
V22113 n0_14958_666 n2_14958_666 0.0
V22114 n0_14958_849 n2_14958_849 0.0
V22115 n0_14958_882 n2_14958_882 0.0
V22116 n0_14958_1065 n2_14958_1065 0.0
V22117 n0_14958_1098 n2_14958_1098 0.0
V22118 n0_14958_1281 n2_14958_1281 0.0
V22119 n0_14958_1314 n2_14958_1314 0.0
V22120 n0_14958_1497 n2_14958_1497 0.0
V22121 n0_14958_1530 n2_14958_1530 0.0
V22122 n0_14958_1713 n2_14958_1713 0.0
V22123 n0_14958_1746 n2_14958_1746 0.0
V22124 n0_14958_1783 n2_14958_1783 0.0
V22125 n0_14958_1929 n2_14958_1929 0.0
V22126 n0_14958_1962 n2_14958_1962 0.0
V22127 n0_14958_2145 n2_14958_2145 0.0
V22128 n0_14958_2178 n2_14958_2178 0.0
V22129 n0_14958_2361 n2_14958_2361 0.0
V22130 n0_14958_2394 n2_14958_2394 0.0
V22131 n0_14958_2431 n2_14958_2431 0.0
V22132 n0_14958_2577 n2_14958_2577 0.0
V22133 n0_14958_2610 n2_14958_2610 0.0
V22134 n0_14958_2793 n2_14958_2793 0.0
V22135 n0_14958_2826 n2_14958_2826 0.0
V22136 n0_14958_2863 n2_14958_2863 0.0
V22137 n0_14958_3009 n2_14958_3009 0.0
V22138 n0_14958_3042 n2_14958_3042 0.0
V22139 n0_14958_3225 n2_14958_3225 0.0
V22140 n0_14958_3258 n2_14958_3258 0.0
V22141 n0_14958_3295 n2_14958_3295 0.0
V22142 n0_14958_3441 n2_14958_3441 0.0
V22143 n0_14958_3474 n2_14958_3474 0.0
V22144 n0_14958_3511 n2_14958_3511 0.0
V22145 n0_14958_3657 n2_14958_3657 0.0
V22146 n0_14958_3690 n2_14958_3690 0.0
V22147 n0_14958_3873 n2_14958_3873 0.0
V22148 n0_14958_3906 n2_14958_3906 0.0
V22149 n0_14958_3943 n2_14958_3943 0.0
V22150 n0_14958_4089 n2_14958_4089 0.0
V22151 n0_14958_4122 n2_14958_4122 0.0
V22152 n0_14958_4159 n2_14958_4159 0.0
V22153 n0_14958_4305 n2_14958_4305 0.0
V22154 n0_14958_4338 n2_14958_4338 0.0
V22155 n0_14958_4375 n2_14958_4375 0.0
V22156 n0_14958_4521 n2_14958_4521 0.0
V22157 n0_14958_4554 n2_14958_4554 0.0
V22158 n0_14958_4591 n2_14958_4591 0.0
V22159 n0_14958_4737 n2_14958_4737 0.0
V22160 n0_14958_4770 n2_14958_4770 0.0
V22161 n0_14958_4807 n2_14958_4807 0.0
V22162 n0_14958_4953 n2_14958_4953 0.0
V22163 n0_14958_4986 n2_14958_4986 0.0
V22164 n0_14958_5169 n2_14958_5169 0.0
V22165 n0_14958_5202 n2_14958_5202 0.0
V22166 n0_14958_5239 n2_14958_5239 0.0
V22167 n0_14958_5385 n2_14958_5385 0.0
V22168 n0_14958_5418 n2_14958_5418 0.0
V22169 n0_14958_5455 n2_14958_5455 0.0
V22170 n0_14958_5601 n2_14958_5601 0.0
V22171 n0_14958_5634 n2_14958_5634 0.0
V22172 n0_14958_5671 n2_14958_5671 0.0
V22173 n0_14958_5817 n2_14958_5817 0.0
V22174 n0_14958_5850 n2_14958_5850 0.0
V22175 n0_14958_6033 n2_14958_6033 0.0
V22176 n0_14958_6066 n2_14958_6066 0.0
V22177 n0_14958_15105 n2_14958_15105 0.0
V22178 n0_14958_15138 n2_14958_15138 0.0
V22179 n0_14958_15159 n2_14958_15159 0.0
V22180 n0_14958_15321 n2_14958_15321 0.0
V22181 n0_14958_15354 n2_14958_15354 0.0
V22182 n0_14958_15368 n2_14958_15368 0.0
V22183 n0_14958_15537 n2_14958_15537 0.0
V22184 n0_14958_15570 n2_14958_15570 0.0
V22185 n0_14958_15584 n2_14958_15584 0.0
V22186 n0_14958_15753 n2_14958_15753 0.0
V22187 n0_14958_15786 n2_14958_15786 0.0
V22188 n0_14958_15800 n2_14958_15800 0.0
V22189 n0_14958_15969 n2_14958_15969 0.0
V22190 n0_14958_16002 n2_14958_16002 0.0
V22191 n0_14958_16185 n2_14958_16185 0.0
V22192 n0_14958_16218 n2_14958_16218 0.0
V22193 n0_14958_16401 n2_14958_16401 0.0
V22194 n0_14958_16434 n2_14958_16434 0.0
V22195 n0_14958_16448 n2_14958_16448 0.0
V22196 n0_14958_16617 n2_14958_16617 0.0
V22197 n0_14958_16650 n2_14958_16650 0.0
V22198 n0_14958_16687 n2_14958_16687 0.0
V22199 n0_14958_16833 n2_14958_16833 0.0
V22200 n0_14958_16866 n2_14958_16866 0.0
V22201 n0_14958_17049 n2_14958_17049 0.0
V22202 n0_14958_17082 n2_14958_17082 0.0
V22203 n0_14958_17096 n2_14958_17096 0.0
V22204 n0_14958_17265 n2_14958_17265 0.0
V22205 n0_14958_17298 n2_14958_17298 0.0
V22206 n0_14958_17481 n2_14958_17481 0.0
V22207 n0_14958_17514 n2_14958_17514 0.0
V22208 n0_14958_17528 n2_14958_17528 0.0
V22209 n0_14958_17697 n2_14958_17697 0.0
V22210 n0_14958_17730 n2_14958_17730 0.0
V22211 n0_14958_17913 n2_14958_17913 0.0
V22212 n0_14958_17946 n2_14958_17946 0.0
V22213 n0_14958_17983 n2_14958_17983 0.0
V22214 n0_14958_18129 n2_14958_18129 0.0
V22215 n0_14958_18162 n2_14958_18162 0.0
V22216 n0_14958_18176 n2_14958_18176 0.0
V22217 n0_14958_18345 n2_14958_18345 0.0
V22218 n0_14958_18378 n2_14958_18378 0.0
V22219 n0_14958_18561 n2_14958_18561 0.0
V22220 n0_14958_18594 n2_14958_18594 0.0
V22221 n0_14958_18608 n2_14958_18608 0.0
V22222 n0_14958_18777 n2_14958_18777 0.0
V22223 n0_14958_18810 n2_14958_18810 0.0
V22224 n0_14958_18993 n2_14958_18993 0.0
V22225 n0_14958_19026 n2_14958_19026 0.0
V22226 n0_14958_19209 n2_14958_19209 0.0
V22227 n0_14958_19242 n2_14958_19242 0.0
V22228 n0_14958_19256 n2_14958_19256 0.0
V22229 n0_14958_19263 n2_14958_19263 0.0
V22230 n0_14958_19425 n2_14958_19425 0.0
V22231 n0_14958_19458 n2_14958_19458 0.0
V22232 n0_14958_19641 n2_14958_19641 0.0
V22233 n0_14958_19674 n2_14958_19674 0.0
V22234 n0_14958_19857 n2_14958_19857 0.0
V22235 n0_14958_19890 n2_14958_19890 0.0
V22236 n0_14958_20073 n2_14958_20073 0.0
V22237 n0_14958_20106 n2_14958_20106 0.0
V22238 n0_14958_20289 n2_14958_20289 0.0
V22239 n0_14958_20322 n2_14958_20322 0.0
V22240 n0_14958_20505 n2_14958_20505 0.0
V22241 n0_14958_20538 n2_14958_20538 0.0
V22242 n0_14958_20721 n2_14958_20721 0.0
V22243 n0_14958_20754 n2_14958_20754 0.0
V22244 n0_14958_20937 n2_14958_20937 0.0
V22245 n0_14958_20970 n2_14958_20970 0.0
V22246 n0_15005_417 n2_15005_417 0.0
V22247 n0_15005_450 n2_15005_450 0.0
V22248 n0_15005_1530 n2_15005_1530 0.0
V22249 n0_15005_2793 n2_15005_2793 0.0
V22250 n0_15005_3873 n2_15005_3873 0.0
V22251 n0_15005_3906 n2_15005_3906 0.0
V22252 n0_15005_4953 n2_15005_4953 0.0
V22253 n0_15005_4986 n2_15005_4986 0.0
V22254 n0_15005_6033 n2_15005_6033 0.0
V22255 n0_15005_6066 n2_15005_6066 0.0
V22256 n0_15005_8409 n2_15005_8409 0.0
V22257 n0_15005_10569 n2_15005_10569 0.0
V22258 n0_15005_10602 n2_15005_10602 0.0
V22259 n0_15005_12776 n2_15005_12776 0.0
V22260 n0_15005_15105 n2_15005_15105 0.0
V22261 n0_15005_15138 n2_15005_15138 0.0
V22262 n0_15005_15159 n2_15005_15159 0.0
V22263 n0_15005_16185 n2_15005_16185 0.0
V22264 n0_15005_16218 n2_15005_16218 0.0
V22265 n0_15005_17298 n2_15005_17298 0.0
V22266 n0_15005_19641 n2_15005_19641 0.0
V22267 n0_15005_19674 n2_15005_19674 0.0
V22268 n0_15005_20721 n2_15005_20721 0.0
V22269 n0_15005_20754 n2_15005_20754 0.0
V22270 n0_15054_201 n2_15054_201 0.0
V22271 n0_15054_234 n2_15054_234 0.0
V22272 n0_15054_417 n2_15054_417 0.0
V22273 n0_15054_450 n2_15054_450 0.0
V22274 n0_15054_633 n2_15054_633 0.0
V22275 n0_15054_666 n2_15054_666 0.0
V22276 n0_15054_849 n2_15054_849 0.0
V22277 n0_15054_882 n2_15054_882 0.0
V22278 n0_15054_1065 n2_15054_1065 0.0
V22279 n0_15054_1098 n2_15054_1098 0.0
V22280 n0_15054_1281 n2_15054_1281 0.0
V22281 n0_15054_1314 n2_15054_1314 0.0
V22282 n0_15054_1497 n2_15054_1497 0.0
V22283 n0_15054_1530 n2_15054_1530 0.0
V22284 n0_15054_1713 n2_15054_1713 0.0
V22285 n0_15054_1746 n2_15054_1746 0.0
V22286 n0_15054_1783 n2_15054_1783 0.0
V22287 n0_15054_1929 n2_15054_1929 0.0
V22288 n0_15054_1962 n2_15054_1962 0.0
V22289 n0_15054_2145 n2_15054_2145 0.0
V22290 n0_15054_2178 n2_15054_2178 0.0
V22291 n0_15054_2361 n2_15054_2361 0.0
V22292 n0_15054_2394 n2_15054_2394 0.0
V22293 n0_15054_2431 n2_15054_2431 0.0
V22294 n0_15054_2577 n2_15054_2577 0.0
V22295 n0_15054_2610 n2_15054_2610 0.0
V22296 n0_15054_2793 n2_15054_2793 0.0
V22297 n0_15054_2826 n2_15054_2826 0.0
V22298 n0_15054_2863 n2_15054_2863 0.0
V22299 n0_15054_3009 n2_15054_3009 0.0
V22300 n0_15054_3042 n2_15054_3042 0.0
V22301 n0_15054_3225 n2_15054_3225 0.0
V22302 n0_15054_3258 n2_15054_3258 0.0
V22303 n0_15054_3295 n2_15054_3295 0.0
V22304 n0_15054_3441 n2_15054_3441 0.0
V22305 n0_15054_3474 n2_15054_3474 0.0
V22306 n0_15054_3511 n2_15054_3511 0.0
V22307 n0_15054_3657 n2_15054_3657 0.0
V22308 n0_15054_3690 n2_15054_3690 0.0
V22309 n0_15054_3873 n2_15054_3873 0.0
V22310 n0_15054_3906 n2_15054_3906 0.0
V22311 n0_15054_3943 n2_15054_3943 0.0
V22312 n0_15054_4089 n2_15054_4089 0.0
V22313 n0_15054_4122 n2_15054_4122 0.0
V22314 n0_15054_4159 n2_15054_4159 0.0
V22315 n0_15054_4305 n2_15054_4305 0.0
V22316 n0_15054_4338 n2_15054_4338 0.0
V22317 n0_15054_4375 n2_15054_4375 0.0
V22318 n0_15054_4521 n2_15054_4521 0.0
V22319 n0_15054_4554 n2_15054_4554 0.0
V22320 n0_15054_4591 n2_15054_4591 0.0
V22321 n0_15054_4737 n2_15054_4737 0.0
V22322 n0_15054_4770 n2_15054_4770 0.0
V22323 n0_15054_4807 n2_15054_4807 0.0
V22324 n0_15054_4953 n2_15054_4953 0.0
V22325 n0_15054_4986 n2_15054_4986 0.0
V22326 n0_15054_5169 n2_15054_5169 0.0
V22327 n0_15054_5202 n2_15054_5202 0.0
V22328 n0_15054_5239 n2_15054_5239 0.0
V22329 n0_15054_5385 n2_15054_5385 0.0
V22330 n0_15054_5418 n2_15054_5418 0.0
V22331 n0_15054_5455 n2_15054_5455 0.0
V22332 n0_15054_5601 n2_15054_5601 0.0
V22333 n0_15054_5634 n2_15054_5634 0.0
V22334 n0_15054_5671 n2_15054_5671 0.0
V22335 n0_15054_5817 n2_15054_5817 0.0
V22336 n0_15054_5850 n2_15054_5850 0.0
V22337 n0_15054_6033 n2_15054_6033 0.0
V22338 n0_15054_6066 n2_15054_6066 0.0
V22339 n0_15054_6249 n2_15054_6249 0.0
V22340 n0_15054_6282 n2_15054_6282 0.0
V22341 n0_15054_6319 n2_15054_6319 0.0
V22342 n0_15054_6465 n2_15054_6465 0.0
V22343 n0_15054_6498 n2_15054_6498 0.0
V22344 n0_15054_6535 n2_15054_6535 0.0
V22345 n0_15054_6681 n2_15054_6681 0.0
V22346 n0_15054_6714 n2_15054_6714 0.0
V22347 n0_15054_6897 n2_15054_6897 0.0
V22348 n0_15054_6930 n2_15054_6930 0.0
V22349 n0_15054_7113 n2_15054_7113 0.0
V22350 n0_15054_7329 n2_15054_7329 0.0
V22351 n0_15054_7362 n2_15054_7362 0.0
V22352 n0_15054_7545 n2_15054_7545 0.0
V22353 n0_15054_7578 n2_15054_7578 0.0
V22354 n0_15054_7761 n2_15054_7761 0.0
V22355 n0_15054_7794 n2_15054_7794 0.0
V22356 n0_15054_7831 n2_15054_7831 0.0
V22357 n0_15054_7977 n2_15054_7977 0.0
V22358 n0_15054_8010 n2_15054_8010 0.0
V22359 n0_15054_8193 n2_15054_8193 0.0
V22360 n0_15054_8226 n2_15054_8226 0.0
V22361 n0_15054_8409 n2_15054_8409 0.0
V22362 n0_15054_8442 n2_15054_8442 0.0
V22363 n0_15054_8625 n2_15054_8625 0.0
V22364 n0_15054_8658 n2_15054_8658 0.0
V22365 n0_15054_8841 n2_15054_8841 0.0
V22366 n0_15054_8874 n2_15054_8874 0.0
V22367 n0_15054_8911 n2_15054_8911 0.0
V22368 n0_15054_9057 n2_15054_9057 0.0
V22369 n0_15054_9090 n2_15054_9090 0.0
V22370 n0_15054_9273 n2_15054_9273 0.0
V22371 n0_15054_9306 n2_15054_9306 0.0
V22372 n0_15054_9705 n2_15054_9705 0.0
V22373 n0_15054_9738 n2_15054_9738 0.0
V22374 n0_15054_9921 n2_15054_9921 0.0
V22375 n0_15054_9954 n2_15054_9954 0.0
V22376 n0_15054_9991 n2_15054_9991 0.0
V22377 n0_15054_10137 n2_15054_10137 0.0
V22378 n0_15054_10170 n2_15054_10170 0.0
V22379 n0_15054_10353 n2_15054_10353 0.0
V22380 n0_15054_10386 n2_15054_10386 0.0
V22381 n0_15054_10569 n2_15054_10569 0.0
V22382 n0_15054_10602 n2_15054_10602 0.0
V22383 n0_15054_10785 n2_15054_10785 0.0
V22384 n0_15054_10818 n2_15054_10818 0.0
V22385 n0_15054_11001 n2_15054_11001 0.0
V22386 n0_15054_11034 n2_15054_11034 0.0
V22387 n0_15054_11048 n2_15054_11048 0.0
V22388 n0_15054_11217 n2_15054_11217 0.0
V22389 n0_15054_11250 n2_15054_11250 0.0
V22390 n0_15054_11433 n2_15054_11433 0.0
V22391 n0_15054_11466 n2_15054_11466 0.0
V22392 n0_15054_11865 n2_15054_11865 0.0
V22393 n0_15054_11898 n2_15054_11898 0.0
V22394 n0_15054_12081 n2_15054_12081 0.0
V22395 n0_15054_12114 n2_15054_12114 0.0
V22396 n0_15054_12128 n2_15054_12128 0.0
V22397 n0_15054_12135 n2_15054_12135 0.0
V22398 n0_15054_12297 n2_15054_12297 0.0
V22399 n0_15054_12330 n2_15054_12330 0.0
V22400 n0_15054_12513 n2_15054_12513 0.0
V22401 n0_15054_12546 n2_15054_12546 0.0
V22402 n0_15054_12729 n2_15054_12729 0.0
V22403 n0_15054_12762 n2_15054_12762 0.0
V22404 n0_15054_12776 n2_15054_12776 0.0
V22405 n0_15054_12945 n2_15054_12945 0.0
V22406 n0_15054_12978 n2_15054_12978 0.0
V22407 n0_15054_12992 n2_15054_12992 0.0
V22408 n0_15054_13161 n2_15054_13161 0.0
V22409 n0_15054_13194 n2_15054_13194 0.0
V22410 n0_15054_13377 n2_15054_13377 0.0
V22411 n0_15054_13410 n2_15054_13410 0.0
V22412 n0_15054_13423 n2_15054_13423 0.0
V22413 n0_15054_13593 n2_15054_13593 0.0
V22414 n0_15054_13626 n2_15054_13626 0.0
V22415 n0_15054_13809 n2_15054_13809 0.0
V22416 n0_15054_13842 n2_15054_13842 0.0
V22417 n0_15054_14241 n2_15054_14241 0.0
V22418 n0_15054_14274 n2_15054_14274 0.0
V22419 n0_15054_14457 n2_15054_14457 0.0
V22420 n0_15054_14490 n2_15054_14490 0.0
V22421 n0_15054_14511 n2_15054_14511 0.0
V22422 n0_15054_14673 n2_15054_14673 0.0
V22423 n0_15054_14706 n2_15054_14706 0.0
V22424 n0_15054_14889 n2_15054_14889 0.0
V22425 n0_15054_14922 n2_15054_14922 0.0
V22426 n0_15054_14943 n2_15054_14943 0.0
V22427 n0_15054_15105 n2_15054_15105 0.0
V22428 n0_15054_15138 n2_15054_15138 0.0
V22429 n0_15054_15159 n2_15054_15159 0.0
V22430 n0_15054_15321 n2_15054_15321 0.0
V22431 n0_15054_15354 n2_15054_15354 0.0
V22432 n0_15054_15368 n2_15054_15368 0.0
V22433 n0_15054_15537 n2_15054_15537 0.0
V22434 n0_15054_15570 n2_15054_15570 0.0
V22435 n0_15054_15584 n2_15054_15584 0.0
V22436 n0_15054_15753 n2_15054_15753 0.0
V22437 n0_15054_15786 n2_15054_15786 0.0
V22438 n0_15054_15800 n2_15054_15800 0.0
V22439 n0_15054_15969 n2_15054_15969 0.0
V22440 n0_15054_16002 n2_15054_16002 0.0
V22441 n0_15054_16185 n2_15054_16185 0.0
V22442 n0_15054_16218 n2_15054_16218 0.0
V22443 n0_15054_16401 n2_15054_16401 0.0
V22444 n0_15054_16434 n2_15054_16434 0.0
V22445 n0_15054_16448 n2_15054_16448 0.0
V22446 n0_15054_16617 n2_15054_16617 0.0
V22447 n0_15054_16650 n2_15054_16650 0.0
V22448 n0_15054_16687 n2_15054_16687 0.0
V22449 n0_15054_16833 n2_15054_16833 0.0
V22450 n0_15054_16866 n2_15054_16866 0.0
V22451 n0_15054_17049 n2_15054_17049 0.0
V22452 n0_15054_17082 n2_15054_17082 0.0
V22453 n0_15054_17096 n2_15054_17096 0.0
V22454 n0_15054_17265 n2_15054_17265 0.0
V22455 n0_15054_17298 n2_15054_17298 0.0
V22456 n0_15054_17481 n2_15054_17481 0.0
V22457 n0_15054_17514 n2_15054_17514 0.0
V22458 n0_15054_17528 n2_15054_17528 0.0
V22459 n0_15054_17697 n2_15054_17697 0.0
V22460 n0_15054_17730 n2_15054_17730 0.0
V22461 n0_15054_17913 n2_15054_17913 0.0
V22462 n0_15054_17946 n2_15054_17946 0.0
V22463 n0_15054_17983 n2_15054_17983 0.0
V22464 n0_15054_18129 n2_15054_18129 0.0
V22465 n0_15054_18162 n2_15054_18162 0.0
V22466 n0_15054_18176 n2_15054_18176 0.0
V22467 n0_15054_18345 n2_15054_18345 0.0
V22468 n0_15054_18378 n2_15054_18378 0.0
V22469 n0_15054_18561 n2_15054_18561 0.0
V22470 n0_15054_18594 n2_15054_18594 0.0
V22471 n0_15054_18608 n2_15054_18608 0.0
V22472 n0_15054_18777 n2_15054_18777 0.0
V22473 n0_15054_18810 n2_15054_18810 0.0
V22474 n0_15054_18993 n2_15054_18993 0.0
V22475 n0_15054_19026 n2_15054_19026 0.0
V22476 n0_15054_19209 n2_15054_19209 0.0
V22477 n0_15054_19242 n2_15054_19242 0.0
V22478 n0_15054_19256 n2_15054_19256 0.0
V22479 n0_15054_19263 n2_15054_19263 0.0
V22480 n0_15054_19425 n2_15054_19425 0.0
V22481 n0_15054_19458 n2_15054_19458 0.0
V22482 n0_15054_19641 n2_15054_19641 0.0
V22483 n0_15054_19674 n2_15054_19674 0.0
V22484 n0_15054_19857 n2_15054_19857 0.0
V22485 n0_15054_19890 n2_15054_19890 0.0
V22486 n0_15054_20073 n2_15054_20073 0.0
V22487 n0_15054_20106 n2_15054_20106 0.0
V22488 n0_15054_20289 n2_15054_20289 0.0
V22489 n0_15054_20322 n2_15054_20322 0.0
V22490 n0_15054_20505 n2_15054_20505 0.0
V22491 n0_15054_20538 n2_15054_20538 0.0
V22492 n0_15054_20721 n2_15054_20721 0.0
V22493 n0_15054_20754 n2_15054_20754 0.0
V22494 n0_15054_20937 n2_15054_20937 0.0
V22495 n0_15054_20970 n2_15054_20970 0.0
V22496 n0_15146_201 n2_15146_201 0.0
V22497 n0_15146_234 n2_15146_234 0.0
V22498 n0_15146_417 n2_15146_417 0.0
V22499 n0_15146_450 n2_15146_450 0.0
V22500 n0_15146_633 n2_15146_633 0.0
V22501 n0_15146_666 n2_15146_666 0.0
V22502 n0_15146_849 n2_15146_849 0.0
V22503 n0_15146_882 n2_15146_882 0.0
V22504 n0_15146_1065 n2_15146_1065 0.0
V22505 n0_15146_1098 n2_15146_1098 0.0
V22506 n0_15146_1281 n2_15146_1281 0.0
V22507 n0_15146_1314 n2_15146_1314 0.0
V22508 n0_15146_1497 n2_15146_1497 0.0
V22509 n0_15146_1530 n2_15146_1530 0.0
V22510 n0_15146_1713 n2_15146_1713 0.0
V22511 n0_15146_1746 n2_15146_1746 0.0
V22512 n0_15146_1783 n2_15146_1783 0.0
V22513 n0_15146_1929 n2_15146_1929 0.0
V22514 n0_15146_1962 n2_15146_1962 0.0
V22515 n0_15146_2145 n2_15146_2145 0.0
V22516 n0_15146_2178 n2_15146_2178 0.0
V22517 n0_15146_2361 n2_15146_2361 0.0
V22518 n0_15146_2394 n2_15146_2394 0.0
V22519 n0_15146_2431 n2_15146_2431 0.0
V22520 n0_15146_2577 n2_15146_2577 0.0
V22521 n0_15146_2610 n2_15146_2610 0.0
V22522 n0_15146_2793 n2_15146_2793 0.0
V22523 n0_15146_2826 n2_15146_2826 0.0
V22524 n0_15146_2863 n2_15146_2863 0.0
V22525 n0_15146_3009 n2_15146_3009 0.0
V22526 n0_15146_3042 n2_15146_3042 0.0
V22527 n0_15146_3225 n2_15146_3225 0.0
V22528 n0_15146_3258 n2_15146_3258 0.0
V22529 n0_15146_3295 n2_15146_3295 0.0
V22530 n0_15146_3441 n2_15146_3441 0.0
V22531 n0_15146_3474 n2_15146_3474 0.0
V22532 n0_15146_3511 n2_15146_3511 0.0
V22533 n0_15146_3657 n2_15146_3657 0.0
V22534 n0_15146_3690 n2_15146_3690 0.0
V22535 n0_15146_3873 n2_15146_3873 0.0
V22536 n0_15146_3906 n2_15146_3906 0.0
V22537 n0_15146_3943 n2_15146_3943 0.0
V22538 n0_15146_4089 n2_15146_4089 0.0
V22539 n0_15146_4122 n2_15146_4122 0.0
V22540 n0_15146_4159 n2_15146_4159 0.0
V22541 n0_15146_4305 n2_15146_4305 0.0
V22542 n0_15146_4338 n2_15146_4338 0.0
V22543 n0_15146_4375 n2_15146_4375 0.0
V22544 n0_15146_4521 n2_15146_4521 0.0
V22545 n0_15146_4554 n2_15146_4554 0.0
V22546 n0_15146_4591 n2_15146_4591 0.0
V22547 n0_15146_4737 n2_15146_4737 0.0
V22548 n0_15146_4770 n2_15146_4770 0.0
V22549 n0_15146_4807 n2_15146_4807 0.0
V22550 n0_15146_4953 n2_15146_4953 0.0
V22551 n0_15146_5169 n2_15146_5169 0.0
V22552 n0_15146_5202 n2_15146_5202 0.0
V22553 n0_15146_5239 n2_15146_5239 0.0
V22554 n0_15146_5385 n2_15146_5385 0.0
V22555 n0_15146_5418 n2_15146_5418 0.0
V22556 n0_15146_5455 n2_15146_5455 0.0
V22557 n0_15146_5601 n2_15146_5601 0.0
V22558 n0_15146_5634 n2_15146_5634 0.0
V22559 n0_15146_5671 n2_15146_5671 0.0
V22560 n0_15146_5817 n2_15146_5817 0.0
V22561 n0_15146_5850 n2_15146_5850 0.0
V22562 n0_15146_6033 n2_15146_6033 0.0
V22563 n0_15146_6066 n2_15146_6066 0.0
V22564 n0_15146_15138 n2_15146_15138 0.0
V22565 n0_15146_15159 n2_15146_15159 0.0
V22566 n0_15146_15321 n2_15146_15321 0.0
V22567 n0_15146_15354 n2_15146_15354 0.0
V22568 n0_15146_15368 n2_15146_15368 0.0
V22569 n0_15146_15537 n2_15146_15537 0.0
V22570 n0_15146_15570 n2_15146_15570 0.0
V22571 n0_15146_15584 n2_15146_15584 0.0
V22572 n0_15146_15753 n2_15146_15753 0.0
V22573 n0_15146_15786 n2_15146_15786 0.0
V22574 n0_15146_15800 n2_15146_15800 0.0
V22575 n0_15146_15969 n2_15146_15969 0.0
V22576 n0_15146_16002 n2_15146_16002 0.0
V22577 n0_15146_16185 n2_15146_16185 0.0
V22578 n0_15146_16401 n2_15146_16401 0.0
V22579 n0_15146_16434 n2_15146_16434 0.0
V22580 n0_15146_16448 n2_15146_16448 0.0
V22581 n0_15146_16617 n2_15146_16617 0.0
V22582 n0_15146_16650 n2_15146_16650 0.0
V22583 n0_15146_16687 n2_15146_16687 0.0
V22584 n0_15146_16833 n2_15146_16833 0.0
V22585 n0_15146_16866 n2_15146_16866 0.0
V22586 n0_15146_17049 n2_15146_17049 0.0
V22587 n0_15146_17082 n2_15146_17082 0.0
V22588 n0_15146_17096 n2_15146_17096 0.0
V22589 n0_15146_17265 n2_15146_17265 0.0
V22590 n0_15146_17298 n2_15146_17298 0.0
V22591 n0_15146_17481 n2_15146_17481 0.0
V22592 n0_15146_17514 n2_15146_17514 0.0
V22593 n0_15146_17528 n2_15146_17528 0.0
V22594 n0_15146_17697 n2_15146_17697 0.0
V22595 n0_15146_17730 n2_15146_17730 0.0
V22596 n0_15146_17913 n2_15146_17913 0.0
V22597 n0_15146_17946 n2_15146_17946 0.0
V22598 n0_15146_17983 n2_15146_17983 0.0
V22599 n0_15146_18129 n2_15146_18129 0.0
V22600 n0_15146_18162 n2_15146_18162 0.0
V22601 n0_15146_18176 n2_15146_18176 0.0
V22602 n0_15146_18345 n2_15146_18345 0.0
V22603 n0_15146_18378 n2_15146_18378 0.0
V22604 n0_15146_18561 n2_15146_18561 0.0
V22605 n0_15146_18594 n2_15146_18594 0.0
V22606 n0_15146_18608 n2_15146_18608 0.0
V22607 n0_15146_18777 n2_15146_18777 0.0
V22608 n0_15146_18810 n2_15146_18810 0.0
V22609 n0_15146_18993 n2_15146_18993 0.0
V22610 n0_15146_19026 n2_15146_19026 0.0
V22611 n0_15146_19209 n2_15146_19209 0.0
V22612 n0_15146_19242 n2_15146_19242 0.0
V22613 n0_15146_19256 n2_15146_19256 0.0
V22614 n0_15146_19263 n2_15146_19263 0.0
V22615 n0_15146_19425 n2_15146_19425 0.0
V22616 n0_15146_19458 n2_15146_19458 0.0
V22617 n0_15146_19641 n2_15146_19641 0.0
V22618 n0_15146_19674 n2_15146_19674 0.0
V22619 n0_15146_19857 n2_15146_19857 0.0
V22620 n0_15146_19890 n2_15146_19890 0.0
V22621 n0_15146_20073 n2_15146_20073 0.0
V22622 n0_15146_20106 n2_15146_20106 0.0
V22623 n0_15146_20289 n2_15146_20289 0.0
V22624 n0_15146_20322 n2_15146_20322 0.0
V22625 n0_15146_20505 n2_15146_20505 0.0
V22626 n0_15146_20538 n2_15146_20538 0.0
V22627 n0_15146_20754 n2_15146_20754 0.0
V22628 n0_15146_20937 n2_15146_20937 0.0
V22629 n0_15146_20970 n2_15146_20970 0.0
V22630 n0_15991_5023 n2_15991_5023 0.0
V22631 n0_15991_5169 n2_15991_5169 0.0
V22632 n0_15991_5202 n2_15991_5202 0.0
V22633 n0_15991_5239 n2_15991_5239 0.0
V22634 n0_15991_5385 n2_15991_5385 0.0
V22635 n0_15991_5418 n2_15991_5418 0.0
V22636 n0_15991_5455 n2_15991_5455 0.0
V22637 n0_15991_5601 n2_15991_5601 0.0
V22638 n0_15991_5634 n2_15991_5634 0.0
V22639 n0_15991_5817 n2_15991_5817 0.0
V22640 n0_15991_5850 n2_15991_5850 0.0
V22641 n0_15991_6033 n2_15991_6033 0.0
V22642 n0_15991_6066 n2_15991_6066 0.0
V22643 n0_15991_6249 n2_15991_6249 0.0
V22644 n0_15991_6282 n2_15991_6282 0.0
V22645 n0_15991_6319 n2_15991_6319 0.0
V22646 n0_15991_6465 n2_15991_6465 0.0
V22647 n0_15991_6498 n2_15991_6498 0.0
V22648 n0_15991_6681 n2_15991_6681 0.0
V22649 n0_15991_6714 n2_15991_6714 0.0
V22650 n0_15991_6897 n2_15991_6897 0.0
V22651 n0_15991_6930 n2_15991_6930 0.0
V22652 n0_15991_7113 n2_15991_7113 0.0
V22653 n0_15991_7146 n2_15991_7146 0.0
V22654 n0_15991_7329 n2_15991_7329 0.0
V22655 n0_15991_7362 n2_15991_7362 0.0
V22656 n0_15991_7545 n2_15991_7545 0.0
V22657 n0_15991_7578 n2_15991_7578 0.0
V22658 n0_15991_7761 n2_15991_7761 0.0
V22659 n0_15991_7794 n2_15991_7794 0.0
V22660 n0_15991_7831 n2_15991_7831 0.0
V22661 n0_15991_7977 n2_15991_7977 0.0
V22662 n0_15991_8010 n2_15991_8010 0.0
V22663 n0_15991_8193 n2_15991_8193 0.0
V22664 n0_15991_8226 n2_15991_8226 0.0
V22665 n0_15991_8409 n2_15991_8409 0.0
V22666 n0_15991_8442 n2_15991_8442 0.0
V22667 n0_15991_8625 n2_15991_8625 0.0
V22668 n0_15991_8658 n2_15991_8658 0.0
V22669 n0_15991_8841 n2_15991_8841 0.0
V22670 n0_15991_8874 n2_15991_8874 0.0
V22671 n0_15991_8911 n2_15991_8911 0.0
V22672 n0_15991_9057 n2_15991_9057 0.0
V22673 n0_15991_9090 n2_15991_9090 0.0
V22674 n0_15991_9273 n2_15991_9273 0.0
V22675 n0_15991_9306 n2_15991_9306 0.0
V22676 n0_15991_9489 n2_15991_9489 0.0
V22677 n0_15991_9522 n2_15991_9522 0.0
V22678 n0_15991_9705 n2_15991_9705 0.0
V22679 n0_15991_9738 n2_15991_9738 0.0
V22680 n0_15991_9921 n2_15991_9921 0.0
V22681 n0_15991_9954 n2_15991_9954 0.0
V22682 n0_15991_9991 n2_15991_9991 0.0
V22683 n0_15991_10137 n2_15991_10137 0.0
V22684 n0_15991_10170 n2_15991_10170 0.0
V22685 n0_15991_10353 n2_15991_10353 0.0
V22686 n0_15991_10386 n2_15991_10386 0.0
V22687 n0_15991_10569 n2_15991_10569 0.0
V22688 n0_15991_10785 n2_15991_10785 0.0
V22689 n0_15991_10818 n2_15991_10818 0.0
V22690 n0_15991_11001 n2_15991_11001 0.0
V22691 n0_15991_11034 n2_15991_11034 0.0
V22692 n0_15991_11048 n2_15991_11048 0.0
V22693 n0_15991_11217 n2_15991_11217 0.0
V22694 n0_15991_11250 n2_15991_11250 0.0
V22695 n0_15991_11433 n2_15991_11433 0.0
V22696 n0_15991_11466 n2_15991_11466 0.0
V22697 n0_15991_11649 n2_15991_11649 0.0
V22698 n0_15991_11682 n2_15991_11682 0.0
V22699 n0_15991_11865 n2_15991_11865 0.0
V22700 n0_15991_11898 n2_15991_11898 0.0
V22701 n0_15991_12081 n2_15991_12081 0.0
V22702 n0_15991_12114 n2_15991_12114 0.0
V22703 n0_15991_12128 n2_15991_12128 0.0
V22704 n0_15991_12135 n2_15991_12135 0.0
V22705 n0_15991_12297 n2_15991_12297 0.0
V22706 n0_15991_12330 n2_15991_12330 0.0
V22707 n0_15991_12513 n2_15991_12513 0.0
V22708 n0_15991_12546 n2_15991_12546 0.0
V22709 n0_15991_12729 n2_15991_12729 0.0
V22710 n0_15991_12762 n2_15991_12762 0.0
V22711 n0_15991_12776 n2_15991_12776 0.0
V22712 n0_15991_12945 n2_15991_12945 0.0
V22713 n0_15991_12978 n2_15991_12978 0.0
V22714 n0_15991_12992 n2_15991_12992 0.0
V22715 n0_15991_13161 n2_15991_13161 0.0
V22716 n0_15991_13194 n2_15991_13194 0.0
V22717 n0_15991_13377 n2_15991_13377 0.0
V22718 n0_15991_13410 n2_15991_13410 0.0
V22719 n0_15991_13423 n2_15991_13423 0.0
V22720 n0_15991_13593 n2_15991_13593 0.0
V22721 n0_15991_13626 n2_15991_13626 0.0
V22722 n0_15991_13647 n2_15991_13647 0.0
V22723 n0_15991_13809 n2_15991_13809 0.0
V22724 n0_15991_13842 n2_15991_13842 0.0
V22725 n0_15991_14025 n2_15991_14025 0.0
V22726 n0_15991_14058 n2_15991_14058 0.0
V22727 n0_15991_14241 n2_15991_14241 0.0
V22728 n0_15991_14274 n2_15991_14274 0.0
V22729 n0_15991_14457 n2_15991_14457 0.0
V22730 n0_15991_14490 n2_15991_14490 0.0
V22731 n0_15991_14511 n2_15991_14511 0.0
V22732 n0_15991_14673 n2_15991_14673 0.0
V22733 n0_15991_14706 n2_15991_14706 0.0
V22734 n0_15991_14889 n2_15991_14889 0.0
V22735 n0_15991_14922 n2_15991_14922 0.0
V22736 n0_15991_14943 n2_15991_14943 0.0
V22737 n0_15991_15138 n2_15991_15138 0.0
V22738 n0_15991_15159 n2_15991_15159 0.0
V22739 n0_15991_15321 n2_15991_15321 0.0
V22740 n0_15991_15354 n2_15991_15354 0.0
V22741 n0_15991_15537 n2_15991_15537 0.0
V22742 n0_15991_15570 n2_15991_15570 0.0
V22743 n0_15991_15584 n2_15991_15584 0.0
V22744 n0_15991_15753 n2_15991_15753 0.0
V22745 n0_15991_15786 n2_15991_15786 0.0
V22746 n0_15991_15969 n2_15991_15969 0.0
V22747 n0_15991_16002 n2_15991_16002 0.0
V22748 n0_15991_16185 n2_15991_16185 0.0
V22749 n0_16130_6033 n2_16130_6033 0.0
V22750 n0_16130_6066 n2_16130_6066 0.0
V22751 n0_16130_8409 n2_16130_8409 0.0
V22752 n0_16130_10569 n2_16130_10569 0.0
V22753 n0_16130_10602 n2_16130_10602 0.0
V22754 n0_16130_12776 n2_16130_12776 0.0
V22755 n0_16130_15105 n2_16130_15105 0.0
V22756 n0_16130_15138 n2_16130_15138 0.0
V22757 n0_16130_15159 n2_16130_15159 0.0
V22758 n0_16179_5169 n2_16179_5169 0.0
V22759 n0_16179_5202 n2_16179_5202 0.0
V22760 n0_16179_5239 n2_16179_5239 0.0
V22761 n0_16179_5385 n2_16179_5385 0.0
V22762 n0_16179_5418 n2_16179_5418 0.0
V22763 n0_16179_5455 n2_16179_5455 0.0
V22764 n0_16179_5601 n2_16179_5601 0.0
V22765 n0_16179_5634 n2_16179_5634 0.0
V22766 n0_16179_5817 n2_16179_5817 0.0
V22767 n0_16179_5850 n2_16179_5850 0.0
V22768 n0_16179_6033 n2_16179_6033 0.0
V22769 n0_16179_6066 n2_16179_6066 0.0
V22770 n0_16179_6249 n2_16179_6249 0.0
V22771 n0_16179_6282 n2_16179_6282 0.0
V22772 n0_16179_6319 n2_16179_6319 0.0
V22773 n0_16179_6465 n2_16179_6465 0.0
V22774 n0_16179_6498 n2_16179_6498 0.0
V22775 n0_16179_6681 n2_16179_6681 0.0
V22776 n0_16179_6714 n2_16179_6714 0.0
V22777 n0_16179_6897 n2_16179_6897 0.0
V22778 n0_16179_6930 n2_16179_6930 0.0
V22779 n0_16179_7113 n2_16179_7113 0.0
V22780 n0_16179_7329 n2_16179_7329 0.0
V22781 n0_16179_7362 n2_16179_7362 0.0
V22782 n0_16179_7545 n2_16179_7545 0.0
V22783 n0_16179_7578 n2_16179_7578 0.0
V22784 n0_16179_7761 n2_16179_7761 0.0
V22785 n0_16179_7794 n2_16179_7794 0.0
V22786 n0_16179_7831 n2_16179_7831 0.0
V22787 n0_16179_7977 n2_16179_7977 0.0
V22788 n0_16179_8010 n2_16179_8010 0.0
V22789 n0_16179_8193 n2_16179_8193 0.0
V22790 n0_16179_8226 n2_16179_8226 0.0
V22791 n0_16179_8409 n2_16179_8409 0.0
V22792 n0_16179_8442 n2_16179_8442 0.0
V22793 n0_16179_8625 n2_16179_8625 0.0
V22794 n0_16179_8658 n2_16179_8658 0.0
V22795 n0_16179_8841 n2_16179_8841 0.0
V22796 n0_16179_8874 n2_16179_8874 0.0
V22797 n0_16179_8911 n2_16179_8911 0.0
V22798 n0_16179_9057 n2_16179_9057 0.0
V22799 n0_16179_9090 n2_16179_9090 0.0
V22800 n0_16179_9273 n2_16179_9273 0.0
V22801 n0_16179_9306 n2_16179_9306 0.0
V22802 n0_16179_9705 n2_16179_9705 0.0
V22803 n0_16179_9738 n2_16179_9738 0.0
V22804 n0_16179_9921 n2_16179_9921 0.0
V22805 n0_16179_9954 n2_16179_9954 0.0
V22806 n0_16179_9991 n2_16179_9991 0.0
V22807 n0_16179_10137 n2_16179_10137 0.0
V22808 n0_16179_10170 n2_16179_10170 0.0
V22809 n0_16179_10353 n2_16179_10353 0.0
V22810 n0_16179_10386 n2_16179_10386 0.0
V22811 n0_16179_10569 n2_16179_10569 0.0
V22812 n0_16179_10602 n2_16179_10602 0.0
V22813 n0_16179_10785 n2_16179_10785 0.0
V22814 n0_16179_10818 n2_16179_10818 0.0
V22815 n0_16179_11001 n2_16179_11001 0.0
V22816 n0_16179_11034 n2_16179_11034 0.0
V22817 n0_16179_11048 n2_16179_11048 0.0
V22818 n0_16179_11217 n2_16179_11217 0.0
V22819 n0_16179_11250 n2_16179_11250 0.0
V22820 n0_16179_11433 n2_16179_11433 0.0
V22821 n0_16179_11466 n2_16179_11466 0.0
V22822 n0_16179_11865 n2_16179_11865 0.0
V22823 n0_16179_11898 n2_16179_11898 0.0
V22824 n0_16179_12081 n2_16179_12081 0.0
V22825 n0_16179_12114 n2_16179_12114 0.0
V22826 n0_16179_12128 n2_16179_12128 0.0
V22827 n0_16179_12135 n2_16179_12135 0.0
V22828 n0_16179_12297 n2_16179_12297 0.0
V22829 n0_16179_12330 n2_16179_12330 0.0
V22830 n0_16179_12513 n2_16179_12513 0.0
V22831 n0_16179_12546 n2_16179_12546 0.0
V22832 n0_16179_12729 n2_16179_12729 0.0
V22833 n0_16179_12762 n2_16179_12762 0.0
V22834 n0_16179_12776 n2_16179_12776 0.0
V22835 n0_16179_12945 n2_16179_12945 0.0
V22836 n0_16179_12978 n2_16179_12978 0.0
V22837 n0_16179_12992 n2_16179_12992 0.0
V22838 n0_16179_13161 n2_16179_13161 0.0
V22839 n0_16179_13194 n2_16179_13194 0.0
V22840 n0_16179_13377 n2_16179_13377 0.0
V22841 n0_16179_13410 n2_16179_13410 0.0
V22842 n0_16179_13423 n2_16179_13423 0.0
V22843 n0_16179_13593 n2_16179_13593 0.0
V22844 n0_16179_13626 n2_16179_13626 0.0
V22845 n0_16179_13647 n2_16179_13647 0.0
V22846 n0_16179_13809 n2_16179_13809 0.0
V22847 n0_16179_13842 n2_16179_13842 0.0
V22848 n0_16179_14241 n2_16179_14241 0.0
V22849 n0_16179_14274 n2_16179_14274 0.0
V22850 n0_16179_14457 n2_16179_14457 0.0
V22851 n0_16179_14490 n2_16179_14490 0.0
V22852 n0_16179_14511 n2_16179_14511 0.0
V22853 n0_16179_14673 n2_16179_14673 0.0
V22854 n0_16179_14706 n2_16179_14706 0.0
V22855 n0_16179_14889 n2_16179_14889 0.0
V22856 n0_16179_14922 n2_16179_14922 0.0
V22857 n0_16179_14943 n2_16179_14943 0.0
V22858 n0_16179_15105 n2_16179_15105 0.0
V22859 n0_16179_15138 n2_16179_15138 0.0
V22860 n0_16179_15159 n2_16179_15159 0.0
V22861 n0_16179_15321 n2_16179_15321 0.0
V22862 n0_16179_15354 n2_16179_15354 0.0
V22863 n0_16179_15537 n2_16179_15537 0.0
V22864 n0_16179_15570 n2_16179_15570 0.0
V22865 n0_16179_15584 n2_16179_15584 0.0
V22866 n0_16179_15753 n2_16179_15753 0.0
V22867 n0_16179_15786 n2_16179_15786 0.0
V22868 n0_16179_15969 n2_16179_15969 0.0
V22869 n0_16179_16002 n2_16179_16002 0.0
V22870 n0_17116_201 n2_17116_201 0.0
V22871 n0_17116_234 n2_17116_234 0.0
V22872 n0_17116_417 n2_17116_417 0.0
V22873 n0_17116_450 n2_17116_450 0.0
V22874 n0_17116_633 n2_17116_633 0.0
V22875 n0_17116_666 n2_17116_666 0.0
V22876 n0_17116_849 n2_17116_849 0.0
V22877 n0_17116_882 n2_17116_882 0.0
V22878 n0_17116_1065 n2_17116_1065 0.0
V22879 n0_17116_1098 n2_17116_1098 0.0
V22880 n0_17116_1281 n2_17116_1281 0.0
V22881 n0_17116_1314 n2_17116_1314 0.0
V22882 n0_17116_1497 n2_17116_1497 0.0
V22883 n0_17116_1530 n2_17116_1530 0.0
V22884 n0_17116_1713 n2_17116_1713 0.0
V22885 n0_17116_1746 n2_17116_1746 0.0
V22886 n0_17116_1783 n2_17116_1783 0.0
V22887 n0_17116_1929 n2_17116_1929 0.0
V22888 n0_17116_1962 n2_17116_1962 0.0
V22889 n0_17116_2145 n2_17116_2145 0.0
V22890 n0_17116_2178 n2_17116_2178 0.0
V22891 n0_17116_2361 n2_17116_2361 0.0
V22892 n0_17116_2394 n2_17116_2394 0.0
V22893 n0_17116_2431 n2_17116_2431 0.0
V22894 n0_17116_2577 n2_17116_2577 0.0
V22895 n0_17116_2610 n2_17116_2610 0.0
V22896 n0_17116_2793 n2_17116_2793 0.0
V22897 n0_17116_2826 n2_17116_2826 0.0
V22898 n0_17116_2863 n2_17116_2863 0.0
V22899 n0_17116_3009 n2_17116_3009 0.0
V22900 n0_17116_3042 n2_17116_3042 0.0
V22901 n0_17116_3225 n2_17116_3225 0.0
V22902 n0_17116_3258 n2_17116_3258 0.0
V22903 n0_17116_3295 n2_17116_3295 0.0
V22904 n0_17116_3441 n2_17116_3441 0.0
V22905 n0_17116_3474 n2_17116_3474 0.0
V22906 n0_17116_3657 n2_17116_3657 0.0
V22907 n0_17116_3690 n2_17116_3690 0.0
V22908 n0_17116_3873 n2_17116_3873 0.0
V22909 n0_17116_3906 n2_17116_3906 0.0
V22910 n0_17116_4089 n2_17116_4089 0.0
V22911 n0_17116_4122 n2_17116_4122 0.0
V22912 n0_17116_4305 n2_17116_4305 0.0
V22913 n0_17116_4338 n2_17116_4338 0.0
V22914 n0_17116_4375 n2_17116_4375 0.0
V22915 n0_17116_4521 n2_17116_4521 0.0
V22916 n0_17116_4554 n2_17116_4554 0.0
V22917 n0_17116_4591 n2_17116_4591 0.0
V22918 n0_17116_4737 n2_17116_4737 0.0
V22919 n0_17116_4770 n2_17116_4770 0.0
V22920 n0_17116_4807 n2_17116_4807 0.0
V22921 n0_17116_4953 n2_17116_4953 0.0
V22922 n0_17116_4986 n2_17116_4986 0.0
V22923 n0_17116_5023 n2_17116_5023 0.0
V22924 n0_17116_5169 n2_17116_5169 0.0
V22925 n0_17116_5202 n2_17116_5202 0.0
V22926 n0_17116_5239 n2_17116_5239 0.0
V22927 n0_17116_5385 n2_17116_5385 0.0
V22928 n0_17116_5418 n2_17116_5418 0.0
V22929 n0_17116_5455 n2_17116_5455 0.0
V22930 n0_17116_5601 n2_17116_5601 0.0
V22931 n0_17116_5634 n2_17116_5634 0.0
V22932 n0_17116_5817 n2_17116_5817 0.0
V22933 n0_17116_5850 n2_17116_5850 0.0
V22934 n0_17116_6033 n2_17116_6033 0.0
V22935 n0_17116_6066 n2_17116_6066 0.0
V22936 n0_17116_6249 n2_17116_6249 0.0
V22937 n0_17116_6282 n2_17116_6282 0.0
V22938 n0_17116_6319 n2_17116_6319 0.0
V22939 n0_17116_6465 n2_17116_6465 0.0
V22940 n0_17116_6498 n2_17116_6498 0.0
V22941 n0_17116_6681 n2_17116_6681 0.0
V22942 n0_17116_6714 n2_17116_6714 0.0
V22943 n0_17116_6897 n2_17116_6897 0.0
V22944 n0_17116_6930 n2_17116_6930 0.0
V22945 n0_17116_7113 n2_17116_7113 0.0
V22946 n0_17116_7146 n2_17116_7146 0.0
V22947 n0_17116_7329 n2_17116_7329 0.0
V22948 n0_17116_7362 n2_17116_7362 0.0
V22949 n0_17116_7545 n2_17116_7545 0.0
V22950 n0_17116_7578 n2_17116_7578 0.0
V22951 n0_17116_7761 n2_17116_7761 0.0
V22952 n0_17116_7794 n2_17116_7794 0.0
V22953 n0_17116_7831 n2_17116_7831 0.0
V22954 n0_17116_7977 n2_17116_7977 0.0
V22955 n0_17116_8010 n2_17116_8010 0.0
V22956 n0_17116_8193 n2_17116_8193 0.0
V22957 n0_17116_8226 n2_17116_8226 0.0
V22958 n0_17116_8409 n2_17116_8409 0.0
V22959 n0_17116_8442 n2_17116_8442 0.0
V22960 n0_17116_8625 n2_17116_8625 0.0
V22961 n0_17116_8658 n2_17116_8658 0.0
V22962 n0_17116_8841 n2_17116_8841 0.0
V22963 n0_17116_8874 n2_17116_8874 0.0
V22964 n0_17116_8911 n2_17116_8911 0.0
V22965 n0_17116_9057 n2_17116_9057 0.0
V22966 n0_17116_9090 n2_17116_9090 0.0
V22967 n0_17116_9273 n2_17116_9273 0.0
V22968 n0_17116_9306 n2_17116_9306 0.0
V22969 n0_17116_9489 n2_17116_9489 0.0
V22970 n0_17116_9522 n2_17116_9522 0.0
V22971 n0_17116_9705 n2_17116_9705 0.0
V22972 n0_17116_9738 n2_17116_9738 0.0
V22973 n0_17116_9921 n2_17116_9921 0.0
V22974 n0_17116_9954 n2_17116_9954 0.0
V22975 n0_17116_9991 n2_17116_9991 0.0
V22976 n0_17116_10137 n2_17116_10137 0.0
V22977 n0_17116_10170 n2_17116_10170 0.0
V22978 n0_17116_10353 n2_17116_10353 0.0
V22979 n0_17116_10386 n2_17116_10386 0.0
V22980 n0_17116_10569 n2_17116_10569 0.0
V22981 n0_17116_10785 n2_17116_10785 0.0
V22982 n0_17116_10818 n2_17116_10818 0.0
V22983 n0_17116_11001 n2_17116_11001 0.0
V22984 n0_17116_11034 n2_17116_11034 0.0
V22985 n0_17116_11048 n2_17116_11048 0.0
V22986 n0_17116_11055 n2_17116_11055 0.0
V22987 n0_17116_11217 n2_17116_11217 0.0
V22988 n0_17116_11250 n2_17116_11250 0.0
V22989 n0_17116_11433 n2_17116_11433 0.0
V22990 n0_17116_11466 n2_17116_11466 0.0
V22991 n0_17116_11649 n2_17116_11649 0.0
V22992 n0_17116_11682 n2_17116_11682 0.0
V22993 n0_17116_11865 n2_17116_11865 0.0
V22994 n0_17116_11898 n2_17116_11898 0.0
V22995 n0_17116_12081 n2_17116_12081 0.0
V22996 n0_17116_12114 n2_17116_12114 0.0
V22997 n0_17116_12128 n2_17116_12128 0.0
V22998 n0_17116_12135 n2_17116_12135 0.0
V22999 n0_17116_12297 n2_17116_12297 0.0
V23000 n0_17116_12330 n2_17116_12330 0.0
V23001 n0_17116_12513 n2_17116_12513 0.0
V23002 n0_17116_12546 n2_17116_12546 0.0
V23003 n0_17116_12729 n2_17116_12729 0.0
V23004 n0_17116_12762 n2_17116_12762 0.0
V23005 n0_17116_12945 n2_17116_12945 0.0
V23006 n0_17116_12978 n2_17116_12978 0.0
V23007 n0_17116_13161 n2_17116_13161 0.0
V23008 n0_17116_13194 n2_17116_13194 0.0
V23009 n0_17116_13377 n2_17116_13377 0.0
V23010 n0_17116_13410 n2_17116_13410 0.0
V23011 n0_17116_13593 n2_17116_13593 0.0
V23012 n0_17116_13626 n2_17116_13626 0.0
V23013 n0_17116_13640 n2_17116_13640 0.0
V23014 n0_17116_13647 n2_17116_13647 0.0
V23015 n0_17116_13809 n2_17116_13809 0.0
V23016 n0_17116_13842 n2_17116_13842 0.0
V23017 n0_17116_14025 n2_17116_14025 0.0
V23018 n0_17116_14058 n2_17116_14058 0.0
V23019 n0_17116_14241 n2_17116_14241 0.0
V23020 n0_17116_14274 n2_17116_14274 0.0
V23021 n0_17116_14457 n2_17116_14457 0.0
V23022 n0_17116_14490 n2_17116_14490 0.0
V23023 n0_17116_14511 n2_17116_14511 0.0
V23024 n0_17116_14673 n2_17116_14673 0.0
V23025 n0_17116_14706 n2_17116_14706 0.0
V23026 n0_17116_14889 n2_17116_14889 0.0
V23027 n0_17116_14922 n2_17116_14922 0.0
V23028 n0_17116_14936 n2_17116_14936 0.0
V23029 n0_17116_14943 n2_17116_14943 0.0
V23030 n0_17116_15138 n2_17116_15138 0.0
V23031 n0_17116_15152 n2_17116_15152 0.0
V23032 n0_17116_15159 n2_17116_15159 0.0
V23033 n0_17116_15321 n2_17116_15321 0.0
V23034 n0_17116_15354 n2_17116_15354 0.0
V23035 n0_17116_15537 n2_17116_15537 0.0
V23036 n0_17116_15570 n2_17116_15570 0.0
V23037 n0_17116_15584 n2_17116_15584 0.0
V23038 n0_17116_15753 n2_17116_15753 0.0
V23039 n0_17116_15786 n2_17116_15786 0.0
V23040 n0_17116_15969 n2_17116_15969 0.0
V23041 n0_17116_16002 n2_17116_16002 0.0
V23042 n0_17116_16185 n2_17116_16185 0.0
V23043 n0_17116_16218 n2_17116_16218 0.0
V23044 n0_17116_16401 n2_17116_16401 0.0
V23045 n0_17116_16434 n2_17116_16434 0.0
V23046 n0_17116_16617 n2_17116_16617 0.0
V23047 n0_17116_16650 n2_17116_16650 0.0
V23048 n0_17116_16664 n2_17116_16664 0.0
V23049 n0_17116_16687 n2_17116_16687 0.0
V23050 n0_17116_16833 n2_17116_16833 0.0
V23051 n0_17116_16866 n2_17116_16866 0.0
V23052 n0_17116_17049 n2_17116_17049 0.0
V23053 n0_17116_17082 n2_17116_17082 0.0
V23054 n0_17116_17119 n2_17116_17119 0.0
V23055 n0_17116_17265 n2_17116_17265 0.0
V23056 n0_17116_17298 n2_17116_17298 0.0
V23057 n0_17116_17481 n2_17116_17481 0.0
V23058 n0_17116_17514 n2_17116_17514 0.0
V23059 n0_17116_17535 n2_17116_17535 0.0
V23060 n0_17116_17697 n2_17116_17697 0.0
V23061 n0_17116_17730 n2_17116_17730 0.0
V23062 n0_17116_17913 n2_17116_17913 0.0
V23063 n0_17116_17946 n2_17116_17946 0.0
V23064 n0_17116_18129 n2_17116_18129 0.0
V23065 n0_17116_18162 n2_17116_18162 0.0
V23066 n0_17116_18176 n2_17116_18176 0.0
V23067 n0_17116_18345 n2_17116_18345 0.0
V23068 n0_17116_18378 n2_17116_18378 0.0
V23069 n0_17116_18561 n2_17116_18561 0.0
V23070 n0_17116_18594 n2_17116_18594 0.0
V23071 n0_17116_18777 n2_17116_18777 0.0
V23072 n0_17116_18810 n2_17116_18810 0.0
V23073 n0_17116_18993 n2_17116_18993 0.0
V23074 n0_17116_19026 n2_17116_19026 0.0
V23075 n0_17116_19040 n2_17116_19040 0.0
V23076 n0_17116_19209 n2_17116_19209 0.0
V23077 n0_17116_19242 n2_17116_19242 0.0
V23078 n0_17116_19425 n2_17116_19425 0.0
V23079 n0_17116_19458 n2_17116_19458 0.0
V23080 n0_17116_19641 n2_17116_19641 0.0
V23081 n0_17116_19674 n2_17116_19674 0.0
V23082 n0_17116_19857 n2_17116_19857 0.0
V23083 n0_17116_19890 n2_17116_19890 0.0
V23084 n0_17116_20073 n2_17116_20073 0.0
V23085 n0_17116_20106 n2_17116_20106 0.0
V23086 n0_17116_20289 n2_17116_20289 0.0
V23087 n0_17116_20322 n2_17116_20322 0.0
V23088 n0_17116_20505 n2_17116_20505 0.0
V23089 n0_17116_20538 n2_17116_20538 0.0
V23090 n0_17116_20754 n2_17116_20754 0.0
V23091 n0_17116_20937 n2_17116_20937 0.0
V23092 n0_17116_20970 n2_17116_20970 0.0
V23093 n0_17208_201 n2_17208_201 0.0
V23094 n0_17208_234 n2_17208_234 0.0
V23095 n0_17208_417 n2_17208_417 0.0
V23096 n0_17208_450 n2_17208_450 0.0
V23097 n0_17208_633 n2_17208_633 0.0
V23098 n0_17208_666 n2_17208_666 0.0
V23099 n0_17208_849 n2_17208_849 0.0
V23100 n0_17208_882 n2_17208_882 0.0
V23101 n0_17208_1065 n2_17208_1065 0.0
V23102 n0_17208_1098 n2_17208_1098 0.0
V23103 n0_17208_1281 n2_17208_1281 0.0
V23104 n0_17208_1314 n2_17208_1314 0.0
V23105 n0_17208_1497 n2_17208_1497 0.0
V23106 n0_17208_1530 n2_17208_1530 0.0
V23107 n0_17208_1713 n2_17208_1713 0.0
V23108 n0_17208_1746 n2_17208_1746 0.0
V23109 n0_17208_1783 n2_17208_1783 0.0
V23110 n0_17208_1929 n2_17208_1929 0.0
V23111 n0_17208_1962 n2_17208_1962 0.0
V23112 n0_17208_2145 n2_17208_2145 0.0
V23113 n0_17208_2178 n2_17208_2178 0.0
V23114 n0_17208_2361 n2_17208_2361 0.0
V23115 n0_17208_2394 n2_17208_2394 0.0
V23116 n0_17208_2431 n2_17208_2431 0.0
V23117 n0_17208_2577 n2_17208_2577 0.0
V23118 n0_17208_2610 n2_17208_2610 0.0
V23119 n0_17208_2793 n2_17208_2793 0.0
V23120 n0_17208_2826 n2_17208_2826 0.0
V23121 n0_17208_2863 n2_17208_2863 0.0
V23122 n0_17208_3009 n2_17208_3009 0.0
V23123 n0_17208_3042 n2_17208_3042 0.0
V23124 n0_17208_3225 n2_17208_3225 0.0
V23125 n0_17208_3258 n2_17208_3258 0.0
V23126 n0_17208_3295 n2_17208_3295 0.0
V23127 n0_17208_3441 n2_17208_3441 0.0
V23128 n0_17208_3474 n2_17208_3474 0.0
V23129 n0_17208_3657 n2_17208_3657 0.0
V23130 n0_17208_3690 n2_17208_3690 0.0
V23131 n0_17208_3873 n2_17208_3873 0.0
V23132 n0_17208_3906 n2_17208_3906 0.0
V23133 n0_17208_17265 n2_17208_17265 0.0
V23134 n0_17208_17298 n2_17208_17298 0.0
V23135 n0_17208_17481 n2_17208_17481 0.0
V23136 n0_17208_17514 n2_17208_17514 0.0
V23137 n0_17208_17535 n2_17208_17535 0.0
V23138 n0_17208_17697 n2_17208_17697 0.0
V23139 n0_17208_17730 n2_17208_17730 0.0
V23140 n0_17208_17913 n2_17208_17913 0.0
V23141 n0_17208_17946 n2_17208_17946 0.0
V23142 n0_17208_18129 n2_17208_18129 0.0
V23143 n0_17208_18162 n2_17208_18162 0.0
V23144 n0_17208_18176 n2_17208_18176 0.0
V23145 n0_17208_18345 n2_17208_18345 0.0
V23146 n0_17208_18378 n2_17208_18378 0.0
V23147 n0_17208_18561 n2_17208_18561 0.0
V23148 n0_17208_18594 n2_17208_18594 0.0
V23149 n0_17208_18777 n2_17208_18777 0.0
V23150 n0_17208_18810 n2_17208_18810 0.0
V23151 n0_17208_18993 n2_17208_18993 0.0
V23152 n0_17208_19026 n2_17208_19026 0.0
V23153 n0_17208_19040 n2_17208_19040 0.0
V23154 n0_17208_19209 n2_17208_19209 0.0
V23155 n0_17208_19242 n2_17208_19242 0.0
V23156 n0_17208_19425 n2_17208_19425 0.0
V23157 n0_17208_19458 n2_17208_19458 0.0
V23158 n0_17208_19641 n2_17208_19641 0.0
V23159 n0_17208_19674 n2_17208_19674 0.0
V23160 n0_17208_19857 n2_17208_19857 0.0
V23161 n0_17208_19890 n2_17208_19890 0.0
V23162 n0_17208_20073 n2_17208_20073 0.0
V23163 n0_17208_20106 n2_17208_20106 0.0
V23164 n0_17208_20289 n2_17208_20289 0.0
V23165 n0_17208_20322 n2_17208_20322 0.0
V23166 n0_17208_20505 n2_17208_20505 0.0
V23167 n0_17208_20538 n2_17208_20538 0.0
V23168 n0_17208_20721 n2_17208_20721 0.0
V23169 n0_17208_20754 n2_17208_20754 0.0
V23170 n0_17208_20937 n2_17208_20937 0.0
V23171 n0_17208_20970 n2_17208_20970 0.0
V23172 n0_17255_417 n2_17255_417 0.0
V23173 n0_17255_450 n2_17255_450 0.0
V23174 n0_17255_1530 n2_17255_1530 0.0
V23175 n0_17255_2793 n2_17255_2793 0.0
V23176 n0_17255_3873 n2_17255_3873 0.0
V23177 n0_17255_3906 n2_17255_3906 0.0
V23178 n0_17255_6033 n2_17255_6033 0.0
V23179 n0_17255_6066 n2_17255_6066 0.0
V23180 n0_17255_8409 n2_17255_8409 0.0
V23181 n0_17255_10569 n2_17255_10569 0.0
V23182 n0_17255_10602 n2_17255_10602 0.0
V23183 n0_17255_15105 n2_17255_15105 0.0
V23184 n0_17255_15138 n2_17255_15138 0.0
V23185 n0_17255_15152 n2_17255_15152 0.0
V23186 n0_17255_15159 n2_17255_15159 0.0
V23187 n0_17255_17298 n2_17255_17298 0.0
V23188 n0_17255_19641 n2_17255_19641 0.0
V23189 n0_17255_19674 n2_17255_19674 0.0
V23190 n0_17255_20721 n2_17255_20721 0.0
V23191 n0_17255_20754 n2_17255_20754 0.0
V23192 n0_17304_201 n2_17304_201 0.0
V23193 n0_17304_234 n2_17304_234 0.0
V23194 n0_17304_417 n2_17304_417 0.0
V23195 n0_17304_450 n2_17304_450 0.0
V23196 n0_17304_633 n2_17304_633 0.0
V23197 n0_17304_666 n2_17304_666 0.0
V23198 n0_17304_849 n2_17304_849 0.0
V23199 n0_17304_882 n2_17304_882 0.0
V23200 n0_17304_1065 n2_17304_1065 0.0
V23201 n0_17304_1098 n2_17304_1098 0.0
V23202 n0_17304_1281 n2_17304_1281 0.0
V23203 n0_17304_1314 n2_17304_1314 0.0
V23204 n0_17304_1497 n2_17304_1497 0.0
V23205 n0_17304_1530 n2_17304_1530 0.0
V23206 n0_17304_1713 n2_17304_1713 0.0
V23207 n0_17304_1746 n2_17304_1746 0.0
V23208 n0_17304_1783 n2_17304_1783 0.0
V23209 n0_17304_1929 n2_17304_1929 0.0
V23210 n0_17304_1962 n2_17304_1962 0.0
V23211 n0_17304_2145 n2_17304_2145 0.0
V23212 n0_17304_2178 n2_17304_2178 0.0
V23213 n0_17304_2361 n2_17304_2361 0.0
V23214 n0_17304_2394 n2_17304_2394 0.0
V23215 n0_17304_2431 n2_17304_2431 0.0
V23216 n0_17304_2577 n2_17304_2577 0.0
V23217 n0_17304_2610 n2_17304_2610 0.0
V23218 n0_17304_2793 n2_17304_2793 0.0
V23219 n0_17304_2826 n2_17304_2826 0.0
V23220 n0_17304_2863 n2_17304_2863 0.0
V23221 n0_17304_3009 n2_17304_3009 0.0
V23222 n0_17304_3042 n2_17304_3042 0.0
V23223 n0_17304_3225 n2_17304_3225 0.0
V23224 n0_17304_3258 n2_17304_3258 0.0
V23225 n0_17304_3295 n2_17304_3295 0.0
V23226 n0_17304_3441 n2_17304_3441 0.0
V23227 n0_17304_3474 n2_17304_3474 0.0
V23228 n0_17304_3657 n2_17304_3657 0.0
V23229 n0_17304_3690 n2_17304_3690 0.0
V23230 n0_17304_3873 n2_17304_3873 0.0
V23231 n0_17304_3906 n2_17304_3906 0.0
V23232 n0_17304_4089 n2_17304_4089 0.0
V23233 n0_17304_4122 n2_17304_4122 0.0
V23234 n0_17304_4305 n2_17304_4305 0.0
V23235 n0_17304_4338 n2_17304_4338 0.0
V23236 n0_17304_4375 n2_17304_4375 0.0
V23237 n0_17304_4521 n2_17304_4521 0.0
V23238 n0_17304_4554 n2_17304_4554 0.0
V23239 n0_17304_4591 n2_17304_4591 0.0
V23240 n0_17304_4737 n2_17304_4737 0.0
V23241 n0_17304_4770 n2_17304_4770 0.0
V23242 n0_17304_4807 n2_17304_4807 0.0
V23243 n0_17304_5169 n2_17304_5169 0.0
V23244 n0_17304_5202 n2_17304_5202 0.0
V23245 n0_17304_5239 n2_17304_5239 0.0
V23246 n0_17304_5385 n2_17304_5385 0.0
V23247 n0_17304_5418 n2_17304_5418 0.0
V23248 n0_17304_5455 n2_17304_5455 0.0
V23249 n0_17304_5601 n2_17304_5601 0.0
V23250 n0_17304_5634 n2_17304_5634 0.0
V23251 n0_17304_5817 n2_17304_5817 0.0
V23252 n0_17304_5850 n2_17304_5850 0.0
V23253 n0_17304_6033 n2_17304_6033 0.0
V23254 n0_17304_6066 n2_17304_6066 0.0
V23255 n0_17304_6249 n2_17304_6249 0.0
V23256 n0_17304_6282 n2_17304_6282 0.0
V23257 n0_17304_6319 n2_17304_6319 0.0
V23258 n0_17304_6465 n2_17304_6465 0.0
V23259 n0_17304_6498 n2_17304_6498 0.0
V23260 n0_17304_6681 n2_17304_6681 0.0
V23261 n0_17304_6714 n2_17304_6714 0.0
V23262 n0_17304_6897 n2_17304_6897 0.0
V23263 n0_17304_6930 n2_17304_6930 0.0
V23264 n0_17304_7113 n2_17304_7113 0.0
V23265 n0_17304_7329 n2_17304_7329 0.0
V23266 n0_17304_7362 n2_17304_7362 0.0
V23267 n0_17304_7545 n2_17304_7545 0.0
V23268 n0_17304_7578 n2_17304_7578 0.0
V23269 n0_17304_7761 n2_17304_7761 0.0
V23270 n0_17304_7794 n2_17304_7794 0.0
V23271 n0_17304_7831 n2_17304_7831 0.0
V23272 n0_17304_7977 n2_17304_7977 0.0
V23273 n0_17304_8010 n2_17304_8010 0.0
V23274 n0_17304_8193 n2_17304_8193 0.0
V23275 n0_17304_8226 n2_17304_8226 0.0
V23276 n0_17304_8409 n2_17304_8409 0.0
V23277 n0_17304_8442 n2_17304_8442 0.0
V23278 n0_17304_8625 n2_17304_8625 0.0
V23279 n0_17304_8658 n2_17304_8658 0.0
V23280 n0_17304_8841 n2_17304_8841 0.0
V23281 n0_17304_8874 n2_17304_8874 0.0
V23282 n0_17304_8911 n2_17304_8911 0.0
V23283 n0_17304_9057 n2_17304_9057 0.0
V23284 n0_17304_9090 n2_17304_9090 0.0
V23285 n0_17304_9273 n2_17304_9273 0.0
V23286 n0_17304_9306 n2_17304_9306 0.0
V23287 n0_17304_9705 n2_17304_9705 0.0
V23288 n0_17304_9738 n2_17304_9738 0.0
V23289 n0_17304_9921 n2_17304_9921 0.0
V23290 n0_17304_9954 n2_17304_9954 0.0
V23291 n0_17304_9991 n2_17304_9991 0.0
V23292 n0_17304_10137 n2_17304_10137 0.0
V23293 n0_17304_10170 n2_17304_10170 0.0
V23294 n0_17304_10353 n2_17304_10353 0.0
V23295 n0_17304_10386 n2_17304_10386 0.0
V23296 n0_17304_10569 n2_17304_10569 0.0
V23297 n0_17304_10602 n2_17304_10602 0.0
V23298 n0_17304_10785 n2_17304_10785 0.0
V23299 n0_17304_10818 n2_17304_10818 0.0
V23300 n0_17304_11001 n2_17304_11001 0.0
V23301 n0_17304_11034 n2_17304_11034 0.0
V23302 n0_17304_11048 n2_17304_11048 0.0
V23303 n0_17304_11055 n2_17304_11055 0.0
V23304 n0_17304_11217 n2_17304_11217 0.0
V23305 n0_17304_11250 n2_17304_11250 0.0
V23306 n0_17304_11433 n2_17304_11433 0.0
V23307 n0_17304_11466 n2_17304_11466 0.0
V23308 n0_17304_11865 n2_17304_11865 0.0
V23309 n0_17304_11898 n2_17304_11898 0.0
V23310 n0_17304_12081 n2_17304_12081 0.0
V23311 n0_17304_12114 n2_17304_12114 0.0
V23312 n0_17304_12128 n2_17304_12128 0.0
V23313 n0_17304_12135 n2_17304_12135 0.0
V23314 n0_17304_12297 n2_17304_12297 0.0
V23315 n0_17304_12330 n2_17304_12330 0.0
V23316 n0_17304_12513 n2_17304_12513 0.0
V23317 n0_17304_12546 n2_17304_12546 0.0
V23318 n0_17304_12729 n2_17304_12729 0.0
V23319 n0_17304_12762 n2_17304_12762 0.0
V23320 n0_17304_12945 n2_17304_12945 0.0
V23321 n0_17304_12978 n2_17304_12978 0.0
V23322 n0_17304_13161 n2_17304_13161 0.0
V23323 n0_17304_13194 n2_17304_13194 0.0
V23324 n0_17304_13377 n2_17304_13377 0.0
V23325 n0_17304_13410 n2_17304_13410 0.0
V23326 n0_17304_13423 n2_17304_13423 0.0
V23327 n0_17304_13593 n2_17304_13593 0.0
V23328 n0_17304_13626 n2_17304_13626 0.0
V23329 n0_17304_13640 n2_17304_13640 0.0
V23330 n0_17304_13647 n2_17304_13647 0.0
V23331 n0_17304_13809 n2_17304_13809 0.0
V23332 n0_17304_13842 n2_17304_13842 0.0
V23333 n0_17304_14241 n2_17304_14241 0.0
V23334 n0_17304_14274 n2_17304_14274 0.0
V23335 n0_17304_14457 n2_17304_14457 0.0
V23336 n0_17304_14490 n2_17304_14490 0.0
V23337 n0_17304_14511 n2_17304_14511 0.0
V23338 n0_17304_14673 n2_17304_14673 0.0
V23339 n0_17304_14706 n2_17304_14706 0.0
V23340 n0_17304_14889 n2_17304_14889 0.0
V23341 n0_17304_14922 n2_17304_14922 0.0
V23342 n0_17304_14936 n2_17304_14936 0.0
V23343 n0_17304_14943 n2_17304_14943 0.0
V23344 n0_17304_15105 n2_17304_15105 0.0
V23345 n0_17304_15138 n2_17304_15138 0.0
V23346 n0_17304_15152 n2_17304_15152 0.0
V23347 n0_17304_15159 n2_17304_15159 0.0
V23348 n0_17304_15321 n2_17304_15321 0.0
V23349 n0_17304_15354 n2_17304_15354 0.0
V23350 n0_17304_15537 n2_17304_15537 0.0
V23351 n0_17304_15570 n2_17304_15570 0.0
V23352 n0_17304_15584 n2_17304_15584 0.0
V23353 n0_17304_15753 n2_17304_15753 0.0
V23354 n0_17304_15786 n2_17304_15786 0.0
V23355 n0_17304_15969 n2_17304_15969 0.0
V23356 n0_17304_16002 n2_17304_16002 0.0
V23357 n0_17304_16401 n2_17304_16401 0.0
V23358 n0_17304_16434 n2_17304_16434 0.0
V23359 n0_17304_16617 n2_17304_16617 0.0
V23360 n0_17304_16650 n2_17304_16650 0.0
V23361 n0_17304_16664 n2_17304_16664 0.0
V23362 n0_17304_16687 n2_17304_16687 0.0
V23363 n0_17304_16833 n2_17304_16833 0.0
V23364 n0_17304_16866 n2_17304_16866 0.0
V23365 n0_17304_17049 n2_17304_17049 0.0
V23366 n0_17304_17082 n2_17304_17082 0.0
V23367 n0_17304_17119 n2_17304_17119 0.0
V23368 n0_17304_17265 n2_17304_17265 0.0
V23369 n0_17304_17298 n2_17304_17298 0.0
V23370 n0_17304_17481 n2_17304_17481 0.0
V23371 n0_17304_17514 n2_17304_17514 0.0
V23372 n0_17304_17535 n2_17304_17535 0.0
V23373 n0_17304_17697 n2_17304_17697 0.0
V23374 n0_17304_17730 n2_17304_17730 0.0
V23375 n0_17304_17913 n2_17304_17913 0.0
V23376 n0_17304_17946 n2_17304_17946 0.0
V23377 n0_17304_18129 n2_17304_18129 0.0
V23378 n0_17304_18162 n2_17304_18162 0.0
V23379 n0_17304_18176 n2_17304_18176 0.0
V23380 n0_17304_18345 n2_17304_18345 0.0
V23381 n0_17304_18378 n2_17304_18378 0.0
V23382 n0_17304_18561 n2_17304_18561 0.0
V23383 n0_17304_18594 n2_17304_18594 0.0
V23384 n0_17304_18777 n2_17304_18777 0.0
V23385 n0_17304_18810 n2_17304_18810 0.0
V23386 n0_17304_18993 n2_17304_18993 0.0
V23387 n0_17304_19026 n2_17304_19026 0.0
V23388 n0_17304_19040 n2_17304_19040 0.0
V23389 n0_17304_19209 n2_17304_19209 0.0
V23390 n0_17304_19242 n2_17304_19242 0.0
V23391 n0_17304_19425 n2_17304_19425 0.0
V23392 n0_17304_19458 n2_17304_19458 0.0
V23393 n0_17304_19641 n2_17304_19641 0.0
V23394 n0_17304_19674 n2_17304_19674 0.0
V23395 n0_17304_19857 n2_17304_19857 0.0
V23396 n0_17304_19890 n2_17304_19890 0.0
V23397 n0_17304_20073 n2_17304_20073 0.0
V23398 n0_17304_20106 n2_17304_20106 0.0
V23399 n0_17304_20289 n2_17304_20289 0.0
V23400 n0_17304_20322 n2_17304_20322 0.0
V23401 n0_17304_20505 n2_17304_20505 0.0
V23402 n0_17304_20538 n2_17304_20538 0.0
V23403 n0_17304_20721 n2_17304_20721 0.0
V23404 n0_17304_20754 n2_17304_20754 0.0
V23405 n0_17304_20937 n2_17304_20937 0.0
V23406 n0_17304_20970 n2_17304_20970 0.0
V23407 n0_17396_201 n2_17396_201 0.0
V23408 n0_17396_234 n2_17396_234 0.0
V23409 n0_17396_417 n2_17396_417 0.0
V23410 n0_17396_450 n2_17396_450 0.0
V23411 n0_17396_633 n2_17396_633 0.0
V23412 n0_17396_666 n2_17396_666 0.0
V23413 n0_17396_849 n2_17396_849 0.0
V23414 n0_17396_882 n2_17396_882 0.0
V23415 n0_17396_1065 n2_17396_1065 0.0
V23416 n0_17396_1098 n2_17396_1098 0.0
V23417 n0_17396_1281 n2_17396_1281 0.0
V23418 n0_17396_1314 n2_17396_1314 0.0
V23419 n0_17396_1497 n2_17396_1497 0.0
V23420 n0_17396_1530 n2_17396_1530 0.0
V23421 n0_17396_1713 n2_17396_1713 0.0
V23422 n0_17396_1746 n2_17396_1746 0.0
V23423 n0_17396_1783 n2_17396_1783 0.0
V23424 n0_17396_1929 n2_17396_1929 0.0
V23425 n0_17396_1962 n2_17396_1962 0.0
V23426 n0_17396_2145 n2_17396_2145 0.0
V23427 n0_17396_2178 n2_17396_2178 0.0
V23428 n0_17396_2361 n2_17396_2361 0.0
V23429 n0_17396_2394 n2_17396_2394 0.0
V23430 n0_17396_2431 n2_17396_2431 0.0
V23431 n0_17396_2577 n2_17396_2577 0.0
V23432 n0_17396_2610 n2_17396_2610 0.0
V23433 n0_17396_2793 n2_17396_2793 0.0
V23434 n0_17396_2826 n2_17396_2826 0.0
V23435 n0_17396_2863 n2_17396_2863 0.0
V23436 n0_17396_3009 n2_17396_3009 0.0
V23437 n0_17396_3042 n2_17396_3042 0.0
V23438 n0_17396_3225 n2_17396_3225 0.0
V23439 n0_17396_3258 n2_17396_3258 0.0
V23440 n0_17396_3295 n2_17396_3295 0.0
V23441 n0_17396_3441 n2_17396_3441 0.0
V23442 n0_17396_3474 n2_17396_3474 0.0
V23443 n0_17396_3657 n2_17396_3657 0.0
V23444 n0_17396_3690 n2_17396_3690 0.0
V23445 n0_17396_17481 n2_17396_17481 0.0
V23446 n0_17396_17514 n2_17396_17514 0.0
V23447 n0_17396_17535 n2_17396_17535 0.0
V23448 n0_17396_17697 n2_17396_17697 0.0
V23449 n0_17396_17730 n2_17396_17730 0.0
V23450 n0_17396_17913 n2_17396_17913 0.0
V23451 n0_17396_17946 n2_17396_17946 0.0
V23452 n0_17396_18129 n2_17396_18129 0.0
V23453 n0_17396_18162 n2_17396_18162 0.0
V23454 n0_17396_18176 n2_17396_18176 0.0
V23455 n0_17396_18345 n2_17396_18345 0.0
V23456 n0_17396_18378 n2_17396_18378 0.0
V23457 n0_17396_18561 n2_17396_18561 0.0
V23458 n0_17396_18594 n2_17396_18594 0.0
V23459 n0_17396_18777 n2_17396_18777 0.0
V23460 n0_17396_18810 n2_17396_18810 0.0
V23461 n0_17396_18993 n2_17396_18993 0.0
V23462 n0_17396_19026 n2_17396_19026 0.0
V23463 n0_17396_19040 n2_17396_19040 0.0
V23464 n0_17396_19209 n2_17396_19209 0.0
V23465 n0_17396_19242 n2_17396_19242 0.0
V23466 n0_17396_19425 n2_17396_19425 0.0
V23467 n0_17396_19458 n2_17396_19458 0.0
V23468 n0_17396_19641 n2_17396_19641 0.0
V23469 n0_17396_19674 n2_17396_19674 0.0
V23470 n0_17396_19857 n2_17396_19857 0.0
V23471 n0_17396_19890 n2_17396_19890 0.0
V23472 n0_17396_20073 n2_17396_20073 0.0
V23473 n0_17396_20106 n2_17396_20106 0.0
V23474 n0_17396_20289 n2_17396_20289 0.0
V23475 n0_17396_20322 n2_17396_20322 0.0
V23476 n0_17396_20505 n2_17396_20505 0.0
V23477 n0_17396_20538 n2_17396_20538 0.0
V23478 n0_17396_20754 n2_17396_20754 0.0
V23479 n0_17396_20937 n2_17396_20937 0.0
V23480 n0_17396_20970 n2_17396_20970 0.0
V23481 n0_18241_2793 n2_18241_2793 0.0
V23482 n0_18241_2826 n2_18241_2826 0.0
V23483 n0_18241_3009 n2_18241_3009 0.0
V23484 n0_18241_3042 n2_18241_3042 0.0
V23485 n0_18241_3225 n2_18241_3225 0.0
V23486 n0_18241_3258 n2_18241_3258 0.0
V23487 n0_18241_3295 n2_18241_3295 0.0
V23488 n0_18241_3441 n2_18241_3441 0.0
V23489 n0_18241_3474 n2_18241_3474 0.0
V23490 n0_18241_3657 n2_18241_3657 0.0
V23491 n0_18241_3690 n2_18241_3690 0.0
V23492 n0_18241_3873 n2_18241_3873 0.0
V23493 n0_18241_3906 n2_18241_3906 0.0
V23494 n0_18241_4089 n2_18241_4089 0.0
V23495 n0_18241_4122 n2_18241_4122 0.0
V23496 n0_18241_4305 n2_18241_4305 0.0
V23497 n0_18241_4338 n2_18241_4338 0.0
V23498 n0_18241_4375 n2_18241_4375 0.0
V23499 n0_18241_4521 n2_18241_4521 0.0
V23500 n0_18241_4554 n2_18241_4554 0.0
V23501 n0_18241_4591 n2_18241_4591 0.0
V23502 n0_18241_4737 n2_18241_4737 0.0
V23503 n0_18241_4770 n2_18241_4770 0.0
V23504 n0_18241_4807 n2_18241_4807 0.0
V23505 n0_18241_4953 n2_18241_4953 0.0
V23506 n0_18241_4986 n2_18241_4986 0.0
V23507 n0_18241_5023 n2_18241_5023 0.0
V23508 n0_18241_5169 n2_18241_5169 0.0
V23509 n0_18241_5202 n2_18241_5202 0.0
V23510 n0_18241_5239 n2_18241_5239 0.0
V23511 n0_18241_5385 n2_18241_5385 0.0
V23512 n0_18241_5418 n2_18241_5418 0.0
V23513 n0_18241_5455 n2_18241_5455 0.0
V23514 n0_18241_5601 n2_18241_5601 0.0
V23515 n0_18241_5634 n2_18241_5634 0.0
V23516 n0_18241_5817 n2_18241_5817 0.0
V23517 n0_18241_5850 n2_18241_5850 0.0
V23518 n0_18241_6033 n2_18241_6033 0.0
V23519 n0_18241_6066 n2_18241_6066 0.0
V23520 n0_18241_6249 n2_18241_6249 0.0
V23521 n0_18241_6282 n2_18241_6282 0.0
V23522 n0_18241_6319 n2_18241_6319 0.0
V23523 n0_18241_6465 n2_18241_6465 0.0
V23524 n0_18241_6498 n2_18241_6498 0.0
V23525 n0_18241_6681 n2_18241_6681 0.0
V23526 n0_18241_6714 n2_18241_6714 0.0
V23527 n0_18241_6897 n2_18241_6897 0.0
V23528 n0_18241_6930 n2_18241_6930 0.0
V23529 n0_18241_7113 n2_18241_7113 0.0
V23530 n0_18241_7146 n2_18241_7146 0.0
V23531 n0_18241_7329 n2_18241_7329 0.0
V23532 n0_18241_7362 n2_18241_7362 0.0
V23533 n0_18241_7545 n2_18241_7545 0.0
V23534 n0_18241_7578 n2_18241_7578 0.0
V23535 n0_18241_7761 n2_18241_7761 0.0
V23536 n0_18241_7794 n2_18241_7794 0.0
V23537 n0_18241_7831 n2_18241_7831 0.0
V23538 n0_18241_7977 n2_18241_7977 0.0
V23539 n0_18241_8010 n2_18241_8010 0.0
V23540 n0_18241_8193 n2_18241_8193 0.0
V23541 n0_18241_8226 n2_18241_8226 0.0
V23542 n0_18241_8409 n2_18241_8409 0.0
V23543 n0_18241_8442 n2_18241_8442 0.0
V23544 n0_18241_8625 n2_18241_8625 0.0
V23545 n0_18241_8658 n2_18241_8658 0.0
V23546 n0_18241_8841 n2_18241_8841 0.0
V23547 n0_18241_8874 n2_18241_8874 0.0
V23548 n0_18241_8911 n2_18241_8911 0.0
V23549 n0_18241_9057 n2_18241_9057 0.0
V23550 n0_18241_9090 n2_18241_9090 0.0
V23551 n0_18241_9273 n2_18241_9273 0.0
V23552 n0_18241_9306 n2_18241_9306 0.0
V23553 n0_18241_9489 n2_18241_9489 0.0
V23554 n0_18241_9522 n2_18241_9522 0.0
V23555 n0_18241_9705 n2_18241_9705 0.0
V23556 n0_18241_9738 n2_18241_9738 0.0
V23557 n0_18241_9921 n2_18241_9921 0.0
V23558 n0_18241_9954 n2_18241_9954 0.0
V23559 n0_18241_9991 n2_18241_9991 0.0
V23560 n0_18241_10137 n2_18241_10137 0.0
V23561 n0_18241_10170 n2_18241_10170 0.0
V23562 n0_18241_10353 n2_18241_10353 0.0
V23563 n0_18241_10386 n2_18241_10386 0.0
V23564 n0_18241_10569 n2_18241_10569 0.0
V23565 n0_18241_10785 n2_18241_10785 0.0
V23566 n0_18241_10818 n2_18241_10818 0.0
V23567 n0_18241_11001 n2_18241_11001 0.0
V23568 n0_18241_11034 n2_18241_11034 0.0
V23569 n0_18241_11055 n2_18241_11055 0.0
V23570 n0_18241_11217 n2_18241_11217 0.0
V23571 n0_18241_11250 n2_18241_11250 0.0
V23572 n0_18241_11433 n2_18241_11433 0.0
V23573 n0_18241_11466 n2_18241_11466 0.0
V23574 n0_18241_11649 n2_18241_11649 0.0
V23575 n0_18241_11682 n2_18241_11682 0.0
V23576 n0_18241_11865 n2_18241_11865 0.0
V23577 n0_18241_11898 n2_18241_11898 0.0
V23578 n0_18241_12081 n2_18241_12081 0.0
V23579 n0_18241_12114 n2_18241_12114 0.0
V23580 n0_18241_12128 n2_18241_12128 0.0
V23581 n0_18241_12297 n2_18241_12297 0.0
V23582 n0_18241_12330 n2_18241_12330 0.0
V23583 n0_18241_12513 n2_18241_12513 0.0
V23584 n0_18241_12546 n2_18241_12546 0.0
V23585 n0_18241_12729 n2_18241_12729 0.0
V23586 n0_18241_12762 n2_18241_12762 0.0
V23587 n0_18241_12945 n2_18241_12945 0.0
V23588 n0_18241_12978 n2_18241_12978 0.0
V23589 n0_18241_13161 n2_18241_13161 0.0
V23590 n0_18241_13194 n2_18241_13194 0.0
V23591 n0_18241_13377 n2_18241_13377 0.0
V23592 n0_18241_13410 n2_18241_13410 0.0
V23593 n0_18241_13593 n2_18241_13593 0.0
V23594 n0_18241_13626 n2_18241_13626 0.0
V23595 n0_18241_13640 n2_18241_13640 0.0
V23596 n0_18241_13647 n2_18241_13647 0.0
V23597 n0_18241_13809 n2_18241_13809 0.0
V23598 n0_18241_13842 n2_18241_13842 0.0
V23599 n0_18241_14025 n2_18241_14025 0.0
V23600 n0_18241_14058 n2_18241_14058 0.0
V23601 n0_18241_14241 n2_18241_14241 0.0
V23602 n0_18241_14274 n2_18241_14274 0.0
V23603 n0_18241_14457 n2_18241_14457 0.0
V23604 n0_18241_14490 n2_18241_14490 0.0
V23605 n0_18241_14504 n2_18241_14504 0.0
V23606 n0_18241_14511 n2_18241_14511 0.0
V23607 n0_18241_14673 n2_18241_14673 0.0
V23608 n0_18241_14706 n2_18241_14706 0.0
V23609 n0_18241_14889 n2_18241_14889 0.0
V23610 n0_18241_14922 n2_18241_14922 0.0
V23611 n0_18241_14936 n2_18241_14936 0.0
V23612 n0_18241_15138 n2_18241_15138 0.0
V23613 n0_18241_15152 n2_18241_15152 0.0
V23614 n0_18241_15321 n2_18241_15321 0.0
V23615 n0_18241_15354 n2_18241_15354 0.0
V23616 n0_18241_15537 n2_18241_15537 0.0
V23617 n0_18241_15570 n2_18241_15570 0.0
V23618 n0_18241_15584 n2_18241_15584 0.0
V23619 n0_18241_15753 n2_18241_15753 0.0
V23620 n0_18241_15786 n2_18241_15786 0.0
V23621 n0_18241_15969 n2_18241_15969 0.0
V23622 n0_18241_16002 n2_18241_16002 0.0
V23623 n0_18241_16185 n2_18241_16185 0.0
V23624 n0_18241_16218 n2_18241_16218 0.0
V23625 n0_18241_16401 n2_18241_16401 0.0
V23626 n0_18241_16434 n2_18241_16434 0.0
V23627 n0_18241_16617 n2_18241_16617 0.0
V23628 n0_18241_16650 n2_18241_16650 0.0
V23629 n0_18241_16664 n2_18241_16664 0.0
V23630 n0_18241_16671 n2_18241_16671 0.0
V23631 n0_18241_16833 n2_18241_16833 0.0
V23632 n0_18241_16866 n2_18241_16866 0.0
V23633 n0_18241_17049 n2_18241_17049 0.0
V23634 n0_18241_17082 n2_18241_17082 0.0
V23635 n0_18241_17119 n2_18241_17119 0.0
V23636 n0_18241_17265 n2_18241_17265 0.0
V23637 n0_18241_17298 n2_18241_17298 0.0
V23638 n0_18241_17481 n2_18241_17481 0.0
V23639 n0_18241_17514 n2_18241_17514 0.0
V23640 n0_18241_17697 n2_18241_17697 0.0
V23641 n0_18241_17730 n2_18241_17730 0.0
V23642 n0_18241_17744 n2_18241_17744 0.0
V23643 n0_18241_17913 n2_18241_17913 0.0
V23644 n0_18241_17946 n2_18241_17946 0.0
V23645 n0_18241_18129 n2_18241_18129 0.0
V23646 n0_18241_18162 n2_18241_18162 0.0
V23647 n0_18241_18345 n2_18241_18345 0.0
V23648 n0_18241_18378 n2_18241_18378 0.0
V23649 n0_18380_3873 n2_18380_3873 0.0
V23650 n0_18380_3906 n2_18380_3906 0.0
V23651 n0_18380_6033 n2_18380_6033 0.0
V23652 n0_18380_6066 n2_18380_6066 0.0
V23653 n0_18380_8409 n2_18380_8409 0.0
V23654 n0_18380_10569 n2_18380_10569 0.0
V23655 n0_18380_10602 n2_18380_10602 0.0
V23656 n0_18380_15105 n2_18380_15105 0.0
V23657 n0_18380_15138 n2_18380_15138 0.0
V23658 n0_18380_15152 n2_18380_15152 0.0
V23659 n0_18380_17298 n2_18380_17298 0.0
V23660 n0_18429_2826 n2_18429_2826 0.0
V23661 n0_18429_3009 n2_18429_3009 0.0
V23662 n0_18429_3042 n2_18429_3042 0.0
V23663 n0_18429_3225 n2_18429_3225 0.0
V23664 n0_18429_3258 n2_18429_3258 0.0
V23665 n0_18429_3295 n2_18429_3295 0.0
V23666 n0_18429_3441 n2_18429_3441 0.0
V23667 n0_18429_3474 n2_18429_3474 0.0
V23668 n0_18429_3657 n2_18429_3657 0.0
V23669 n0_18429_3690 n2_18429_3690 0.0
V23670 n0_18429_3873 n2_18429_3873 0.0
V23671 n0_18429_3906 n2_18429_3906 0.0
V23672 n0_18429_4089 n2_18429_4089 0.0
V23673 n0_18429_4122 n2_18429_4122 0.0
V23674 n0_18429_4305 n2_18429_4305 0.0
V23675 n0_18429_4338 n2_18429_4338 0.0
V23676 n0_18429_4375 n2_18429_4375 0.0
V23677 n0_18429_4521 n2_18429_4521 0.0
V23678 n0_18429_4554 n2_18429_4554 0.0
V23679 n0_18429_4591 n2_18429_4591 0.0
V23680 n0_18429_4737 n2_18429_4737 0.0
V23681 n0_18429_4770 n2_18429_4770 0.0
V23682 n0_18429_4807 n2_18429_4807 0.0
V23683 n0_18429_5169 n2_18429_5169 0.0
V23684 n0_18429_5202 n2_18429_5202 0.0
V23685 n0_18429_5239 n2_18429_5239 0.0
V23686 n0_18429_5385 n2_18429_5385 0.0
V23687 n0_18429_5418 n2_18429_5418 0.0
V23688 n0_18429_5455 n2_18429_5455 0.0
V23689 n0_18429_5601 n2_18429_5601 0.0
V23690 n0_18429_5634 n2_18429_5634 0.0
V23691 n0_18429_5817 n2_18429_5817 0.0
V23692 n0_18429_5850 n2_18429_5850 0.0
V23693 n0_18429_6033 n2_18429_6033 0.0
V23694 n0_18429_6066 n2_18429_6066 0.0
V23695 n0_18429_6249 n2_18429_6249 0.0
V23696 n0_18429_6282 n2_18429_6282 0.0
V23697 n0_18429_6319 n2_18429_6319 0.0
V23698 n0_18429_6465 n2_18429_6465 0.0
V23699 n0_18429_6498 n2_18429_6498 0.0
V23700 n0_18429_6681 n2_18429_6681 0.0
V23701 n0_18429_6714 n2_18429_6714 0.0
V23702 n0_18429_6897 n2_18429_6897 0.0
V23703 n0_18429_6930 n2_18429_6930 0.0
V23704 n0_18429_7113 n2_18429_7113 0.0
V23705 n0_18429_7329 n2_18429_7329 0.0
V23706 n0_18429_7362 n2_18429_7362 0.0
V23707 n0_18429_7545 n2_18429_7545 0.0
V23708 n0_18429_7578 n2_18429_7578 0.0
V23709 n0_18429_7761 n2_18429_7761 0.0
V23710 n0_18429_7794 n2_18429_7794 0.0
V23711 n0_18429_7831 n2_18429_7831 0.0
V23712 n0_18429_7977 n2_18429_7977 0.0
V23713 n0_18429_8010 n2_18429_8010 0.0
V23714 n0_18429_8193 n2_18429_8193 0.0
V23715 n0_18429_8226 n2_18429_8226 0.0
V23716 n0_18429_8409 n2_18429_8409 0.0
V23717 n0_18429_8442 n2_18429_8442 0.0
V23718 n0_18429_8625 n2_18429_8625 0.0
V23719 n0_18429_8658 n2_18429_8658 0.0
V23720 n0_18429_8841 n2_18429_8841 0.0
V23721 n0_18429_8874 n2_18429_8874 0.0
V23722 n0_18429_8911 n2_18429_8911 0.0
V23723 n0_18429_9057 n2_18429_9057 0.0
V23724 n0_18429_9090 n2_18429_9090 0.0
V23725 n0_18429_9273 n2_18429_9273 0.0
V23726 n0_18429_9306 n2_18429_9306 0.0
V23727 n0_18429_9705 n2_18429_9705 0.0
V23728 n0_18429_9738 n2_18429_9738 0.0
V23729 n0_18429_9921 n2_18429_9921 0.0
V23730 n0_18429_9954 n2_18429_9954 0.0
V23731 n0_18429_9991 n2_18429_9991 0.0
V23732 n0_18429_10137 n2_18429_10137 0.0
V23733 n0_18429_10170 n2_18429_10170 0.0
V23734 n0_18429_10353 n2_18429_10353 0.0
V23735 n0_18429_10386 n2_18429_10386 0.0
V23736 n0_18429_10569 n2_18429_10569 0.0
V23737 n0_18429_10602 n2_18429_10602 0.0
V23738 n0_18429_10785 n2_18429_10785 0.0
V23739 n0_18429_10818 n2_18429_10818 0.0
V23740 n0_18429_11001 n2_18429_11001 0.0
V23741 n0_18429_11034 n2_18429_11034 0.0
V23742 n0_18429_11055 n2_18429_11055 0.0
V23743 n0_18429_11217 n2_18429_11217 0.0
V23744 n0_18429_11250 n2_18429_11250 0.0
V23745 n0_18429_11433 n2_18429_11433 0.0
V23746 n0_18429_11466 n2_18429_11466 0.0
V23747 n0_18429_11865 n2_18429_11865 0.0
V23748 n0_18429_11898 n2_18429_11898 0.0
V23749 n0_18429_12081 n2_18429_12081 0.0
V23750 n0_18429_12114 n2_18429_12114 0.0
V23751 n0_18429_12128 n2_18429_12128 0.0
V23752 n0_18429_12297 n2_18429_12297 0.0
V23753 n0_18429_12330 n2_18429_12330 0.0
V23754 n0_18429_12513 n2_18429_12513 0.0
V23755 n0_18429_12546 n2_18429_12546 0.0
V23756 n0_18429_12729 n2_18429_12729 0.0
V23757 n0_18429_12762 n2_18429_12762 0.0
V23758 n0_18429_12945 n2_18429_12945 0.0
V23759 n0_18429_12978 n2_18429_12978 0.0
V23760 n0_18429_13161 n2_18429_13161 0.0
V23761 n0_18429_13194 n2_18429_13194 0.0
V23762 n0_18429_13377 n2_18429_13377 0.0
V23763 n0_18429_13410 n2_18429_13410 0.0
V23764 n0_18429_13423 n2_18429_13423 0.0
V23765 n0_18429_13593 n2_18429_13593 0.0
V23766 n0_18429_13626 n2_18429_13626 0.0
V23767 n0_18429_13640 n2_18429_13640 0.0
V23768 n0_18429_13647 n2_18429_13647 0.0
V23769 n0_18429_13809 n2_18429_13809 0.0
V23770 n0_18429_13842 n2_18429_13842 0.0
V23771 n0_18429_14241 n2_18429_14241 0.0
V23772 n0_18429_14274 n2_18429_14274 0.0
V23773 n0_18429_14457 n2_18429_14457 0.0
V23774 n0_18429_14490 n2_18429_14490 0.0
V23775 n0_18429_14504 n2_18429_14504 0.0
V23776 n0_18429_14511 n2_18429_14511 0.0
V23777 n0_18429_14673 n2_18429_14673 0.0
V23778 n0_18429_14706 n2_18429_14706 0.0
V23779 n0_18429_14889 n2_18429_14889 0.0
V23780 n0_18429_14922 n2_18429_14922 0.0
V23781 n0_18429_14936 n2_18429_14936 0.0
V23782 n0_18429_15105 n2_18429_15105 0.0
V23783 n0_18429_15138 n2_18429_15138 0.0
V23784 n0_18429_15152 n2_18429_15152 0.0
V23785 n0_18429_15321 n2_18429_15321 0.0
V23786 n0_18429_15354 n2_18429_15354 0.0
V23787 n0_18429_15537 n2_18429_15537 0.0
V23788 n0_18429_15570 n2_18429_15570 0.0
V23789 n0_18429_15584 n2_18429_15584 0.0
V23790 n0_18429_15753 n2_18429_15753 0.0
V23791 n0_18429_15786 n2_18429_15786 0.0
V23792 n0_18429_15969 n2_18429_15969 0.0
V23793 n0_18429_16002 n2_18429_16002 0.0
V23794 n0_18429_16401 n2_18429_16401 0.0
V23795 n0_18429_16434 n2_18429_16434 0.0
V23796 n0_18429_16617 n2_18429_16617 0.0
V23797 n0_18429_16650 n2_18429_16650 0.0
V23798 n0_18429_16664 n2_18429_16664 0.0
V23799 n0_18429_16671 n2_18429_16671 0.0
V23800 n0_18429_16833 n2_18429_16833 0.0
V23801 n0_18429_16866 n2_18429_16866 0.0
V23802 n0_18429_17049 n2_18429_17049 0.0
V23803 n0_18429_17082 n2_18429_17082 0.0
V23804 n0_18429_17119 n2_18429_17119 0.0
V23805 n0_18429_17265 n2_18429_17265 0.0
V23806 n0_18429_17298 n2_18429_17298 0.0
V23807 n0_18429_17481 n2_18429_17481 0.0
V23808 n0_18429_17514 n2_18429_17514 0.0
V23809 n0_18429_17697 n2_18429_17697 0.0
V23810 n0_18429_17730 n2_18429_17730 0.0
V23811 n0_18429_17744 n2_18429_17744 0.0
V23812 n0_18429_17913 n2_18429_17913 0.0
V23813 n0_18429_17946 n2_18429_17946 0.0
V23814 n0_18429_18129 n2_18429_18129 0.0
V23815 n0_18429_18162 n2_18429_18162 0.0
V23816 n0_18429_18345 n2_18429_18345 0.0
V23817 n0_19366_201 n2_19366_201 0.0
V23818 n0_19366_234 n2_19366_234 0.0
V23819 n0_19366_417 n2_19366_417 0.0
V23820 n0_19366_450 n2_19366_450 0.0
V23821 n0_19366_633 n2_19366_633 0.0
V23822 n0_19366_666 n2_19366_666 0.0
V23823 n0_19366_849 n2_19366_849 0.0
V23824 n0_19366_882 n2_19366_882 0.0
V23825 n0_19366_1065 n2_19366_1065 0.0
V23826 n0_19366_1098 n2_19366_1098 0.0
V23827 n0_19366_1281 n2_19366_1281 0.0
V23828 n0_19366_1314 n2_19366_1314 0.0
V23829 n0_19366_1497 n2_19366_1497 0.0
V23830 n0_19366_1530 n2_19366_1530 0.0
V23831 n0_19366_1713 n2_19366_1713 0.0
V23832 n0_19366_1746 n2_19366_1746 0.0
V23833 n0_19366_1929 n2_19366_1929 0.0
V23834 n0_19366_1962 n2_19366_1962 0.0
V23835 n0_19366_1976 n2_19366_1976 0.0
V23836 n0_19366_1999 n2_19366_1999 0.0
V23837 n0_19366_2145 n2_19366_2145 0.0
V23838 n0_19366_2178 n2_19366_2178 0.0
V23839 n0_19366_2361 n2_19366_2361 0.0
V23840 n0_19366_2394 n2_19366_2394 0.0
V23841 n0_19366_2577 n2_19366_2577 0.0
V23842 n0_19366_2610 n2_19366_2610 0.0
V23843 n0_19366_2793 n2_19366_2793 0.0
V23844 n0_19366_2826 n2_19366_2826 0.0
V23845 n0_19366_3009 n2_19366_3009 0.0
V23846 n0_19366_3042 n2_19366_3042 0.0
V23847 n0_19366_3225 n2_19366_3225 0.0
V23848 n0_19366_3258 n2_19366_3258 0.0
V23849 n0_19366_3295 n2_19366_3295 0.0
V23850 n0_19366_3441 n2_19366_3441 0.0
V23851 n0_19366_3474 n2_19366_3474 0.0
V23852 n0_19366_3657 n2_19366_3657 0.0
V23853 n0_19366_3690 n2_19366_3690 0.0
V23854 n0_19366_3873 n2_19366_3873 0.0
V23855 n0_19366_3906 n2_19366_3906 0.0
V23856 n0_19366_4089 n2_19366_4089 0.0
V23857 n0_19366_4122 n2_19366_4122 0.0
V23858 n0_19366_4305 n2_19366_4305 0.0
V23859 n0_19366_4338 n2_19366_4338 0.0
V23860 n0_19366_4375 n2_19366_4375 0.0
V23861 n0_19366_4521 n2_19366_4521 0.0
V23862 n0_19366_4554 n2_19366_4554 0.0
V23863 n0_19366_4737 n2_19366_4737 0.0
V23864 n0_19366_4770 n2_19366_4770 0.0
V23865 n0_19366_4953 n2_19366_4953 0.0
V23866 n0_19366_4986 n2_19366_4986 0.0
V23867 n0_19366_5169 n2_19366_5169 0.0
V23868 n0_19366_5202 n2_19366_5202 0.0
V23869 n0_19366_5239 n2_19366_5239 0.0
V23870 n0_19366_5385 n2_19366_5385 0.0
V23871 n0_19366_5418 n2_19366_5418 0.0
V23872 n0_19366_5455 n2_19366_5455 0.0
V23873 n0_19366_5601 n2_19366_5601 0.0
V23874 n0_19366_5634 n2_19366_5634 0.0
V23875 n0_19366_5671 n2_19366_5671 0.0
V23876 n0_19366_5817 n2_19366_5817 0.0
V23877 n0_19366_5850 n2_19366_5850 0.0
V23878 n0_19366_6033 n2_19366_6033 0.0
V23879 n0_19366_6066 n2_19366_6066 0.0
V23880 n0_19366_6249 n2_19366_6249 0.0
V23881 n0_19366_6282 n2_19366_6282 0.0
V23882 n0_19366_6319 n2_19366_6319 0.0
V23883 n0_19366_6465 n2_19366_6465 0.0
V23884 n0_19366_6498 n2_19366_6498 0.0
V23885 n0_19366_6681 n2_19366_6681 0.0
V23886 n0_19366_6714 n2_19366_6714 0.0
V23887 n0_19366_6897 n2_19366_6897 0.0
V23888 n0_19366_6930 n2_19366_6930 0.0
V23889 n0_19366_7113 n2_19366_7113 0.0
V23890 n0_19366_7146 n2_19366_7146 0.0
V23891 n0_19366_7329 n2_19366_7329 0.0
V23892 n0_19366_7362 n2_19366_7362 0.0
V23893 n0_19366_7545 n2_19366_7545 0.0
V23894 n0_19366_7578 n2_19366_7578 0.0
V23895 n0_19366_7761 n2_19366_7761 0.0
V23896 n0_19366_7794 n2_19366_7794 0.0
V23897 n0_19366_7831 n2_19366_7831 0.0
V23898 n0_19366_7977 n2_19366_7977 0.0
V23899 n0_19366_8010 n2_19366_8010 0.0
V23900 n0_19366_8193 n2_19366_8193 0.0
V23901 n0_19366_8226 n2_19366_8226 0.0
V23902 n0_19366_8409 n2_19366_8409 0.0
V23903 n0_19366_8442 n2_19366_8442 0.0
V23904 n0_19366_8625 n2_19366_8625 0.0
V23905 n0_19366_8658 n2_19366_8658 0.0
V23906 n0_19366_8841 n2_19366_8841 0.0
V23907 n0_19366_8874 n2_19366_8874 0.0
V23908 n0_19366_8911 n2_19366_8911 0.0
V23909 n0_19366_9057 n2_19366_9057 0.0
V23910 n0_19366_9090 n2_19366_9090 0.0
V23911 n0_19366_9273 n2_19366_9273 0.0
V23912 n0_19366_9306 n2_19366_9306 0.0
V23913 n0_19366_9489 n2_19366_9489 0.0
V23914 n0_19366_9522 n2_19366_9522 0.0
V23915 n0_19366_9705 n2_19366_9705 0.0
V23916 n0_19366_9738 n2_19366_9738 0.0
V23917 n0_19366_9921 n2_19366_9921 0.0
V23918 n0_19366_9954 n2_19366_9954 0.0
V23919 n0_19366_9991 n2_19366_9991 0.0
V23920 n0_19366_10137 n2_19366_10137 0.0
V23921 n0_19366_10170 n2_19366_10170 0.0
V23922 n0_19366_10353 n2_19366_10353 0.0
V23923 n0_19366_10386 n2_19366_10386 0.0
V23924 n0_19366_10569 n2_19366_10569 0.0
V23925 n0_19366_10785 n2_19366_10785 0.0
V23926 n0_19366_10818 n2_19366_10818 0.0
V23927 n0_19366_11001 n2_19366_11001 0.0
V23928 n0_19366_11034 n2_19366_11034 0.0
V23929 n0_19366_11055 n2_19366_11055 0.0
V23930 n0_19366_11217 n2_19366_11217 0.0
V23931 n0_19366_11250 n2_19366_11250 0.0
V23932 n0_19366_11433 n2_19366_11433 0.0
V23933 n0_19366_11466 n2_19366_11466 0.0
V23934 n0_19366_11649 n2_19366_11649 0.0
V23935 n0_19366_11682 n2_19366_11682 0.0
V23936 n0_19366_11865 n2_19366_11865 0.0
V23937 n0_19366_11898 n2_19366_11898 0.0
V23938 n0_19366_12081 n2_19366_12081 0.0
V23939 n0_19366_12114 n2_19366_12114 0.0
V23940 n0_19366_12128 n2_19366_12128 0.0
V23941 n0_19366_12297 n2_19366_12297 0.0
V23942 n0_19366_12330 n2_19366_12330 0.0
V23943 n0_19366_12513 n2_19366_12513 0.0
V23944 n0_19366_12546 n2_19366_12546 0.0
V23945 n0_19366_12729 n2_19366_12729 0.0
V23946 n0_19366_12762 n2_19366_12762 0.0
V23947 n0_19366_12945 n2_19366_12945 0.0
V23948 n0_19366_12978 n2_19366_12978 0.0
V23949 n0_19366_13161 n2_19366_13161 0.0
V23950 n0_19366_13194 n2_19366_13194 0.0
V23951 n0_19366_13377 n2_19366_13377 0.0
V23952 n0_19366_13410 n2_19366_13410 0.0
V23953 n0_19366_13593 n2_19366_13593 0.0
V23954 n0_19366_13626 n2_19366_13626 0.0
V23955 n0_19366_13647 n2_19366_13647 0.0
V23956 n0_19366_13809 n2_19366_13809 0.0
V23957 n0_19366_13842 n2_19366_13842 0.0
V23958 n0_19366_14025 n2_19366_14025 0.0
V23959 n0_19366_14058 n2_19366_14058 0.0
V23960 n0_19366_14241 n2_19366_14241 0.0
V23961 n0_19366_14274 n2_19366_14274 0.0
V23962 n0_19366_14457 n2_19366_14457 0.0
V23963 n0_19366_14490 n2_19366_14490 0.0
V23964 n0_19366_14504 n2_19366_14504 0.0
V23965 n0_19366_14511 n2_19366_14511 0.0
V23966 n0_19366_14673 n2_19366_14673 0.0
V23967 n0_19366_14706 n2_19366_14706 0.0
V23968 n0_19366_14889 n2_19366_14889 0.0
V23969 n0_19366_14922 n2_19366_14922 0.0
V23970 n0_19366_14936 n2_19366_14936 0.0
V23971 n0_19366_15138 n2_19366_15138 0.0
V23972 n0_19366_15152 n2_19366_15152 0.0
V23973 n0_19366_15321 n2_19366_15321 0.0
V23974 n0_19366_15354 n2_19366_15354 0.0
V23975 n0_19366_15537 n2_19366_15537 0.0
V23976 n0_19366_15570 n2_19366_15570 0.0
V23977 n0_19366_15584 n2_19366_15584 0.0
V23978 n0_19366_15753 n2_19366_15753 0.0
V23979 n0_19366_15786 n2_19366_15786 0.0
V23980 n0_19366_15969 n2_19366_15969 0.0
V23981 n0_19366_16002 n2_19366_16002 0.0
V23982 n0_19366_16185 n2_19366_16185 0.0
V23983 n0_19366_16218 n2_19366_16218 0.0
V23984 n0_19366_16401 n2_19366_16401 0.0
V23985 n0_19366_16434 n2_19366_16434 0.0
V23986 n0_19366_16617 n2_19366_16617 0.0
V23987 n0_19366_16650 n2_19366_16650 0.0
V23988 n0_19366_16664 n2_19366_16664 0.0
V23989 n0_19366_16671 n2_19366_16671 0.0
V23990 n0_19366_16687 n2_19366_16687 0.0
V23991 n0_19366_16833 n2_19366_16833 0.0
V23992 n0_19366_16866 n2_19366_16866 0.0
V23993 n0_19366_17049 n2_19366_17049 0.0
V23994 n0_19366_17082 n2_19366_17082 0.0
V23995 n0_19366_17119 n2_19366_17119 0.0
V23996 n0_19366_17265 n2_19366_17265 0.0
V23997 n0_19366_17298 n2_19366_17298 0.0
V23998 n0_19366_17481 n2_19366_17481 0.0
V23999 n0_19366_17514 n2_19366_17514 0.0
V24000 n0_19366_17697 n2_19366_17697 0.0
V24001 n0_19366_17730 n2_19366_17730 0.0
V24002 n0_19366_17744 n2_19366_17744 0.0
V24003 n0_19366_17913 n2_19366_17913 0.0
V24004 n0_19366_17946 n2_19366_17946 0.0
V24005 n0_19366_18129 n2_19366_18129 0.0
V24006 n0_19366_18162 n2_19366_18162 0.0
V24007 n0_19366_18345 n2_19366_18345 0.0
V24008 n0_19366_18378 n2_19366_18378 0.0
V24009 n0_19366_18561 n2_19366_18561 0.0
V24010 n0_19366_18594 n2_19366_18594 0.0
V24011 n0_19366_18777 n2_19366_18777 0.0
V24012 n0_19366_18810 n2_19366_18810 0.0
V24013 n0_19366_18932 n2_19366_18932 0.0
V24014 n0_19366_18993 n2_19366_18993 0.0
V24015 n0_19366_19026 n2_19366_19026 0.0
V24016 n0_19366_19040 n2_19366_19040 0.0
V24017 n0_19366_19209 n2_19366_19209 0.0
V24018 n0_19366_19242 n2_19366_19242 0.0
V24019 n0_19366_19425 n2_19366_19425 0.0
V24020 n0_19366_19458 n2_19366_19458 0.0
V24021 n0_19366_19641 n2_19366_19641 0.0
V24022 n0_19366_19674 n2_19366_19674 0.0
V24023 n0_19366_19857 n2_19366_19857 0.0
V24024 n0_19366_19890 n2_19366_19890 0.0
V24025 n0_19366_20073 n2_19366_20073 0.0
V24026 n0_19366_20106 n2_19366_20106 0.0
V24027 n0_19366_20289 n2_19366_20289 0.0
V24028 n0_19366_20322 n2_19366_20322 0.0
V24029 n0_19366_20505 n2_19366_20505 0.0
V24030 n0_19366_20538 n2_19366_20538 0.0
V24031 n0_19366_20754 n2_19366_20754 0.0
V24032 n0_19366_20937 n2_19366_20937 0.0
V24033 n0_19366_20970 n2_19366_20970 0.0
V24034 n0_19458_201 n2_19458_201 0.0
V24035 n0_19458_234 n2_19458_234 0.0
V24036 n0_19458_417 n2_19458_417 0.0
V24037 n0_19458_450 n2_19458_450 0.0
V24038 n0_19458_633 n2_19458_633 0.0
V24039 n0_19458_666 n2_19458_666 0.0
V24040 n0_19458_849 n2_19458_849 0.0
V24041 n0_19458_882 n2_19458_882 0.0
V24042 n0_19458_1065 n2_19458_1065 0.0
V24043 n0_19458_1098 n2_19458_1098 0.0
V24044 n0_19458_1281 n2_19458_1281 0.0
V24045 n0_19458_1314 n2_19458_1314 0.0
V24046 n0_19458_1497 n2_19458_1497 0.0
V24047 n0_19458_19857 n2_19458_19857 0.0
V24048 n0_19458_19890 n2_19458_19890 0.0
V24049 n0_19458_20073 n2_19458_20073 0.0
V24050 n0_19458_20106 n2_19458_20106 0.0
V24051 n0_19458_20289 n2_19458_20289 0.0
V24052 n0_19458_20322 n2_19458_20322 0.0
V24053 n0_19458_20505 n2_19458_20505 0.0
V24054 n0_19458_20538 n2_19458_20538 0.0
V24055 n0_19458_20721 n2_19458_20721 0.0
V24056 n0_19458_20754 n2_19458_20754 0.0
V24057 n0_19458_20937 n2_19458_20937 0.0
V24058 n0_19458_20970 n2_19458_20970 0.0
V24059 n0_19505_417 n2_19505_417 0.0
V24060 n0_19505_450 n2_19505_450 0.0
V24061 n0_19505_3873 n2_19505_3873 0.0
V24062 n0_19505_3906 n2_19505_3906 0.0
V24063 n0_19505_6033 n2_19505_6033 0.0
V24064 n0_19505_6066 n2_19505_6066 0.0
V24065 n0_19505_8409 n2_19505_8409 0.0
V24066 n0_19505_10569 n2_19505_10569 0.0
V24067 n0_19505_10602 n2_19505_10602 0.0
V24068 n0_19505_15105 n2_19505_15105 0.0
V24069 n0_19505_15138 n2_19505_15138 0.0
V24070 n0_19505_15152 n2_19505_15152 0.0
V24071 n0_19505_17298 n2_19505_17298 0.0
V24072 n0_19505_20721 n2_19505_20721 0.0
V24073 n0_19505_20754 n2_19505_20754 0.0
V24074 n0_19554_201 n2_19554_201 0.0
V24075 n0_19554_234 n2_19554_234 0.0
V24076 n0_19554_417 n2_19554_417 0.0
V24077 n0_19554_450 n2_19554_450 0.0
V24078 n0_19554_633 n2_19554_633 0.0
V24079 n0_19554_666 n2_19554_666 0.0
V24080 n0_19554_849 n2_19554_849 0.0
V24081 n0_19554_882 n2_19554_882 0.0
V24082 n0_19554_1065 n2_19554_1065 0.0
V24083 n0_19554_1098 n2_19554_1098 0.0
V24084 n0_19554_1281 n2_19554_1281 0.0
V24085 n0_19554_1314 n2_19554_1314 0.0
V24086 n0_19554_1497 n2_19554_1497 0.0
V24087 n0_19554_1713 n2_19554_1713 0.0
V24088 n0_19554_1746 n2_19554_1746 0.0
V24089 n0_19554_1929 n2_19554_1929 0.0
V24090 n0_19554_1962 n2_19554_1962 0.0
V24091 n0_19554_1976 n2_19554_1976 0.0
V24092 n0_19554_1999 n2_19554_1999 0.0
V24093 n0_19554_2145 n2_19554_2145 0.0
V24094 n0_19554_2178 n2_19554_2178 0.0
V24095 n0_19554_2361 n2_19554_2361 0.0
V24096 n0_19554_2394 n2_19554_2394 0.0
V24097 n0_19554_2577 n2_19554_2577 0.0
V24098 n0_19554_2610 n2_19554_2610 0.0
V24099 n0_19554_2826 n2_19554_2826 0.0
V24100 n0_19554_3009 n2_19554_3009 0.0
V24101 n0_19554_3042 n2_19554_3042 0.0
V24102 n0_19554_3225 n2_19554_3225 0.0
V24103 n0_19554_3258 n2_19554_3258 0.0
V24104 n0_19554_3295 n2_19554_3295 0.0
V24105 n0_19554_3441 n2_19554_3441 0.0
V24106 n0_19554_3474 n2_19554_3474 0.0
V24107 n0_19554_3657 n2_19554_3657 0.0
V24108 n0_19554_3690 n2_19554_3690 0.0
V24109 n0_19554_3873 n2_19554_3873 0.0
V24110 n0_19554_3906 n2_19554_3906 0.0
V24111 n0_19554_4089 n2_19554_4089 0.0
V24112 n0_19554_4122 n2_19554_4122 0.0
V24113 n0_19554_4305 n2_19554_4305 0.0
V24114 n0_19554_4338 n2_19554_4338 0.0
V24115 n0_19554_4375 n2_19554_4375 0.0
V24116 n0_19554_4521 n2_19554_4521 0.0
V24117 n0_19554_4554 n2_19554_4554 0.0
V24118 n0_19554_4737 n2_19554_4737 0.0
V24119 n0_19554_4770 n2_19554_4770 0.0
V24120 n0_19554_5169 n2_19554_5169 0.0
V24121 n0_19554_5202 n2_19554_5202 0.0
V24122 n0_19554_5239 n2_19554_5239 0.0
V24123 n0_19554_5385 n2_19554_5385 0.0
V24124 n0_19554_5418 n2_19554_5418 0.0
V24125 n0_19554_5455 n2_19554_5455 0.0
V24126 n0_19554_5601 n2_19554_5601 0.0
V24127 n0_19554_5634 n2_19554_5634 0.0
V24128 n0_19554_5671 n2_19554_5671 0.0
V24129 n0_19554_5817 n2_19554_5817 0.0
V24130 n0_19554_5850 n2_19554_5850 0.0
V24131 n0_19554_6033 n2_19554_6033 0.0
V24132 n0_19554_6066 n2_19554_6066 0.0
V24133 n0_19554_6249 n2_19554_6249 0.0
V24134 n0_19554_6282 n2_19554_6282 0.0
V24135 n0_19554_6319 n2_19554_6319 0.0
V24136 n0_19554_6465 n2_19554_6465 0.0
V24137 n0_19554_6498 n2_19554_6498 0.0
V24138 n0_19554_6681 n2_19554_6681 0.0
V24139 n0_19554_6714 n2_19554_6714 0.0
V24140 n0_19554_6897 n2_19554_6897 0.0
V24141 n0_19554_6930 n2_19554_6930 0.0
V24142 n0_19554_7113 n2_19554_7113 0.0
V24143 n0_19554_7329 n2_19554_7329 0.0
V24144 n0_19554_7362 n2_19554_7362 0.0
V24145 n0_19554_7545 n2_19554_7545 0.0
V24146 n0_19554_7578 n2_19554_7578 0.0
V24147 n0_19554_7761 n2_19554_7761 0.0
V24148 n0_19554_7794 n2_19554_7794 0.0
V24149 n0_19554_7831 n2_19554_7831 0.0
V24150 n0_19554_7977 n2_19554_7977 0.0
V24151 n0_19554_8010 n2_19554_8010 0.0
V24152 n0_19554_8193 n2_19554_8193 0.0
V24153 n0_19554_8226 n2_19554_8226 0.0
V24154 n0_19554_8409 n2_19554_8409 0.0
V24155 n0_19554_8442 n2_19554_8442 0.0
V24156 n0_19554_8625 n2_19554_8625 0.0
V24157 n0_19554_8658 n2_19554_8658 0.0
V24158 n0_19554_8841 n2_19554_8841 0.0
V24159 n0_19554_8874 n2_19554_8874 0.0
V24160 n0_19554_8911 n2_19554_8911 0.0
V24161 n0_19554_9057 n2_19554_9057 0.0
V24162 n0_19554_9090 n2_19554_9090 0.0
V24163 n0_19554_9273 n2_19554_9273 0.0
V24164 n0_19554_9306 n2_19554_9306 0.0
V24165 n0_19554_9705 n2_19554_9705 0.0
V24166 n0_19554_9738 n2_19554_9738 0.0
V24167 n0_19554_9921 n2_19554_9921 0.0
V24168 n0_19554_9954 n2_19554_9954 0.0
V24169 n0_19554_9991 n2_19554_9991 0.0
V24170 n0_19554_10137 n2_19554_10137 0.0
V24171 n0_19554_10170 n2_19554_10170 0.0
V24172 n0_19554_10353 n2_19554_10353 0.0
V24173 n0_19554_10386 n2_19554_10386 0.0
V24174 n0_19554_10569 n2_19554_10569 0.0
V24175 n0_19554_10602 n2_19554_10602 0.0
V24176 n0_19554_10785 n2_19554_10785 0.0
V24177 n0_19554_10818 n2_19554_10818 0.0
V24178 n0_19554_11001 n2_19554_11001 0.0
V24179 n0_19554_11034 n2_19554_11034 0.0
V24180 n0_19554_11055 n2_19554_11055 0.0
V24181 n0_19554_11217 n2_19554_11217 0.0
V24182 n0_19554_11250 n2_19554_11250 0.0
V24183 n0_19554_11433 n2_19554_11433 0.0
V24184 n0_19554_11466 n2_19554_11466 0.0
V24185 n0_19554_11865 n2_19554_11865 0.0
V24186 n0_19554_11898 n2_19554_11898 0.0
V24187 n0_19554_12081 n2_19554_12081 0.0
V24188 n0_19554_12114 n2_19554_12114 0.0
V24189 n0_19554_12128 n2_19554_12128 0.0
V24190 n0_19554_12297 n2_19554_12297 0.0
V24191 n0_19554_12330 n2_19554_12330 0.0
V24192 n0_19554_12513 n2_19554_12513 0.0
V24193 n0_19554_12546 n2_19554_12546 0.0
V24194 n0_19554_12729 n2_19554_12729 0.0
V24195 n0_19554_12762 n2_19554_12762 0.0
V24196 n0_19554_12945 n2_19554_12945 0.0
V24197 n0_19554_12978 n2_19554_12978 0.0
V24198 n0_19554_13161 n2_19554_13161 0.0
V24199 n0_19554_13194 n2_19554_13194 0.0
V24200 n0_19554_13377 n2_19554_13377 0.0
V24201 n0_19554_13410 n2_19554_13410 0.0
V24202 n0_19554_13593 n2_19554_13593 0.0
V24203 n0_19554_13626 n2_19554_13626 0.0
V24204 n0_19554_13647 n2_19554_13647 0.0
V24205 n0_19554_13809 n2_19554_13809 0.0
V24206 n0_19554_13842 n2_19554_13842 0.0
V24207 n0_19554_14241 n2_19554_14241 0.0
V24208 n0_19554_14274 n2_19554_14274 0.0
V24209 n0_19554_14457 n2_19554_14457 0.0
V24210 n0_19554_14490 n2_19554_14490 0.0
V24211 n0_19554_14504 n2_19554_14504 0.0
V24212 n0_19554_14511 n2_19554_14511 0.0
V24213 n0_19554_14673 n2_19554_14673 0.0
V24214 n0_19554_14706 n2_19554_14706 0.0
V24215 n0_19554_14889 n2_19554_14889 0.0
V24216 n0_19554_14922 n2_19554_14922 0.0
V24217 n0_19554_14936 n2_19554_14936 0.0
V24218 n0_19554_15105 n2_19554_15105 0.0
V24219 n0_19554_15138 n2_19554_15138 0.0
V24220 n0_19554_15152 n2_19554_15152 0.0
V24221 n0_19554_15321 n2_19554_15321 0.0
V24222 n0_19554_15354 n2_19554_15354 0.0
V24223 n0_19554_15537 n2_19554_15537 0.0
V24224 n0_19554_15570 n2_19554_15570 0.0
V24225 n0_19554_15584 n2_19554_15584 0.0
V24226 n0_19554_15753 n2_19554_15753 0.0
V24227 n0_19554_15786 n2_19554_15786 0.0
V24228 n0_19554_15969 n2_19554_15969 0.0
V24229 n0_19554_16002 n2_19554_16002 0.0
V24230 n0_19554_16401 n2_19554_16401 0.0
V24231 n0_19554_16434 n2_19554_16434 0.0
V24232 n0_19554_16617 n2_19554_16617 0.0
V24233 n0_19554_16650 n2_19554_16650 0.0
V24234 n0_19554_16664 n2_19554_16664 0.0
V24235 n0_19554_16671 n2_19554_16671 0.0
V24236 n0_19554_16687 n2_19554_16687 0.0
V24237 n0_19554_16833 n2_19554_16833 0.0
V24238 n0_19554_16866 n2_19554_16866 0.0
V24239 n0_19554_17049 n2_19554_17049 0.0
V24240 n0_19554_17082 n2_19554_17082 0.0
V24241 n0_19554_17119 n2_19554_17119 0.0
V24242 n0_19554_17265 n2_19554_17265 0.0
V24243 n0_19554_17298 n2_19554_17298 0.0
V24244 n0_19554_17481 n2_19554_17481 0.0
V24245 n0_19554_17514 n2_19554_17514 0.0
V24246 n0_19554_17697 n2_19554_17697 0.0
V24247 n0_19554_17730 n2_19554_17730 0.0
V24248 n0_19554_17744 n2_19554_17744 0.0
V24249 n0_19554_17913 n2_19554_17913 0.0
V24250 n0_19554_17946 n2_19554_17946 0.0
V24251 n0_19554_18129 n2_19554_18129 0.0
V24252 n0_19554_18162 n2_19554_18162 0.0
V24253 n0_19554_18345 n2_19554_18345 0.0
V24254 n0_19554_18594 n2_19554_18594 0.0
V24255 n0_19554_18777 n2_19554_18777 0.0
V24256 n0_19554_18810 n2_19554_18810 0.0
V24257 n0_19554_18932 n2_19554_18932 0.0
V24258 n0_19554_18993 n2_19554_18993 0.0
V24259 n0_19554_19026 n2_19554_19026 0.0
V24260 n0_19554_19040 n2_19554_19040 0.0
V24261 n0_19554_19209 n2_19554_19209 0.0
V24262 n0_19554_19242 n2_19554_19242 0.0
V24263 n0_19554_19425 n2_19554_19425 0.0
V24264 n0_19554_19458 n2_19554_19458 0.0
V24265 n0_19554_19857 n2_19554_19857 0.0
V24266 n0_19554_19890 n2_19554_19890 0.0
V24267 n0_19554_20073 n2_19554_20073 0.0
V24268 n0_19554_20106 n2_19554_20106 0.0
V24269 n0_19554_20289 n2_19554_20289 0.0
V24270 n0_19554_20322 n2_19554_20322 0.0
V24271 n0_19554_20505 n2_19554_20505 0.0
V24272 n0_19554_20538 n2_19554_20538 0.0
V24273 n0_19554_20721 n2_19554_20721 0.0
V24274 n0_19554_20754 n2_19554_20754 0.0
V24275 n0_19554_20937 n2_19554_20937 0.0
V24276 n0_19554_20970 n2_19554_20970 0.0
V24277 n0_19646_201 n2_19646_201 0.0
V24278 n0_19646_234 n2_19646_234 0.0
V24279 n0_19646_417 n2_19646_417 0.0
V24280 n0_19646_450 n2_19646_450 0.0
V24281 n0_19646_633 n2_19646_633 0.0
V24282 n0_19646_666 n2_19646_666 0.0
V24283 n0_19646_849 n2_19646_849 0.0
V24284 n0_19646_882 n2_19646_882 0.0
V24285 n0_19646_1065 n2_19646_1065 0.0
V24286 n0_19646_1098 n2_19646_1098 0.0
V24287 n0_19646_1281 n2_19646_1281 0.0
V24288 n0_19646_1314 n2_19646_1314 0.0
V24289 n0_19646_1497 n2_19646_1497 0.0
V24290 n0_19646_1530 n2_19646_1530 0.0
V24291 n0_19646_19641 n2_19646_19641 0.0
V24292 n0_19646_19674 n2_19646_19674 0.0
V24293 n0_19646_19857 n2_19646_19857 0.0
V24294 n0_19646_19890 n2_19646_19890 0.0
V24295 n0_19646_20073 n2_19646_20073 0.0
V24296 n0_19646_20106 n2_19646_20106 0.0
V24297 n0_19646_20289 n2_19646_20289 0.0
V24298 n0_19646_20322 n2_19646_20322 0.0
V24299 n0_19646_20505 n2_19646_20505 0.0
V24300 n0_19646_20538 n2_19646_20538 0.0
V24301 n0_19646_20754 n2_19646_20754 0.0
V24302 n0_19646_20937 n2_19646_20937 0.0
V24303 n0_19646_20970 n2_19646_20970 0.0
V24304 n0_20491_633 n2_20491_633 0.0
V24305 n0_20491_666 n2_20491_666 0.0
V24306 n0_20491_849 n2_20491_849 0.0
V24307 n0_20491_882 n2_20491_882 0.0
V24308 n0_20491_1065 n2_20491_1065 0.0
V24309 n0_20491_1098 n2_20491_1098 0.0
V24310 n0_20491_1281 n2_20491_1281 0.0
V24311 n0_20491_1314 n2_20491_1314 0.0
V24312 n0_20491_1497 n2_20491_1497 0.0
V24313 n0_20491_1530 n2_20491_1530 0.0
V24314 n0_20491_1713 n2_20491_1713 0.0
V24315 n0_20491_1746 n2_20491_1746 0.0
V24316 n0_20491_1929 n2_20491_1929 0.0
V24317 n0_20491_1962 n2_20491_1962 0.0
V24318 n0_20491_1976 n2_20491_1976 0.0
V24319 n0_20491_2145 n2_20491_2145 0.0
V24320 n0_20491_2178 n2_20491_2178 0.0
V24321 n0_20491_2361 n2_20491_2361 0.0
V24322 n0_20491_2394 n2_20491_2394 0.0
V24323 n0_20491_2577 n2_20491_2577 0.0
V24324 n0_20491_2610 n2_20491_2610 0.0
V24325 n0_20491_2793 n2_20491_2793 0.0
V24326 n0_20491_2826 n2_20491_2826 0.0
V24327 n0_20491_3009 n2_20491_3009 0.0
V24328 n0_20491_3042 n2_20491_3042 0.0
V24329 n0_20491_3225 n2_20491_3225 0.0
V24330 n0_20491_3258 n2_20491_3258 0.0
V24331 n0_20491_3441 n2_20491_3441 0.0
V24332 n0_20491_3474 n2_20491_3474 0.0
V24333 n0_20491_3657 n2_20491_3657 0.0
V24334 n0_20491_3690 n2_20491_3690 0.0
V24335 n0_20491_3873 n2_20491_3873 0.0
V24336 n0_20491_3906 n2_20491_3906 0.0
V24337 n0_20491_4089 n2_20491_4089 0.0
V24338 n0_20491_4122 n2_20491_4122 0.0
V24339 n0_20491_4305 n2_20491_4305 0.0
V24340 n0_20491_4338 n2_20491_4338 0.0
V24341 n0_20491_4521 n2_20491_4521 0.0
V24342 n0_20491_4554 n2_20491_4554 0.0
V24343 n0_20491_4737 n2_20491_4737 0.0
V24344 n0_20491_4770 n2_20491_4770 0.0
V24345 n0_20491_4953 n2_20491_4953 0.0
V24346 n0_20491_4986 n2_20491_4986 0.0
V24347 n0_20491_5169 n2_20491_5169 0.0
V24348 n0_20491_5202 n2_20491_5202 0.0
V24349 n0_20491_5385 n2_20491_5385 0.0
V24350 n0_20491_5418 n2_20491_5418 0.0
V24351 n0_20491_5601 n2_20491_5601 0.0
V24352 n0_20491_5634 n2_20491_5634 0.0
V24353 n0_20491_5671 n2_20491_5671 0.0
V24354 n0_20491_5817 n2_20491_5817 0.0
V24355 n0_20491_5850 n2_20491_5850 0.0
V24356 n0_20491_6033 n2_20491_6033 0.0
V24357 n0_20491_6066 n2_20491_6066 0.0
V24358 n0_20491_6249 n2_20491_6249 0.0
V24359 n0_20491_6282 n2_20491_6282 0.0
V24360 n0_20491_6319 n2_20491_6319 0.0
V24361 n0_20491_6465 n2_20491_6465 0.0
V24362 n0_20491_6498 n2_20491_6498 0.0
V24363 n0_20491_6681 n2_20491_6681 0.0
V24364 n0_20491_6714 n2_20491_6714 0.0
V24365 n0_20491_6897 n2_20491_6897 0.0
V24366 n0_20491_6930 n2_20491_6930 0.0
V24367 n0_20491_7113 n2_20491_7113 0.0
V24368 n0_20491_7146 n2_20491_7146 0.0
V24369 n0_20491_7329 n2_20491_7329 0.0
V24370 n0_20491_7362 n2_20491_7362 0.0
V24371 n0_20491_7545 n2_20491_7545 0.0
V24372 n0_20491_7578 n2_20491_7578 0.0
V24373 n0_20491_7761 n2_20491_7761 0.0
V24374 n0_20491_7794 n2_20491_7794 0.0
V24375 n0_20491_7977 n2_20491_7977 0.0
V24376 n0_20491_8010 n2_20491_8010 0.0
V24377 n0_20491_8193 n2_20491_8193 0.0
V24378 n0_20491_8226 n2_20491_8226 0.0
V24379 n0_20491_8409 n2_20491_8409 0.0
V24380 n0_20491_8442 n2_20491_8442 0.0
V24381 n0_20491_8625 n2_20491_8625 0.0
V24382 n0_20491_8658 n2_20491_8658 0.0
V24383 n0_20491_8841 n2_20491_8841 0.0
V24384 n0_20491_8874 n2_20491_8874 0.0
V24385 n0_20491_9057 n2_20491_9057 0.0
V24386 n0_20491_9090 n2_20491_9090 0.0
V24387 n0_20491_9213 n2_20491_9213 0.0
V24388 n0_20491_11956 n2_20491_11956 0.0
V24389 n0_20491_12081 n2_20491_12081 0.0
V24390 n0_20491_12114 n2_20491_12114 0.0
V24391 n0_20491_12297 n2_20491_12297 0.0
V24392 n0_20491_12330 n2_20491_12330 0.0
V24393 n0_20491_12513 n2_20491_12513 0.0
V24394 n0_20491_12546 n2_20491_12546 0.0
V24395 n0_20491_12729 n2_20491_12729 0.0
V24396 n0_20491_12762 n2_20491_12762 0.0
V24397 n0_20491_12945 n2_20491_12945 0.0
V24398 n0_20491_12978 n2_20491_12978 0.0
V24399 n0_20491_13161 n2_20491_13161 0.0
V24400 n0_20491_13194 n2_20491_13194 0.0
V24401 n0_20491_13377 n2_20491_13377 0.0
V24402 n0_20491_13410 n2_20491_13410 0.0
V24403 n0_20491_13593 n2_20491_13593 0.0
V24404 n0_20491_13626 n2_20491_13626 0.0
V24405 n0_20491_13809 n2_20491_13809 0.0
V24406 n0_20491_13842 n2_20491_13842 0.0
V24407 n0_20491_14025 n2_20491_14025 0.0
V24408 n0_20491_14058 n2_20491_14058 0.0
V24409 n0_20491_14241 n2_20491_14241 0.0
V24410 n0_20491_14274 n2_20491_14274 0.0
V24411 n0_20491_14457 n2_20491_14457 0.0
V24412 n0_20491_14490 n2_20491_14490 0.0
V24413 n0_20491_14673 n2_20491_14673 0.0
V24414 n0_20491_14706 n2_20491_14706 0.0
V24415 n0_20491_14889 n2_20491_14889 0.0
V24416 n0_20491_14922 n2_20491_14922 0.0
V24417 n0_20491_14936 n2_20491_14936 0.0
V24418 n0_20491_15138 n2_20491_15138 0.0
V24419 n0_20491_15152 n2_20491_15152 0.0
V24420 n0_20491_15321 n2_20491_15321 0.0
V24421 n0_20491_15354 n2_20491_15354 0.0
V24422 n0_20491_15537 n2_20491_15537 0.0
V24423 n0_20491_15570 n2_20491_15570 0.0
V24424 n0_20491_15753 n2_20491_15753 0.0
V24425 n0_20491_15786 n2_20491_15786 0.0
V24426 n0_20491_15969 n2_20491_15969 0.0
V24427 n0_20491_16002 n2_20491_16002 0.0
V24428 n0_20491_16185 n2_20491_16185 0.0
V24429 n0_20491_16218 n2_20491_16218 0.0
V24430 n0_20491_16401 n2_20491_16401 0.0
V24431 n0_20491_16434 n2_20491_16434 0.0
V24432 n0_20491_16617 n2_20491_16617 0.0
V24433 n0_20491_16650 n2_20491_16650 0.0
V24434 n0_20491_16687 n2_20491_16687 0.0
V24435 n0_20491_16833 n2_20491_16833 0.0
V24436 n0_20491_16866 n2_20491_16866 0.0
V24437 n0_20491_17049 n2_20491_17049 0.0
V24438 n0_20491_17082 n2_20491_17082 0.0
V24439 n0_20491_17265 n2_20491_17265 0.0
V24440 n0_20491_17298 n2_20491_17298 0.0
V24441 n0_20491_17481 n2_20491_17481 0.0
V24442 n0_20491_17514 n2_20491_17514 0.0
V24443 n0_20491_17697 n2_20491_17697 0.0
V24444 n0_20491_17730 n2_20491_17730 0.0
V24445 n0_20491_17913 n2_20491_17913 0.0
V24446 n0_20491_17946 n2_20491_17946 0.0
V24447 n0_20491_18129 n2_20491_18129 0.0
V24448 n0_20491_18162 n2_20491_18162 0.0
V24449 n0_20491_18345 n2_20491_18345 0.0
V24450 n0_20491_18378 n2_20491_18378 0.0
V24451 n0_20491_18561 n2_20491_18561 0.0
V24452 n0_20491_18594 n2_20491_18594 0.0
V24453 n0_20491_18777 n2_20491_18777 0.0
V24454 n0_20491_18810 n2_20491_18810 0.0
V24455 n0_20491_18993 n2_20491_18993 0.0
V24456 n0_20491_19026 n2_20491_19026 0.0
V24457 n0_20491_19040 n2_20491_19040 0.0
V24458 n0_20491_19209 n2_20491_19209 0.0
V24459 n0_20491_19242 n2_20491_19242 0.0
V24460 n0_20491_19425 n2_20491_19425 0.0
V24461 n0_20491_19458 n2_20491_19458 0.0
V24462 n0_20491_19641 n2_20491_19641 0.0
V24463 n0_20491_19674 n2_20491_19674 0.0
V24464 n0_20491_19857 n2_20491_19857 0.0
V24465 n0_20491_19890 n2_20491_19890 0.0
V24466 n0_20491_20073 n2_20491_20073 0.0
V24467 n0_20491_20106 n2_20491_20106 0.0
V24468 n0_20491_20289 n2_20491_20289 0.0
V24469 n0_20491_20322 n2_20491_20322 0.0
V24470 n0_20491_20505 n2_20491_20505 0.0
V24471 n0_20491_20538 n2_20491_20538 0.0
V24472 n0_20630_1530 n2_20630_1530 0.0
V24473 n0_20630_3873 n2_20630_3873 0.0
V24474 n0_20630_3906 n2_20630_3906 0.0
V24475 n0_20630_6033 n2_20630_6033 0.0
V24476 n0_20630_6066 n2_20630_6066 0.0
V24477 n0_20630_8409 n2_20630_8409 0.0
V24478 n0_20630_15105 n2_20630_15105 0.0
V24479 n0_20630_15138 n2_20630_15138 0.0
V24480 n0_20630_15152 n2_20630_15152 0.0
V24481 n0_20630_17298 n2_20630_17298 0.0
V24482 n0_20630_19641 n2_20630_19641 0.0
V24483 n0_20630_19674 n2_20630_19674 0.0
V24484 n0_20679_633 n2_20679_633 0.0
V24485 n0_20679_666 n2_20679_666 0.0
V24486 n0_20679_849 n2_20679_849 0.0
V24487 n0_20679_882 n2_20679_882 0.0
V24488 n0_20679_1065 n2_20679_1065 0.0
V24489 n0_20679_1098 n2_20679_1098 0.0
V24490 n0_20679_1281 n2_20679_1281 0.0
V24491 n0_20679_1314 n2_20679_1314 0.0
V24492 n0_20679_1497 n2_20679_1497 0.0
V24493 n0_20679_1530 n2_20679_1530 0.0
V24494 n0_20679_1713 n2_20679_1713 0.0
V24495 n0_20679_1746 n2_20679_1746 0.0
V24496 n0_20679_1929 n2_20679_1929 0.0
V24497 n0_20679_1962 n2_20679_1962 0.0
V24498 n0_20679_1976 n2_20679_1976 0.0
V24499 n0_20679_2145 n2_20679_2145 0.0
V24500 n0_20679_2178 n2_20679_2178 0.0
V24501 n0_20679_2361 n2_20679_2361 0.0
V24502 n0_20679_2394 n2_20679_2394 0.0
V24503 n0_20679_2577 n2_20679_2577 0.0
V24504 n0_20679_2610 n2_20679_2610 0.0
V24505 n0_20679_2826 n2_20679_2826 0.0
V24506 n0_20679_3009 n2_20679_3009 0.0
V24507 n0_20679_3042 n2_20679_3042 0.0
V24508 n0_20679_3225 n2_20679_3225 0.0
V24509 n0_20679_3258 n2_20679_3258 0.0
V24510 n0_20679_3441 n2_20679_3441 0.0
V24511 n0_20679_3474 n2_20679_3474 0.0
V24512 n0_20679_3657 n2_20679_3657 0.0
V24513 n0_20679_3690 n2_20679_3690 0.0
V24514 n0_20679_3873 n2_20679_3873 0.0
V24515 n0_20679_3906 n2_20679_3906 0.0
V24516 n0_20679_4089 n2_20679_4089 0.0
V24517 n0_20679_4122 n2_20679_4122 0.0
V24518 n0_20679_4305 n2_20679_4305 0.0
V24519 n0_20679_4338 n2_20679_4338 0.0
V24520 n0_20679_4521 n2_20679_4521 0.0
V24521 n0_20679_4554 n2_20679_4554 0.0
V24522 n0_20679_4737 n2_20679_4737 0.0
V24523 n0_20679_4770 n2_20679_4770 0.0
V24524 n0_20679_5169 n2_20679_5169 0.0
V24525 n0_20679_5202 n2_20679_5202 0.0
V24526 n0_20679_5385 n2_20679_5385 0.0
V24527 n0_20679_5418 n2_20679_5418 0.0
V24528 n0_20679_5601 n2_20679_5601 0.0
V24529 n0_20679_5634 n2_20679_5634 0.0
V24530 n0_20679_5671 n2_20679_5671 0.0
V24531 n0_20679_5817 n2_20679_5817 0.0
V24532 n0_20679_5850 n2_20679_5850 0.0
V24533 n0_20679_6033 n2_20679_6033 0.0
V24534 n0_20679_6066 n2_20679_6066 0.0
V24535 n0_20679_6249 n2_20679_6249 0.0
V24536 n0_20679_6282 n2_20679_6282 0.0
V24537 n0_20679_6319 n2_20679_6319 0.0
V24538 n0_20679_6465 n2_20679_6465 0.0
V24539 n0_20679_6498 n2_20679_6498 0.0
V24540 n0_20679_6681 n2_20679_6681 0.0
V24541 n0_20679_6714 n2_20679_6714 0.0
V24542 n0_20679_6897 n2_20679_6897 0.0
V24543 n0_20679_6930 n2_20679_6930 0.0
V24544 n0_20679_7113 n2_20679_7113 0.0
V24545 n0_20679_7329 n2_20679_7329 0.0
V24546 n0_20679_7362 n2_20679_7362 0.0
V24547 n0_20679_7545 n2_20679_7545 0.0
V24548 n0_20679_7578 n2_20679_7578 0.0
V24549 n0_20679_7761 n2_20679_7761 0.0
V24550 n0_20679_7794 n2_20679_7794 0.0
V24551 n0_20679_7977 n2_20679_7977 0.0
V24552 n0_20679_8010 n2_20679_8010 0.0
V24553 n0_20679_8193 n2_20679_8193 0.0
V24554 n0_20679_8226 n2_20679_8226 0.0
V24555 n0_20679_8409 n2_20679_8409 0.0
V24556 n0_20679_8442 n2_20679_8442 0.0
V24557 n0_20679_8625 n2_20679_8625 0.0
V24558 n0_20679_8658 n2_20679_8658 0.0
V24559 n0_20679_8841 n2_20679_8841 0.0
V24560 n0_20679_8874 n2_20679_8874 0.0
V24561 n0_20679_9057 n2_20679_9057 0.0
V24562 n0_20679_9090 n2_20679_9090 0.0
V24563 n0_20679_9213 n2_20679_9213 0.0
V24564 n0_20679_11956 n2_20679_11956 0.0
V24565 n0_20679_12081 n2_20679_12081 0.0
V24566 n0_20679_12114 n2_20679_12114 0.0
V24567 n0_20679_12297 n2_20679_12297 0.0
V24568 n0_20679_12330 n2_20679_12330 0.0
V24569 n0_20679_12513 n2_20679_12513 0.0
V24570 n0_20679_12546 n2_20679_12546 0.0
V24571 n0_20679_12729 n2_20679_12729 0.0
V24572 n0_20679_12762 n2_20679_12762 0.0
V24573 n0_20679_12945 n2_20679_12945 0.0
V24574 n0_20679_12978 n2_20679_12978 0.0
V24575 n0_20679_13161 n2_20679_13161 0.0
V24576 n0_20679_13194 n2_20679_13194 0.0
V24577 n0_20679_13377 n2_20679_13377 0.0
V24578 n0_20679_13410 n2_20679_13410 0.0
V24579 n0_20679_13593 n2_20679_13593 0.0
V24580 n0_20679_13626 n2_20679_13626 0.0
V24581 n0_20679_13809 n2_20679_13809 0.0
V24582 n0_20679_13842 n2_20679_13842 0.0
V24583 n0_20679_14241 n2_20679_14241 0.0
V24584 n0_20679_14274 n2_20679_14274 0.0
V24585 n0_20679_14457 n2_20679_14457 0.0
V24586 n0_20679_14490 n2_20679_14490 0.0
V24587 n0_20679_14673 n2_20679_14673 0.0
V24588 n0_20679_14706 n2_20679_14706 0.0
V24589 n0_20679_14889 n2_20679_14889 0.0
V24590 n0_20679_14922 n2_20679_14922 0.0
V24591 n0_20679_14936 n2_20679_14936 0.0
V24592 n0_20679_15105 n2_20679_15105 0.0
V24593 n0_20679_15138 n2_20679_15138 0.0
V24594 n0_20679_15152 n2_20679_15152 0.0
V24595 n0_20679_15321 n2_20679_15321 0.0
V24596 n0_20679_15354 n2_20679_15354 0.0
V24597 n0_20679_15537 n2_20679_15537 0.0
V24598 n0_20679_15570 n2_20679_15570 0.0
V24599 n0_20679_15753 n2_20679_15753 0.0
V24600 n0_20679_15786 n2_20679_15786 0.0
V24601 n0_20679_15969 n2_20679_15969 0.0
V24602 n0_20679_16002 n2_20679_16002 0.0
V24603 n0_20679_16401 n2_20679_16401 0.0
V24604 n0_20679_16434 n2_20679_16434 0.0
V24605 n0_20679_16617 n2_20679_16617 0.0
V24606 n0_20679_16650 n2_20679_16650 0.0
V24607 n0_20679_16687 n2_20679_16687 0.0
V24608 n0_20679_16833 n2_20679_16833 0.0
V24609 n0_20679_16866 n2_20679_16866 0.0
V24610 n0_20679_17049 n2_20679_17049 0.0
V24611 n0_20679_17082 n2_20679_17082 0.0
V24612 n0_20679_17265 n2_20679_17265 0.0
V24613 n0_20679_17298 n2_20679_17298 0.0
V24614 n0_20679_17481 n2_20679_17481 0.0
V24615 n0_20679_17514 n2_20679_17514 0.0
V24616 n0_20679_17697 n2_20679_17697 0.0
V24617 n0_20679_17730 n2_20679_17730 0.0
V24618 n0_20679_17913 n2_20679_17913 0.0
V24619 n0_20679_17946 n2_20679_17946 0.0
V24620 n0_20679_18129 n2_20679_18129 0.0
V24621 n0_20679_18162 n2_20679_18162 0.0
V24622 n0_20679_18345 n2_20679_18345 0.0
V24623 n0_20679_18594 n2_20679_18594 0.0
V24624 n0_20679_18777 n2_20679_18777 0.0
V24625 n0_20679_18810 n2_20679_18810 0.0
V24626 n0_20679_18993 n2_20679_18993 0.0
V24627 n0_20679_19026 n2_20679_19026 0.0
V24628 n0_20679_19040 n2_20679_19040 0.0
V24629 n0_20679_19209 n2_20679_19209 0.0
V24630 n0_20679_19242 n2_20679_19242 0.0
V24631 n0_20679_19425 n2_20679_19425 0.0
V24632 n0_20679_19458 n2_20679_19458 0.0
V24633 n0_20679_19641 n2_20679_19641 0.0
V24634 n0_20679_19674 n2_20679_19674 0.0
V24635 n0_20679_19857 n2_20679_19857 0.0
V24636 n0_20679_19890 n2_20679_19890 0.0
V24637 n0_20679_20073 n2_20679_20073 0.0
V24638 n0_20679_20106 n2_20679_20106 0.0
V24639 n0_20679_20289 n2_20679_20289 0.0
V24640 n0_20679_20322 n2_20679_20322 0.0
V24641 n0_20679_20505 n2_20679_20505 0.0
V24642 n0_20679_20538 n2_20679_20538 0.0
v153 _X_n2_1505_6096 0 0
v5d _X_n2_8255_18471 0 0
v155 _X_n2_2630_6096 0 0
v10b _X_n2_3755_471 0 0
v5f _X_n2_8255_17346 0 0
v157 _X_n2_3755_6096 0 0
v10d _X_n2_3755_1596 0 0
v159 _X_n2_4880_6096 0 0
v10f _X_n2_3755_2721 0 0
v161 _X_n2_380_1596 0 0
v6b _X_n2_6005_18471 0 0
v163 _X_n3_9380_20721 0 1.8
v6d _X_n2_6005_17346 0 0
v165 _X_n3_9380_18471 0 1.8
v11b _X_n2_6005_4971 0 0
v6f _X_n2_6005_16221 0 0
v167 _X_n3_9380_16221 0 1.8
v11d _X_n2_6005_6096 0 0
v169 _X_n3_9380_13971 0 1.8
v11f _X_n2_8255_471 0 0
v171 _X_n3_4880_20721 0 1.8
v7b _X_n2_380_17346 0 0
v173 _X_n3_4880_18471 0 1.8
v7d _X_n2_1505_17346 0 0
v175 _X_n3_2630_20721 0 1.8
v12b _X_n2_8255_7221 0 0
v7f _X_n2_2630_17346 0 0
rra0 n2_1505_10596 _X_n2_1505_10596 2.500000e-01
v177 _X_n3_380_20721 0 1.8
v12d _X_n2_8255_8346 0 0
rra2 n2_2630_10596 _X_n2_2630_10596 2.500000e-01
v179 _X_n3_380_18471 0 1.8
v12f _X_n2_10505_471 0 0
rra4 n2_3755_10596 _X_n2_3755_10596 2.500000e-01
v181 _X_n3_4880_16221 0 1.8
v8b _X_n2_4880_15096 0 0
* vias from: 3 to 3
rra6 n2_4880_10596 _X_n2_4880_10596 2.500000e-01
v183 _X_n3_380_13971 0 1.8
v8d _X_n2_6005_15096 0 0
rra8 n2_6005_10596 _X_n2_6005_10596 2.500000e-01
v185 _X_n3_2630_13971 0 1.8
v13b _X_n2_10505_7221 0 0
v8f _X_n2_380_12846 0 0
rrb0 n2_12755_471 _X_n2_12755_471 2.500000e-01
v187 _X_n3_4880_13971 0 1.8
v13d _X_n2_10505_8346 0 0
rrb2 n2_12755_1596 _X_n2_12755_1596 2.500000e-01
iB33_0_v n1_16083_15983 0  0.0218725 
iB33_0_g 0 n0_15991_15969  0.0218725 
iB33_1_v n1_16083_16016 0  0.0218725 
iB33_1_g 0 n0_15991_16002  0.0218725 
iB33_2_v n1_16083_16199 0  0.0218725 
iB33_2_g 0 n0_15991_16185  0.0218725 
iB33_3_v n1_16083_16232 0  0.0218725 
iB33_3_g 0 n0_15991_16185  0.0218725 
iB33_4_v n1_16130_16199 0  0.0218725 
iB33_4_g 0 n0_15991_16185  0.0218725 
iB33_5_v n1_16130_16232 0  0.0218725 
iB33_5_g 0 n0_15991_16185  0.0218725 
iB33_6_v n1_16083_16415 0  0.0218725 
iB33_6_g 0 n0_15991_16185  0.0218725 
iB33_7_v n1_16083_16448 0  0.0218725 
iB33_7_g 0 n0_15991_16185  0.0218725 
iB33_8_v n1_16083_16604 0  0.0218725 
iB33_8_g 0 n0_15991_16185  0.0218725 
iB33_9_v n1_16083_16631 0  0.0218725 
iB33_9_g 0 n0_15991_16185  0.0218725 
iB33_10_v n1_16083_16664 0  0.0218725 
iB33_10_g 0 n0_15991_16185  0.0218725 
iB33_11_v n1_16083_16798 0  0.0218725 
iB33_11_g 0 n0_15991_16185  0.0218725 
iB33_12_v n1_16083_16820 0  0.0218725 
iB33_12_g 0 n0_15991_16185  0.0218725 
iB33_13_v n1_16083_16847 0  0.0218725 
iB33_13_g 0 n0_15991_16185  0.0218725 
iB33_14_v n1_16083_16880 0  0.0218725 
iB33_14_g 0 n0_15991_16185  0.0218725 
iB33_15_v n1_16083_17063 0  0.0218725 
iB33_15_g 0 n0_15146_17049  0.0218725 
iB33_16_v n1_16083_17096 0  0.0218725 
iB33_16_g 0 n0_15146_17096  0.0218725 
iB33_17_v n1_16083_17495 0  0.0218725 
iB33_17_g 0 n0_15146_17481  0.0218725 
iB33_18_v n1_16083_17528 0  0.0218725 
iB33_18_g 0 n0_15146_17528  0.0218725 
iB33_19_v n1_16083_17676 0  0.0218725 
iB33_19_g 0 n0_15146_17697  0.0218725 
iB33_20_v n1_16083_17684 0  0.0218725 
iB33_20_g 0 n0_15146_17697  0.0218725 
iB33_21_v n1_16083_17711 0  0.0218725 
iB33_21_g 0 n0_15146_17697  0.0218725 
iB33_22_v n1_16083_17744 0  0.0218725 
iB33_22_g 0 n0_15146_17730  0.0218725 
iB33_23_v n1_16083_17927 0  0.0218725 
iB33_23_g 0 n0_15146_17913  0.0218725 
iB33_24_v n1_16083_17960 0  0.0218725 
iB33_24_g 0 n0_15146_17946  0.0218725 
iB33_25_v n1_16083_18143 0  0.0218725 
iB33_25_g 0 n0_15146_18129  0.0218725 
iB33_26_v n1_16083_18176 0  0.0218725 
iB33_26_g 0 n0_15146_18176  0.0218725 
iB33_27_v n1_16083_18332 0  0.0218725 
iB33_27_g 0 n0_15146_18345  0.0218725 
iB33_28_v n1_16083_18359 0  0.0218725 
iB33_28_g 0 n0_15146_18345  0.0218725 
iB33_29_v n1_16083_18392 0  0.0218725 
iB33_29_g 0 n0_15146_18378  0.0218725 
iB33_30_v n1_16083_18527 0  0.0218725 
iB33_30_g 0 n0_15146_18561  0.0218725 
iB33_31_v n1_16083_18575 0  0.0218725 
iB33_31_g 0 n0_15146_18561  0.0218725 
iB33_32_v n1_16083_18608 0  0.0218725 
iB33_32_g 0 n0_15146_18608  0.0218725 
iB33_33_v n1_16130_18392 0  0.0218725 
iB33_33_g 0 n0_17116_18378  0.0218725 
iB33_34_v n1_16130_18527 0  0.0218725 
iB33_34_g 0 n0_17116_18561  0.0218725 
iB33_35_v n1_16083_18764 0  0.0218725 
iB33_35_g 0 n0_15146_18777  0.0218725 
iB33_36_v n1_16083_18791 0  0.0218725 
iB33_36_g 0 n0_15146_18777  0.0218725 
iB33_37_v n1_16083_18824 0  0.0218725 
iB33_37_g 0 n0_15146_18810  0.0218725 
iB33_38_v n1_16083_19007 0  0.0218725 
iB33_38_g 0 n0_15146_18993  0.0218725 
iB33_39_v n1_16083_19040 0  0.0218725 
iB33_39_g 0 n0_15146_19026  0.0218725 
iB33_40_v n1_16083_19196 0  0.0218725 
iB33_40_g 0 n0_15146_19209  0.0218725 
iB33_41_v n1_16083_19223 0  0.0218725 
iB33_41_g 0 n0_15146_19209  0.0218725 
iB33_42_v n1_16083_19256 0  0.0218725 
iB33_42_g 0 n0_15146_19256  0.0218725 
iB33_43_v n1_16083_19412 0  0.0218725 
iB33_43_g 0 n0_15146_19425  0.0218725 
iB33_44_v n1_16083_19439 0  0.0218725 
iB33_44_g 0 n0_15146_19425  0.0218725 
iB33_45_v n1_16083_19472 0  0.0218725 
iB33_45_g 0 n0_15146_19458  0.0218725 
iB33_46_v n1_16083_19871 0  0.0218725 
iB33_46_g 0 n0_15146_19857  0.0218725 
iB33_47_v n1_16083_19904 0  0.0218725 
iB33_47_g 0 n0_15146_19890  0.0218725 
iB33_48_v n1_16083_20087 0  0.0218725 
iB33_48_g 0 n0_15146_20073  0.0218725 
iB33_49_v n1_16083_20120 0  0.0218725 
iB33_49_g 0 n0_15146_20106  0.0218725 
iB33_50_v n1_16083_20303 0  0.0218725 
iB33_50_g 0 n0_15146_20289  0.0218725 
iB33_51_v n1_16083_20336 0  0.0218725 
iB33_51_g 0 n0_15146_20322  0.0218725 
iB33_52_v n1_16083_20519 0  0.0218725 
iB33_52_g 0 n0_15146_20505  0.0218725 
iB33_53_v n1_16083_20552 0  0.0218725 
iB33_53_g 0 n0_15146_20538  0.0218725 
iB33_54_v n1_16083_20687 0  0.0218725 
iB33_54_g 0 n0_15146_20754  0.0218725 
iB33_55_v n1_16083_20735 0  0.0218725 
iB33_55_g 0 n0_15146_20754  0.0218725 
iB33_56_v n1_16083_20768 0  0.0218725 
iB33_56_g 0 n0_15146_20754  0.0218725 
iB33_57_v n1_16130_20687 0  0.0218725 
iB33_57_g 0 n0_17116_20754  0.0218725 
iB33_58_v n1_16130_20735 0  0.0218725 
iB33_58_g 0 n0_17116_20754  0.0218725 
iB33_59_v n1_16130_20768 0  0.0218725 
iB33_59_g 0 n0_17116_20754  0.0218725 
iB33_60_v n1_16083_20951 0  0.0218725 
iB33_60_g 0 n0_15146_20937  0.0218725 
iB33_61_v n1_16083_20984 0  0.0218725 
iB33_61_g 0 n0_15146_20970  0.0218725 
iB33_62_v n1_16271_15983 0  0.0218725 
iB33_62_g 0 n0_16179_15969  0.0218725 
iB33_63_v n1_16271_16016 0  0.0218725 
iB33_63_g 0 n0_16179_16002  0.0218725 
iB33_64_v n1_16271_16199 0  0.0218725 
iB33_64_g 0 n0_16179_16002  0.0218725 
iB33_65_v n1_16271_16415 0  0.0218725 
iB33_65_g 0 n0_15991_16185  0.0218725 
iB33_66_v n1_16271_16448 0  0.0218725 
iB33_66_g 0 n0_15991_16185  0.0218725 
iB33_67_v n1_16271_16604 0  0.0218725 
iB33_67_g 0 n0_15991_16185  0.0218725 
iB33_68_v n1_16271_16631 0  0.0218725 
iB33_68_g 0 n0_15991_16185  0.0218725 
iB33_69_v n1_16271_16664 0  0.0218725 
iB33_69_g 0 n0_15991_16185  0.0218725 
iB33_70_v n1_16271_16798 0  0.0218725 
iB33_70_g 0 n0_15991_16185  0.0218725 
iB33_71_v n1_16271_16820 0  0.0218725 
iB33_71_g 0 n0_15991_16185  0.0218725 
iB33_72_v n1_16271_16847 0  0.0218725 
iB33_72_g 0 n0_15991_16185  0.0218725 
iB33_73_v n1_16271_16880 0  0.0218725 
iB33_73_g 0 n0_15991_16185  0.0218725 
iB33_74_v n1_16271_17063 0  0.0218725 
iB33_74_g 0 n0_17116_17049  0.0218725 
iB33_75_v n1_16271_17096 0  0.0218725 
iB33_75_g 0 n0_17116_17082  0.0218725 
iB33_76_v n1_16271_17252 0  0.0218725 
iB33_76_g 0 n0_17116_17265  0.0218725 
iB33_77_v n1_16271_17279 0  0.0218725 
iB33_77_g 0 n0_17116_17265  0.0218725 
iB33_78_v n1_16271_17312 0  0.0218725 
iB33_78_g 0 n0_17116_17298  0.0218725 
iB33_79_v n1_16271_17495 0  0.0218725 
iB33_79_g 0 n0_17116_17481  0.0218725 
iB33_80_v n1_16271_17528 0  0.0218725 
iB33_80_g 0 n0_17116_17535  0.0218725 
iB33_81_v n1_16271_17676 0  0.0218725 
iB33_81_g 0 n0_17116_17697  0.0218725 
iB33_82_v n1_16271_17684 0  0.0218725 
iB33_82_g 0 n0_17116_17697  0.0218725 
iB33_83_v n1_16271_17711 0  0.0218725 
iB33_83_g 0 n0_17116_17697  0.0218725 
iB33_84_v n1_16271_17744 0  0.0218725 
iB33_84_g 0 n0_17116_17730  0.0218725 
iB33_85_v n1_16271_17927 0  0.0218725 
iB33_85_g 0 n0_17116_17913  0.0218725 
iB33_86_v n1_16271_17960 0  0.0218725 
iB33_86_g 0 n0_17116_17946  0.0218725 
iB33_87_v n1_16271_18143 0  0.0218725 
iB33_87_g 0 n0_17116_18129  0.0218725 
iB33_88_v n1_16271_18176 0  0.0218725 
iB33_88_g 0 n0_17116_18176  0.0218725 
iB33_89_v n1_16271_18332 0  0.0218725 
iB33_89_g 0 n0_17116_18345  0.0218725 
iB33_90_v n1_16271_18359 0  0.0218725 
iB33_90_g 0 n0_17116_18345  0.0218725 
iB33_91_v n1_16271_18392 0  0.0218725 
iB33_91_g 0 n0_17116_18378  0.0218725 
iB33_92_v n1_16271_18527 0  0.0218725 
iB33_92_g 0 n0_17116_18561  0.0218725 
iB33_93_v n1_16271_18575 0  0.0218725 
iB33_93_g 0 n0_17116_18561  0.0218725 
iB33_94_v n1_16271_18608 0  0.0218725 
iB33_94_g 0 n0_17116_18594  0.0218725 
iB33_95_v n1_16364_18527 0  0.0218725 
iB33_95_g 0 n0_17116_18561  0.0218725 
iB33_96_v n1_16364_18575 0  0.0218725 
iB33_96_g 0 n0_17116_18561  0.0218725 
iB33_97_v n1_16364_18608 0  0.0218725 
iB33_97_g 0 n0_17116_18594  0.0218725 
iB33_98_v n1_16271_18764 0  0.0218725 
iB33_98_g 0 n0_17116_18777  0.0218725 
iB33_99_v n1_16271_18791 0  0.0218725 
iB33_99_g 0 n0_17116_18777  0.0218725 
iB33_100_v n1_16271_18824 0  0.0218725 
iB33_100_g 0 n0_17116_18810  0.0218725 
iB33_101_v n1_16271_19007 0  0.0218725 
iB33_101_g 0 n0_17116_18993  0.0218725 
iB33_102_v n1_16271_19040 0  0.0218725 
iB33_102_g 0 n0_17116_19040  0.0218725 
iB33_103_v n1_16364_18791 0  0.0218725 
iB33_103_g 0 n0_17116_18777  0.0218725 
iB33_104_v n1_16364_18824 0  0.0218725 
iB33_104_g 0 n0_17116_18810  0.0218725 
iB33_105_v n1_16364_19007 0  0.0218725 
iB33_105_g 0 n0_17116_18993  0.0218725 
iB33_106_v n1_16364_19040 0  0.0218725 
iB33_106_g 0 n0_17116_19040  0.0218725 
iB33_107_v n1_16271_19196 0  0.0218725 
iB33_107_g 0 n0_17116_19209  0.0218725 
iB33_108_v n1_16271_19223 0  0.0218725 
iB33_108_g 0 n0_17116_19209  0.0218725 
iB33_109_v n1_16271_19256 0  0.0218725 
iB33_109_g 0 n0_17116_19242  0.0218725 
iB33_110_v n1_16271_19412 0  0.0218725 
iB33_110_g 0 n0_17116_19425  0.0218725 
iB33_111_v n1_16271_19439 0  0.0218725 
iB33_111_g 0 n0_17116_19425  0.0218725 
iB33_112_v n1_16271_19472 0  0.0218725 
iB33_112_g 0 n0_17116_19458  0.0218725 
iB33_113_v n1_16364_19196 0  0.0218725 
iB33_113_g 0 n0_17116_19209  0.0218725 
iB33_114_v n1_16364_19223 0  0.0218725 
iB33_114_g 0 n0_17116_19209  0.0218725 
iB33_115_v n1_16364_19256 0  0.0218725 
iB33_115_g 0 n0_17116_19242  0.0218725 
iB33_116_v n1_16364_19439 0  0.0218725 
iB33_116_g 0 n0_17116_19425  0.0218725 
iB33_117_v n1_16364_19472 0  0.0218725 
iB33_117_g 0 n0_17116_19458  0.0218725 
iB33_118_v n1_16271_19655 0  0.0218725 
iB33_118_g 0 n0_17116_19641  0.0218725 
iB33_119_v n1_16271_19688 0  0.0218725 
iB33_119_g 0 n0_17116_19674  0.0218725 
iB33_120_v n1_16271_19871 0  0.0218725 
iB33_120_g 0 n0_17116_19857  0.0218725 
iB33_121_v n1_16271_19904 0  0.0218725 
iB33_121_g 0 n0_17116_19890  0.0218725 
iB33_122_v n1_16364_19655 0  0.0218725 
iB33_122_g 0 n0_17116_19641  0.0218725 
iB33_123_v n1_16364_19688 0  0.0218725 
iB33_123_g 0 n0_17116_19674  0.0218725 
iB33_124_v n1_16364_19871 0  0.0218725 
iB33_124_g 0 n0_17116_19857  0.0218725 
iB33_125_v n1_16364_19904 0  0.0218725 
iB33_125_g 0 n0_17116_19890  0.0218725 
iB33_126_v n1_16271_20087 0  0.0218725 
iB33_126_g 0 n0_17116_20073  0.0218725 
iB33_127_v n1_16271_20120 0  0.0218725 
iB33_127_g 0 n0_17116_20106  0.0218725 
iB33_128_v n1_16271_20303 0  0.0218725 
iB33_128_g 0 n0_17116_20289  0.0218725 
iB33_129_v n1_16271_20336 0  0.0218725 
iB33_129_g 0 n0_17116_20322  0.0218725 
iB33_130_v n1_16364_20087 0  0.0218725 
iB33_130_g 0 n0_17116_20073  0.0218725 
iB33_131_v n1_16364_20120 0  0.0218725 
iB33_131_g 0 n0_17116_20106  0.0218725 
iB33_132_v n1_16364_20303 0  0.0218725 
iB33_132_g 0 n0_17116_20289  0.0218725 
iB33_133_v n1_16364_20336 0  0.0218725 
iB33_133_g 0 n0_17116_20322  0.0218725 
iB33_134_v n1_16271_20519 0  0.0218725 
iB33_134_g 0 n0_17116_20505  0.0218725 
iB33_135_v n1_16271_20552 0  0.0218725 
iB33_135_g 0 n0_17116_20538  0.0218725 
iB33_136_v n1_16271_20687 0  0.0218725 
iB33_136_g 0 n0_17116_20754  0.0218725 
iB33_137_v n1_16271_20768 0  0.0218725 
iB33_137_g 0 n0_17116_20754  0.0218725 
iB33_138_v n1_16364_20519 0  0.0218725 
iB33_138_g 0 n0_17116_20505  0.0218725 
iB33_139_v n1_16364_20552 0  0.0218725 
iB33_139_g 0 n0_17116_20538  0.0218725 
iB33_140_v n1_16364_20687 0  0.0218725 
iB33_140_g 0 n0_17116_20754  0.0218725 
iB33_141_v n1_16364_20735 0  0.0218725 
iB33_141_g 0 n0_17116_20754  0.0218725 
iB33_142_v n1_16364_20768 0  0.0218725 
iB33_142_g 0 n0_17116_20754  0.0218725 
iB33_143_v n1_16271_20951 0  0.0218725 
iB33_143_g 0 n0_17116_20937  0.0218725 
iB33_144_v n1_16271_20984 0  0.0218725 
iB33_144_g 0 n0_17116_20970  0.0218725 
iB33_145_v n1_16364_20951 0  0.0218725 
iB33_145_g 0 n0_17116_20937  0.0218725 
iB33_146_v n1_16364_20984 0  0.0218725 
iB33_146_g 0 n0_17116_20970  0.0218725 
iB33_147_v n1_18150_18527 0  0.0218725 
iB33_147_g 0 n0_18241_18378  0.0218725 
iB33_148_v n1_18150_18575 0  0.0218725 
iB33_148_g 0 n0_18241_18378  0.0218725 
iB33_149_v n1_18150_18608 0  0.0218725 
iB33_149_g 0 n0_18241_18378  0.0218725 
iB33_150_v n1_18150_18791 0  0.0218725 
iB33_150_g 0 n0_18241_18378  0.0218725 
iB33_151_v n1_18150_18824 0  0.0218725 
iB33_151_g 0 n0_18241_18378  0.0218725 
iB33_152_v n1_18150_19007 0  0.0218725 
iB33_152_g 0 n0_18241_18378  0.0218725 
iB33_153_v n1_18150_19040 0  0.0218725 
iB33_153_g 0 n0_18241_18378  0.0218725 
iB33_154_v n1_18150_19223 0  0.0218725 
iB33_154_g 0 n0_17396_19209  0.0218725 
iB33_155_v n1_18150_19256 0  0.0218725 
iB33_155_g 0 n0_17396_19242  0.0218725 
iB33_156_v n1_18150_19439 0  0.0218725 
iB33_156_g 0 n0_17396_19425  0.0218725 
iB33_157_v n1_18150_19472 0  0.0218725 
iB33_157_g 0 n0_17396_19458  0.0218725 
iB33_158_v n1_18150_19655 0  0.0218725 
iB33_158_g 0 n0_17396_19641  0.0218725 
iB33_159_v n1_18150_19688 0  0.0218725 
iB33_159_g 0 n0_17396_19674  0.0218725 
iB33_160_v n1_18150_19871 0  0.0218725 
iB33_160_g 0 n0_17396_19857  0.0218725 
iB33_161_v n1_18150_19904 0  0.0218725 
iB33_161_g 0 n0_17396_19890  0.0218725 
iB33_162_v n1_18150_20087 0  0.0218725 
iB33_162_g 0 n0_17396_20073  0.0218725 
iB33_163_v n1_18150_20120 0  0.0218725 
iB33_163_g 0 n0_17396_20106  0.0218725 
iB33_164_v n1_18150_20303 0  0.0218725 
iB33_164_g 0 n0_17396_20289  0.0218725 
iB33_165_v n1_18150_20336 0  0.0218725 
iB33_165_g 0 n0_17396_20322  0.0218725 
iB33_166_v n1_18150_20519 0  0.0218725 
iB33_166_g 0 n0_17396_20505  0.0218725 
iB33_167_v n1_18150_20552 0  0.0218725 
iB33_167_g 0 n0_17396_20538  0.0218725 
iB33_168_v n1_18150_20687 0  0.0218725 
iB33_168_g 0 n0_17396_20754  0.0218725 
iB33_169_v n1_18150_20735 0  0.0218725 
iB33_169_g 0 n0_17396_20754  0.0218725 
iB33_170_v n1_18150_20768 0  0.0218725 
iB33_170_g 0 n0_17396_20754  0.0218725 
iB33_171_v n1_18150_20951 0  0.0218725 
iB33_171_g 0 n0_17396_20937  0.0218725 
iB33_172_v n1_18150_20984 0  0.0218725 
iB33_172_g 0 n0_17396_20970  0.0218725 
iB33_173_v n1_18333_15983 0  0.0218725 
iB33_173_g 0 n0_18241_15969  0.0218725 
iB33_174_v n1_18333_16016 0  0.0218725 
iB33_174_g 0 n0_18241_16002  0.0218725 
iB33_175_v n1_18333_16199 0  0.0218725 
iB33_175_g 0 n0_18241_16185  0.0218725 
iB33_176_v n1_18333_16232 0  0.0218725 
iB33_176_g 0 n0_18241_16218  0.0218725 
iB33_177_v n1_18380_16199 0  0.0218725 
iB33_177_g 0 n0_18241_16185  0.0218725 
iB33_178_v n1_18380_16232 0  0.0218725 
iB33_178_g 0 n0_18241_16218  0.0218725 
iB33_179_v n1_18521_15983 0  0.0218725 
iB33_179_g 0 n0_18429_15969  0.0218725 
iB33_180_v n1_18521_16016 0  0.0218725 
iB33_180_g 0 n0_18429_16002  0.0218725 
iB33_181_v n1_18521_16199 0  0.0218725 
iB33_181_g 0 n0_18429_16002  0.0218725 
iB33_182_v n1_18333_16415 0  0.0218725 
iB33_182_g 0 n0_18241_16401  0.0218725 
iB33_183_v n1_18333_16448 0  0.0218725 
iB33_183_g 0 n0_18241_16434  0.0218725 
iB33_184_v n1_18333_16631 0  0.0218725 
iB33_184_g 0 n0_18241_16617  0.0218725 
iB33_185_v n1_18333_16664 0  0.0218725 
iB33_185_g 0 n0_18241_16664  0.0218725 
iB33_186_v n1_18521_16415 0  0.0218725 
iB33_186_g 0 n0_18429_16401  0.0218725 
iB33_187_v n1_18521_16448 0  0.0218725 
iB33_187_g 0 n0_18429_16434  0.0218725 
iB33_188_v n1_18521_16631 0  0.0218725 
iB33_188_g 0 n0_18429_16617  0.0218725 
iB33_189_v n1_18521_16664 0  0.0218725 
iB33_189_g 0 n0_18429_16664  0.0218725 
iB33_190_v n1_18333_16812 0  0.0218725 
iB33_190_g 0 n0_18241_16833  0.0218725 
iB33_191_v n1_18333_16820 0  0.0218725 
iB33_191_g 0 n0_18241_16833  0.0218725 
iB33_192_v n1_18333_16847 0  0.0218725 
iB33_192_g 0 n0_18241_16833  0.0218725 
iB33_193_v n1_18333_16880 0  0.0218725 
iB33_193_g 0 n0_18241_16866  0.0218725 
iB33_194_v n1_18333_17063 0  0.0218725 
iB33_194_g 0 n0_18241_17049  0.0218725 
iB33_195_v n1_18333_17096 0  0.0218725 
iB33_195_g 0 n0_18241_17082  0.0218725 
iB33_196_v n1_18521_16812 0  0.0218725 
iB33_196_g 0 n0_18429_16833  0.0218725 
iB33_197_v n1_18521_16820 0  0.0218725 
iB33_197_g 0 n0_18429_16833  0.0218725 
iB33_198_v n1_18521_16847 0  0.0218725 
iB33_198_g 0 n0_18429_16833  0.0218725 
iB33_199_v n1_18521_16880 0  0.0218725 
iB33_199_g 0 n0_18429_16866  0.0218725 
iB33_200_v n1_18521_17063 0  0.0218725 
iB33_200_g 0 n0_18429_17049  0.0218725 
iB33_201_v n1_18521_17096 0  0.0218725 
iB33_201_g 0 n0_18429_17082  0.0218725 
iB33_202_v n1_18333_17230 0  0.0218725 
iB33_202_g 0 n0_18380_17298  0.0218725 
iB33_203_v n1_18333_17495 0  0.0218725 
iB33_203_g 0 n0_18241_17481  0.0218725 
iB33_204_v n1_18521_17230 0  0.0218725 
iB33_204_g 0 n0_18429_17265  0.0218725 
iB33_205_v n1_18521_17279 0  0.0218725 
iB33_205_g 0 n0_18429_17265  0.0218725 
iB33_206_v n1_18521_17312 0  0.0218725 
iB33_206_g 0 n0_18429_17298  0.0218725 
iB33_207_v n1_18521_17495 0  0.0218725 
iB33_207_g 0 n0_18429_17481  0.0218725 
iB33_208_v n1_18333_17528 0  0.0218725 
iB33_208_g 0 n0_18241_17514  0.0218725 
iB33_209_v n1_18333_17711 0  0.0218725 
iB33_209_g 0 n0_18241_17697  0.0218725 
iB33_210_v n1_18333_17744 0  0.0218725 
iB33_210_g 0 n0_18241_17744  0.0218725 
iB33_211_v n1_18333_17900 0  0.0218725 
iB33_211_g 0 n0_18241_17913  0.0218725 
iB33_212_v n1_18333_17927 0  0.0218725 
iB33_212_g 0 n0_18241_17913  0.0218725 
iB33_213_v n1_18521_17528 0  0.0218725 
iB33_213_g 0 n0_18429_17514  0.0218725 
iB33_214_v n1_18521_17711 0  0.0218725 
iB33_214_g 0 n0_18429_17697  0.0218725 
iB33_215_v n1_18521_17744 0  0.0218725 
iB33_215_g 0 n0_18429_17744  0.0218725 
iB33_216_v n1_18521_17900 0  0.0218725 
iB33_216_g 0 n0_18429_17913  0.0218725 
iB33_217_v n1_18521_17927 0  0.0218725 
iB33_217_g 0 n0_18429_17913  0.0218725 
iB33_218_v n1_18333_17960 0  0.0218725 
iB33_218_g 0 n0_18241_17946  0.0218725 
iB33_219_v n1_18333_18143 0  0.0218725 
iB33_219_g 0 n0_18241_18129  0.0218725 
iB33_220_v n1_18333_18176 0  0.0218725 
iB33_220_g 0 n0_18241_18162  0.0218725 
iB33_221_v n1_18521_17960 0  0.0218725 
iB33_221_g 0 n0_18429_17946  0.0218725 
iB33_222_v n1_18521_18143 0  0.0218725 
iB33_222_g 0 n0_18429_18129  0.0218725 
iB33_223_v n1_18521_18176 0  0.0218725 
iB33_223_g 0 n0_18429_18162  0.0218725 
iB33_224_v n1_18333_18359 0  0.0218725 
iB33_224_g 0 n0_18241_18345  0.0218725 
iB33_225_v n1_18333_18392 0  0.0218725 
iB33_225_g 0 n0_18241_18378  0.0218725 
iB33_226_v n1_18333_18527 0  0.0218725 
iB33_226_g 0 n0_18241_18378  0.0218725 
iB33_227_v n1_18333_18575 0  0.0218725 
iB33_227_g 0 n0_18241_18378  0.0218725 
iB33_228_v n1_18333_18608 0  0.0218725 
iB33_228_g 0 n0_18241_18378  0.0218725 
iB33_229_v n1_18380_18392 0  0.0218725 
iB33_229_g 0 n0_18429_18345  0.0218725 
iB33_230_v n1_18380_18527 0  0.0218725 
iB33_230_g 0 n0_18429_18345  0.0218725 
iB33_231_v n1_18521_18359 0  0.0218725 
iB33_231_g 0 n0_18429_18345  0.0218725 
iB33_232_v n1_18521_18392 0  0.0218725 
iB33_232_g 0 n0_18429_18345  0.0218725 
iB33_233_v n1_18521_18527 0  0.0218725 
iB33_233_g 0 n0_18429_18345  0.0218725 
iB33_234_v n1_18521_18575 0  0.0218725 
iB33_234_g 0 n0_18429_18345  0.0218725 
iB33_235_v n1_18521_18608 0  0.0218725 
iB33_235_g 0 n0_18429_18345  0.0218725 
iB33_236_v n1_18333_18791 0  0.0218725 
iB33_236_g 0 n0_18241_18378  0.0218725 
iB33_237_v n1_18333_18824 0  0.0218725 
iB33_237_g 0 n0_18241_18378  0.0218725 
iB33_238_v n1_18333_19007 0  0.0218725 
iB33_238_g 0 n0_18241_18378  0.0218725 
iB33_239_v n1_18333_19040 0  0.0218725 
iB33_239_g 0 n0_18241_18378  0.0218725 
iB33_240_v n1_18521_18791 0  0.0218725 
iB33_240_g 0 n0_18429_18345  0.0218725 
iB33_241_v n1_18521_18824 0  0.0218725 
iB33_241_g 0 n0_18429_18345  0.0218725 
iB33_242_v n1_18521_19007 0  0.0218725 
iB33_242_g 0 n0_18429_18345  0.0218725 
iB33_243_v n1_18521_19040 0  0.0218725 
iB33_243_g 0 n0_18429_18345  0.0218725 
iB33_244_v n1_18333_19223 0  0.0218725 
iB33_244_g 0 n0_18241_18378  0.0218725 
iB33_245_v n1_18333_19256 0  0.0218725 
iB33_245_g 0 n0_17396_19242  0.0218725 
iB33_246_v n1_18333_19439 0  0.0218725 
iB33_246_g 0 n0_17396_19425  0.0218725 
iB33_247_v n1_18333_19472 0  0.0218725 
iB33_247_g 0 n0_17396_19458  0.0218725 
iB33_248_v n1_18521_19223 0  0.0218725 
iB33_248_g 0 n0_19366_19209  0.0218725 
iB33_249_v n1_18521_19256 0  0.0218725 
iB33_249_g 0 n0_19366_19242  0.0218725 
iB33_250_v n1_18521_19439 0  0.0218725 
iB33_250_g 0 n0_19366_19425  0.0218725 
iB33_251_v n1_18521_19472 0  0.0218725 
iB33_251_g 0 n0_19366_19458  0.0218725 
iB33_252_v n1_18333_19871 0  0.0218725 
iB33_252_g 0 n0_17396_19857  0.0218725 
iB33_253_v n1_18333_19904 0  0.0218725 
iB33_253_g 0 n0_17396_19890  0.0218725 
iB33_254_v n1_18521_19655 0  0.0218725 
iB33_254_g 0 n0_19366_19641  0.0218725 
iB33_255_v n1_18521_19688 0  0.0218725 
iB33_255_g 0 n0_19366_19674  0.0218725 
iB33_256_v n1_18521_19871 0  0.0218725 
iB33_256_g 0 n0_19366_19857  0.0218725 
iB33_257_v n1_18521_19904 0  0.0218725 
iB33_257_g 0 n0_19366_19890  0.0218725 
iB33_258_v n1_18333_20087 0  0.0218725 
iB33_258_g 0 n0_17396_20073  0.0218725 
iB33_259_v n1_18333_20120 0  0.0218725 
iB33_259_g 0 n0_17396_20106  0.0218725 
iB33_260_v n1_18333_20303 0  0.0218725 
iB33_260_g 0 n0_17396_20289  0.0218725 
iB33_261_v n1_18333_20336 0  0.0218725 
iB33_261_g 0 n0_17396_20322  0.0218725 
iB33_262_v n1_18521_20087 0  0.0218725 
iB33_262_g 0 n0_19366_20073  0.0218725 
iB33_263_v n1_18521_20120 0  0.0218725 
iB33_263_g 0 n0_19366_20106  0.0218725 
iB33_264_v n1_18521_20303 0  0.0218725 
iB33_264_g 0 n0_19366_20289  0.0218725 
iB33_265_v n1_18521_20336 0  0.0218725 
iB33_265_g 0 n0_19366_20322  0.0218725 
iB33_266_v n1_18333_20519 0  0.0218725 
iB33_266_g 0 n0_17396_20505  0.0218725 
iB33_267_v n1_18333_20552 0  0.0218725 
iB33_267_g 0 n0_17396_20538  0.0218725 
iB33_268_v n1_18333_20687 0  0.0218725 
iB33_268_g 0 n0_17396_20754  0.0218725 
iB33_269_v n1_18333_20735 0  0.0218725 
iB33_269_g 0 n0_17396_20754  0.0218725 
iB33_270_v n1_18333_20768 0  0.0218725 
iB33_270_g 0 n0_17396_20754  0.0218725 
iB33_271_v n1_18380_20687 0  0.0218725 
iB33_271_g 0 n0_17396_20754  0.0218725 
iB33_272_v n1_18380_20735 0  0.0218725 
iB33_272_g 0 n0_17396_20754  0.0218725 
iB33_273_v n1_18380_20768 0  0.0218725 
iB33_273_g 0 n0_17396_20754  0.0218725 
iB33_274_v n1_18521_20519 0  0.0218725 
iB33_274_g 0 n0_19366_20505  0.0218725 
iB33_275_v n1_18521_20552 0  0.0218725 
iB33_275_g 0 n0_19366_20538  0.0218725 
iB33_276_v n1_18521_20687 0  0.0218725 
iB33_276_g 0 n0_19366_20754  0.0218725 
iB33_277_v n1_18521_20768 0  0.0218725 
iB33_277_g 0 n0_19366_20754  0.0218725 
iB33_278_v n1_18333_20951 0  0.0218725 
iB33_278_g 0 n0_17396_20937  0.0218725 
iB33_279_v n1_18333_20984 0  0.0218725 
iB33_279_g 0 n0_17396_20970  0.0218725 
iB33_280_v n1_18521_20951 0  0.0218725 
iB33_280_g 0 n0_19366_20937  0.0218725 
iB33_281_v n1_18521_20984 0  0.0218725 
iB33_281_g 0 n0_19366_20970  0.0218725 
iB33_282_v n1_18614_18527 0  0.0218725 
iB33_282_g 0 n0_18429_18345  0.0218725 
iB33_283_v n1_18614_18575 0  0.0218725 
iB33_283_g 0 n0_18429_18345  0.0218725 
iB33_284_v n1_18614_18608 0  0.0218725 
iB33_284_g 0 n0_18429_18345  0.0218725 
iB33_285_v n1_18614_18791 0  0.0218725 
iB33_285_g 0 n0_18429_18345  0.0218725 
iB33_286_v n1_18614_18824 0  0.0218725 
iB33_286_g 0 n0_18429_18345  0.0218725 
iB33_287_v n1_18614_19007 0  0.0218725 
iB33_287_g 0 n0_18429_18345  0.0218725 
iB33_288_v n1_18614_19040 0  0.0218725 
iB33_288_g 0 n0_18429_18345  0.0218725 
iB33_289_v n1_18614_19223 0  0.0218725 
iB33_289_g 0 n0_19366_19209  0.0218725 
iB33_290_v n1_18614_19256 0  0.0218725 
iB33_290_g 0 n0_19366_19242  0.0218725 
iB33_291_v n1_18614_19439 0  0.0218725 
iB33_291_g 0 n0_19366_19425  0.0218725 
iB33_292_v n1_18614_19472 0  0.0218725 
iB33_292_g 0 n0_19366_19458  0.0218725 
iB33_293_v n1_18614_19655 0  0.0218725 
iB33_293_g 0 n0_19366_19641  0.0218725 
iB33_294_v n1_18614_19688 0  0.0218725 
iB33_294_g 0 n0_19366_19674  0.0218725 
iB33_295_v n1_18614_19871 0  0.0218725 
iB33_295_g 0 n0_19366_19857  0.0218725 
iB33_296_v n1_18614_19904 0  0.0218725 
iB33_296_g 0 n0_19366_19890  0.0218725 
iB33_297_v n1_18614_20087 0  0.0218725 
iB33_297_g 0 n0_19366_20073  0.0218725 
iB33_298_v n1_18614_20120 0  0.0218725 
iB33_298_g 0 n0_19366_20106  0.0218725 
iB33_299_v n1_18614_20303 0  0.0218725 
iB33_299_g 0 n0_19366_20289  0.0218725 
iB33_300_v n1_18614_20336 0  0.0218725 
iB33_300_g 0 n0_19366_20322  0.0218725 
iB33_301_v n1_18614_20519 0  0.0218725 
iB33_301_g 0 n0_19366_20505  0.0218725 
iB33_302_v n1_18614_20552 0  0.0218725 
iB33_302_g 0 n0_19366_20538  0.0218725 
iB33_303_v n1_18614_20687 0  0.0218725 
iB33_303_g 0 n0_19366_20754  0.0218725 
iB33_304_v n1_18614_20735 0  0.0218725 
iB33_304_g 0 n0_19366_20754  0.0218725 
iB33_305_v n1_18614_20768 0  0.0218725 
iB33_305_g 0 n0_19366_20754  0.0218725 
iB33_306_v n1_18614_20951 0  0.0218725 
iB33_306_g 0 n0_19366_20937  0.0218725 
iB33_307_v n1_18614_20984 0  0.0218725 
iB33_307_g 0 n0_19366_20970  0.0218725 
iB33_308_v n1_20583_15983 0  0.0218725 
iB33_308_g 0 n0_20491_15969  0.0218725 
iB33_309_v n1_20583_16016 0  0.0218725 
iB33_309_g 0 n0_20491_16002  0.0218725 
iB33_310_v n1_20583_16199 0  0.0218725 
iB33_310_g 0 n0_20491_16185  0.0218725 
iB33_311_v n1_20583_16232 0  0.0218725 
iB33_311_g 0 n0_20491_16218  0.0218725 
iB33_312_v n1_20630_16199 0  0.0218725 
iB33_312_g 0 n0_20491_16185  0.0218725 
iB33_313_v n1_20630_16232 0  0.0218725 
iB33_313_g 0 n0_20491_16218  0.0218725 
iB33_314_v n1_20771_15983 0  0.0218725 
iB33_314_g 0 n0_20679_15969  0.0218725 
iB33_315_v n1_20771_16016 0  0.0218725 
iB33_315_g 0 n0_20679_16002  0.0218725 
iB33_316_v n1_20771_16199 0  0.0218725 
iB33_316_g 0 n0_20679_16002  0.0218725 
iB33_317_v n1_20583_16415 0  0.0218725 
iB33_317_g 0 n0_20491_16401  0.0218725 
iB33_318_v n1_20583_16448 0  0.0218725 
iB33_318_g 0 n0_20491_16434  0.0218725 
iB33_319_v n1_20583_16631 0  0.0218725 
iB33_319_g 0 n0_20491_16617  0.0218725 
iB33_320_v n1_20583_16664 0  0.0218725 
iB33_320_g 0 n0_20491_16650  0.0218725 
iB33_321_v n1_20771_16415 0  0.0218725 
iB33_321_g 0 n0_20679_16401  0.0218725 
iB33_322_v n1_20771_16448 0  0.0218725 
iB33_322_g 0 n0_20679_16434  0.0218725 
iB33_323_v n1_20771_16631 0  0.0218725 
iB33_323_g 0 n0_20679_16617  0.0218725 
iB33_324_v n1_20771_16664 0  0.0218725 
iB33_324_g 0 n0_20679_16650  0.0218725 
iB33_325_v n1_20583_16798 0  0.0218725 
iB33_325_g 0 n0_20491_16833  0.0218725 
iB33_326_v n1_20583_16847 0  0.0218725 
iB33_326_g 0 n0_20491_16833  0.0218725 
iB33_327_v n1_20583_16880 0  0.0218725 
iB33_327_g 0 n0_20491_16866  0.0218725 
iB33_328_v n1_20583_17063 0  0.0218725 
iB33_328_g 0 n0_20491_17049  0.0218725 
iB33_329_v n1_20583_17096 0  0.0218725 
iB33_329_g 0 n0_20491_17082  0.0218725 
iB33_330_v n1_20771_16798 0  0.0218725 
iB33_330_g 0 n0_20679_16833  0.0218725 
iB33_331_v n1_20771_16847 0  0.0218725 
iB33_331_g 0 n0_20679_16833  0.0218725 
iB33_332_v n1_20771_16880 0  0.0218725 
iB33_332_g 0 n0_20679_16866  0.0218725 
iB33_333_v n1_20771_17063 0  0.0218725 
iB33_333_g 0 n0_20679_17049  0.0218725 
iB33_334_v n1_20771_17096 0  0.0218725 
iB33_334_g 0 n0_20679_17082  0.0218725 
iB33_335_v n1_20583_17495 0  0.0218725 
iB33_335_g 0 n0_20491_17481  0.0218725 
iB33_336_v n1_20771_17279 0  0.0218725 
iB33_336_g 0 n0_20679_17265  0.0218725 
iB33_337_v n1_20771_17312 0  0.0218725 
iB33_337_g 0 n0_20679_17298  0.0218725 
iB33_338_v n1_20771_17495 0  0.0218725 
iB33_338_g 0 n0_20679_17481  0.0218725 
iB33_339_v n1_20583_17528 0  0.0218725 
iB33_339_g 0 n0_20491_17514  0.0218725 
iB33_340_v n1_20583_17711 0  0.0218725 
iB33_340_g 0 n0_20491_17697  0.0218725 
iB33_341_v n1_20583_17744 0  0.0218725 
iB33_341_g 0 n0_20491_17730  0.0218725 
iB33_342_v n1_20583_17927 0  0.0218725 
iB33_342_g 0 n0_20491_17913  0.0218725 
iB33_343_v n1_20771_17528 0  0.0218725 
iB33_343_g 0 n0_20679_17514  0.0218725 
iB33_344_v n1_20771_17711 0  0.0218725 
iB33_344_g 0 n0_20679_17697  0.0218725 
iB33_345_v n1_20771_17744 0  0.0218725 
iB33_345_g 0 n0_20679_17730  0.0218725 
iB33_346_v n1_20771_17927 0  0.0218725 
iB33_346_g 0 n0_20679_17913  0.0218725 
iB33_347_v n1_20583_17960 0  0.0218725 
iB33_347_g 0 n0_20491_17946  0.0218725 
iB33_348_v n1_20583_18143 0  0.0218725 
iB33_348_g 0 n0_20491_18129  0.0218725 
iB33_349_v n1_20583_18176 0  0.0218725 
iB33_349_g 0 n0_20491_18162  0.0218725 
iB33_350_v n1_20771_17960 0  0.0218725 
iB33_350_g 0 n0_20679_17946  0.0218725 
iB33_351_v n1_20771_18143 0  0.0218725 
iB33_351_g 0 n0_20679_18129  0.0218725 
iB33_352_v n1_20771_18176 0  0.0218725 
iB33_352_g 0 n0_20679_18162  0.0218725 
iB33_353_v n1_20583_18359 0  0.0218725 
iB33_353_g 0 n0_20491_18345  0.0218725 
iB33_354_v n1_20583_18392 0  0.0218725 
iB33_354_g 0 n0_20491_18378  0.0218725 
iB33_355_v n1_20583_18527 0  0.0218725 
iB33_355_g 0 n0_20491_18561  0.0218725 
iB33_356_v n1_20583_18575 0  0.0218725 
iB33_356_g 0 n0_20491_18561  0.0218725 
iB33_357_v n1_20583_18608 0  0.0218725 
iB33_357_g 0 n0_20491_18594  0.0218725 
iB33_358_v n1_20630_18392 0  0.0218725 
iB33_358_g 0 n0_20679_18345  0.0218725 
iB33_359_v n1_20630_18527 0  0.0218725 
iB33_359_g 0 n0_20679_18594  0.0218725 
iB33_360_v n1_20771_18359 0  0.0218725 
iB33_360_g 0 n0_20679_18345  0.0218725 
iB33_361_v n1_20771_18392 0  0.0218725 
iB33_361_g 0 n0_20679_18345  0.0218725 
iB33_362_v n1_20771_18527 0  0.0218725 
iB33_362_g 0 n0_20679_18594  0.0218725 
iB33_363_v n1_20771_18575 0  0.0218725 
iB33_363_g 0 n0_20679_18594  0.0218725 
iB33_364_v n1_20771_18608 0  0.0218725 
iB33_364_g 0 n0_20679_18594  0.0218725 
iB33_365_v n1_20583_18791 0  0.0218725 
iB33_365_g 0 n0_20491_18777  0.0218725 
iB33_366_v n1_20583_18824 0  0.0218725 
iB33_366_g 0 n0_20491_18810  0.0218725 
iB33_367_v n1_20583_19007 0  0.0218725 
iB33_367_g 0 n0_20491_18993  0.0218725 
iB33_368_v n1_20583_19040 0  0.0218725 
iB33_368_g 0 n0_20491_19040  0.0218725 
iB33_369_v n1_20771_18791 0  0.0218725 
iB33_369_g 0 n0_20679_18777  0.0218725 
iB33_370_v n1_20771_18824 0  0.0218725 
iB33_370_g 0 n0_20679_18810  0.0218725 
iB33_371_v n1_20771_19007 0  0.0218725 
iB33_371_g 0 n0_20679_18993  0.0218725 
iB33_372_v n1_20771_19040 0  0.0218725 
iB33_372_g 0 n0_20679_19040  0.0218725 
iB33_373_v n1_20583_19223 0  0.0218725 
iB33_373_g 0 n0_20491_19209  0.0218725 
iB33_374_v n1_20583_19256 0  0.0218725 
iB33_374_g 0 n0_20491_19242  0.0218725 
iB33_375_v n1_20583_19439 0  0.0218725 
iB33_375_g 0 n0_20491_19425  0.0218725 
iB33_376_v n1_20583_19472 0  0.0218725 
iB33_376_g 0 n0_20491_19458  0.0218725 
iB33_377_v n1_20771_19223 0  0.0218725 
iB33_377_g 0 n0_20679_19209  0.0218725 
iB33_378_v n1_20771_19256 0  0.0218725 
iB33_378_g 0 n0_20679_19242  0.0218725 
iB33_379_v n1_20771_19439 0  0.0218725 
iB33_379_g 0 n0_20679_19425  0.0218725 
iB33_380_v n1_20771_19472 0  0.0218725 
iB33_380_g 0 n0_20679_19458  0.0218725 
iB33_381_v n1_20583_19871 0  0.0218725 
iB33_381_g 0 n0_20491_19857  0.0218725 
iB33_382_v n1_20583_19904 0  0.0218725 
iB33_382_g 0 n0_20491_19890  0.0218725 
iB33_383_v n1_20771_19655 0  0.0218725 
iB33_383_g 0 n0_20679_19641  0.0218725 
iB33_384_v n1_20771_19688 0  0.0218725 
iB33_384_g 0 n0_20679_19674  0.0218725 
iB33_385_v n1_20771_19871 0  0.0218725 
iB33_385_g 0 n0_20679_19857  0.0218725 
iB33_386_v n1_20771_19904 0  0.0218725 
iB33_386_g 0 n0_20679_19890  0.0218725 
iB33_387_v n1_20583_20087 0  0.0218725 
iB33_387_g 0 n0_20491_20073  0.0218725 
iB33_388_v n1_20583_20120 0  0.0218725 
iB33_388_g 0 n0_20491_20106  0.0218725 
iB33_389_v n1_20583_20303 0  0.0218725 
iB33_389_g 0 n0_20491_20289  0.0218725 
iB33_390_v n1_20583_20336 0  0.0218725 
iB33_390_g 0 n0_20491_20322  0.0218725 
iB33_391_v n1_20771_20087 0  0.0218725 
iB33_391_g 0 n0_20679_20073  0.0218725 
iB33_392_v n1_20771_20120 0  0.0218725 
iB33_392_g 0 n0_20679_20106  0.0218725 
iB33_393_v n1_20771_20303 0  0.0218725 
iB33_393_g 0 n0_20679_20289  0.0218725 
iB33_394_v n1_20771_20336 0  0.0218725 
iB33_394_g 0 n0_20679_20322  0.0218725 
iB33_395_v n1_20583_20519 0  0.0218725 
iB33_395_g 0 n0_20491_20505  0.0218725 
iB33_396_v n1_20583_20552 0  0.0218725 
iB33_396_g 0 n0_20491_20538  0.0218725 
iB33_397_v n1_20583_20687 0  0.0218725 
iB33_397_g 0 n0_20491_20538  0.0218725 
iB33_398_v n1_20583_20735 0  0.0218725 
iB33_398_g 0 n0_20491_20538  0.0218725 
iB33_399_v n1_20583_20768 0  0.0218725 
iB33_399_g 0 n0_20491_20538  0.0218725 
iB33_400_v n1_20630_20687 0  0.0218725 
iB33_400_g 0 n0_20679_20538  0.0218725 
iB33_401_v n1_20630_20735 0  0.0218725 
iB33_401_g 0 n0_20679_20538  0.0218725 
iB33_402_v n1_20630_20768 0  0.0218725 
iB33_402_g 0 n0_20679_20538  0.0218725 
iB33_403_v n1_20771_20519 0  0.0218725 
iB33_403_g 0 n0_20679_20505  0.0218725 
iB33_404_v n1_20771_20552 0  0.0218725 
iB33_404_g 0 n0_20679_20538  0.0218725 
iB33_405_v n1_20771_20687 0  0.0218725 
iB33_405_g 0 n0_20679_20538  0.0218725 
iB33_406_v n1_20583_20951 0  0.0218725 
iB33_406_g 0 n0_20491_20538  0.0218725 
iB33_407_v n1_20583_20984 0  0.0218725 
iB33_407_g 0 n0_20491_20538  0.0218725 
iB00_0_v n1_333_383 0  0.0174842 
iB00_0_g 0 n0_241_633  0.0174842 
iB00_1_v n1_521_215 0  0.0174842 
iB00_1_g 0 n0_429_633  0.0174842 
iB00_2_v n1_521_248 0  0.0174842 
iB00_2_g 0 n0_429_633  0.0174842 
iB00_3_v n1_521_383 0  0.0174842 
iB00_3_g 0 n0_429_633  0.0174842 
iB00_4_v n1_333_431 0  0.0174842 
iB00_4_g 0 n0_241_633  0.0174842 
iB00_5_v n1_333_464 0  0.0174842 
iB00_5_g 0 n0_241_633  0.0174842 
iB00_6_v n1_333_647 0  0.0174842 
iB00_6_g 0 n0_241_633  0.0174842 
iB00_7_v n1_333_680 0  0.0174842 
iB00_7_g 0 n0_241_666  0.0174842 
iB00_8_v n1_380_431 0  0.0174842 
iB00_8_g 0 n0_429_633  0.0174842 
iB00_9_v n1_380_464 0  0.0174842 
iB00_9_g 0 n0_429_633  0.0174842 
iB00_10_v n1_521_431 0  0.0174842 
iB00_10_g 0 n0_429_633  0.0174842 
iB00_11_v n1_521_647 0  0.0174842 
iB00_11_g 0 n0_429_633  0.0174842 
iB00_12_v n1_521_680 0  0.0174842 
iB00_12_g 0 n0_429_666  0.0174842 
iB00_13_v n1_333_863 0  0.0174842 
iB00_13_g 0 n0_241_849  0.0174842 
iB00_14_v n1_333_896 0  0.0174842 
iB00_14_g 0 n0_241_882  0.0174842 
iB00_15_v n1_333_1079 0  0.0174842 
iB00_15_g 0 n0_241_1065  0.0174842 
iB00_16_v n1_333_1112 0  0.0174842 
iB00_16_g 0 n0_241_1098  0.0174842 
iB00_17_v n1_521_863 0  0.0174842 
iB00_17_g 0 n0_429_849  0.0174842 
iB00_18_v n1_521_896 0  0.0174842 
iB00_18_g 0 n0_429_882  0.0174842 
iB00_19_v n1_521_1079 0  0.0174842 
iB00_19_g 0 n0_429_1065  0.0174842 
iB00_20_v n1_521_1112 0  0.0174842 
iB00_20_g 0 n0_429_1098  0.0174842 
iB00_21_v n1_333_1295 0  0.0174842 
iB00_21_g 0 n0_241_1281  0.0174842 
iB00_22_v n1_333_1328 0  0.0174842 
iB00_22_g 0 n0_241_1314  0.0174842 
iB00_23_v n1_521_1295 0  0.0174842 
iB00_23_g 0 n0_429_1281  0.0174842 
iB00_24_v n1_521_1328 0  0.0174842 
iB00_24_g 0 n0_429_1314  0.0174842 
iB00_25_v n1_521_1511 0  0.0174842 
iB00_25_g 0 n0_429_1497  0.0174842 
iB00_26_v n1_521_1544 0  0.0174842 
iB00_26_g 0 n0_429_1530  0.0174842 
iB00_27_v n1_333_1727 0  0.0174842 
iB00_27_g 0 n0_241_1713  0.0174842 
iB00_28_v n1_333_1760 0  0.0174842 
iB00_28_g 0 n0_241_1746  0.0174842 
iB00_29_v n1_333_1943 0  0.0174842 
iB00_29_g 0 n0_241_1929  0.0174842 
iB00_30_v n1_333_1976 0  0.0174842 
iB00_30_g 0 n0_241_1962  0.0174842 
iB00_31_v n1_521_1727 0  0.0174842 
iB00_31_g 0 n0_429_1713  0.0174842 
iB00_32_v n1_521_1760 0  0.0174842 
iB00_32_g 0 n0_429_1746  0.0174842 
iB00_33_v n1_521_1943 0  0.0174842 
iB00_33_g 0 n0_429_1929  0.0174842 
iB00_34_v n1_521_1976 0  0.0174842 
iB00_34_g 0 n0_429_1962  0.0174842 
iB00_35_v n1_333_2159 0  0.0174842 
iB00_35_g 0 n0_241_2145  0.0174842 
iB00_36_v n1_333_2192 0  0.0174842 
iB00_36_g 0 n0_241_2178  0.0174842 
iB00_37_v n1_333_2375 0  0.0174842 
iB00_37_g 0 n0_241_2361  0.0174842 
iB00_38_v n1_333_2408 0  0.0174842 
iB00_38_g 0 n0_241_2394  0.0174842 
iB00_39_v n1_521_2159 0  0.0174842 
iB00_39_g 0 n0_429_2145  0.0174842 
iB00_40_v n1_521_2192 0  0.0174842 
iB00_40_g 0 n0_429_2178  0.0174842 
iB00_41_v n1_521_2375 0  0.0174842 
iB00_41_g 0 n0_429_2361  0.0174842 
iB00_42_v n1_521_2408 0  0.0174842 
iB00_42_g 0 n0_429_2394  0.0174842 
iB00_43_v n1_333_2543 0  0.0174842 
iB00_43_g 0 n0_241_2577  0.0174842 
iB00_44_v n1_333_2591 0  0.0174842 
iB00_44_g 0 n0_241_2577  0.0174842 
iB00_45_v n1_333_2624 0  0.0174842 
iB00_45_g 0 n0_241_2610  0.0174842 
iB00_46_v n1_333_2807 0  0.0174842 
iB00_46_g 0 n0_241_2793  0.0174842 
iB00_47_v n1_333_2840 0  0.0174842 
iB00_47_g 0 n0_241_2826  0.0174842 
iB00_48_v n1_521_2543 0  0.0174842 
iB00_48_g 0 n0_429_2577  0.0174842 
iB00_49_v n1_521_2591 0  0.0174842 
iB00_49_g 0 n0_429_2577  0.0174842 
iB00_50_v n1_521_2624 0  0.0174842 
iB00_50_g 0 n0_429_2610  0.0174842 
iB00_51_v n1_521_2807 0  0.0174842 
iB00_51_g 0 n0_429_2826  0.0174842 
iB00_52_v n1_521_2840 0  0.0174842 
iB00_52_g 0 n0_429_2826  0.0174842 
iB00_53_v n1_333_3023 0  0.0174842 
iB00_53_g 0 n0_241_3009  0.0174842 
iB00_54_v n1_333_3056 0  0.0174842 
iB00_54_g 0 n0_241_3042  0.0174842 
iB00_55_v n1_333_3239 0  0.0174842 
iB00_55_g 0 n0_241_3225  0.0174842 
iB00_56_v n1_521_3023 0  0.0174842 
iB00_56_g 0 n0_429_3009  0.0174842 
iB00_57_v n1_521_3056 0  0.0174842 
iB00_57_g 0 n0_429_3042  0.0174842 
iB00_58_v n1_521_3239 0  0.0174842 
iB00_58_g 0 n0_429_3225  0.0174842 
iB00_59_v n1_333_3272 0  0.0174842 
iB00_59_g 0 n0_241_3258  0.0174842 
iB00_60_v n1_333_3455 0  0.0174842 
iB00_60_g 0 n0_241_3441  0.0174842 
iB00_61_v n1_333_3488 0  0.0174842 
iB00_61_g 0 n0_241_3474  0.0174842 
iB00_62_v n1_333_3671 0  0.0174842 
iB00_62_g 0 n0_241_3657  0.0174842 
iB00_63_v n1_521_3272 0  0.0174842 
iB00_63_g 0 n0_429_3258  0.0174842 
iB00_64_v n1_521_3455 0  0.0174842 
iB00_64_g 0 n0_429_3441  0.0174842 
iB00_65_v n1_521_3488 0  0.0174842 
iB00_65_g 0 n0_429_3474  0.0174842 
iB00_66_v n1_521_3671 0  0.0174842 
iB00_66_g 0 n0_429_3657  0.0174842 
iB00_67_v n1_333_3704 0  0.0174842 
iB00_67_g 0 n0_241_3690  0.0174842 
iB00_68_v n1_521_3704 0  0.0174842 
iB00_68_g 0 n0_429_3690  0.0174842 
iB00_69_v n1_521_3887 0  0.0174842 
iB00_69_g 0 n0_429_3873  0.0174842 
iB00_70_v n1_521_3920 0  0.0174842 
iB00_70_g 0 n0_429_3906  0.0174842 
iB00_71_v n1_333_4103 0  0.0174842 
iB00_71_g 0 n0_241_4089  0.0174842 
iB00_72_v n1_333_4136 0  0.0174842 
iB00_72_g 0 n0_241_4122  0.0174842 
iB00_73_v n1_333_4319 0  0.0174842 
iB00_73_g 0 n0_241_4305  0.0174842 
iB00_74_v n1_333_4352 0  0.0174842 
iB00_74_g 0 n0_241_4338  0.0174842 
iB00_75_v n1_333_4486 0  0.0174842 
iB00_75_g 0 n0_241_4521  0.0174842 
iB00_76_v n1_521_4103 0  0.0174842 
iB00_76_g 0 n0_429_4089  0.0174842 
iB00_77_v n1_521_4136 0  0.0174842 
iB00_77_g 0 n0_429_4122  0.0174842 
iB00_78_v n1_521_4319 0  0.0174842 
iB00_78_g 0 n0_429_4305  0.0174842 
iB00_79_v n1_521_4352 0  0.0174842 
iB00_79_g 0 n0_429_4338  0.0174842 
iB00_80_v n1_521_4486 0  0.0174842 
iB00_80_g 0 n0_429_4521  0.0174842 
iB00_81_v n1_333_4535 0  0.0174842 
iB00_81_g 0 n0_241_4521  0.0174842 
iB00_82_v n1_333_4568 0  0.0174842 
iB00_82_g 0 n0_241_4554  0.0174842 
iB00_83_v n1_333_4751 0  0.0174842 
iB00_83_g 0 n0_241_4737  0.0174842 
iB00_84_v n1_333_4784 0  0.0174842 
iB00_84_g 0 n0_241_4770  0.0174842 
iB00_85_v n1_521_4535 0  0.0174842 
iB00_85_g 0 n0_429_4521  0.0174842 
iB00_86_v n1_521_4568 0  0.0174842 
iB00_86_g 0 n0_429_4554  0.0174842 
iB00_87_v n1_521_4751 0  0.0174842 
iB00_87_g 0 n0_429_4737  0.0174842 
iB00_88_v n1_521_4784 0  0.0174842 
iB00_88_g 0 n0_429_4770  0.0174842 
iB00_89_v n1_333_4967 0  0.0174842 
iB00_89_g 0 n0_241_4953  0.0174842 
iB00_90_v n1_333_5000 0  0.0174842 
iB00_90_g 0 n0_241_4986  0.0174842 
iB00_91_v n1_333_5183 0  0.0174842 
iB00_91_g 0 n0_241_5169  0.0174842 
iB00_92_v n1_333_5216 0  0.0174842 
iB00_92_g 0 n0_241_5202  0.0174842 
iB00_93_v n1_380_4967 0  0.0174842 
iB00_93_g 0 n0_241_4953  0.0174842 
iB00_94_v n1_380_5000 0  0.0174842 
iB00_94_g 0 n0_241_4986  0.0174842 
iB00_95_v n1_521_5000 0  0.0174842 
iB00_95_g 0 n0_429_5169  0.0174842 
iB00_96_v n1_521_5183 0  0.0174842 
iB00_96_g 0 n0_429_5169  0.0174842 
iB00_97_v n1_521_5216 0  0.0174842 
iB00_97_g 0 n0_429_5202  0.0174842 
iB00_98_v n1_2400_215 0  0.0174842 
iB00_98_g 0 n0_1646_201  0.0174842 
iB00_99_v n1_2400_248 0  0.0174842 
iB00_99_g 0 n0_1646_234  0.0174842 
iB00_100_v n1_2400_383 0  0.0174842 
iB00_100_g 0 n0_1646_417  0.0174842 
iB00_101_v n1_2400_431 0  0.0174842 
iB00_101_g 0 n0_1646_417  0.0174842 
iB00_102_v n1_2400_464 0  0.0174842 
iB00_102_g 0 n0_1646_450  0.0174842 
iB00_103_v n1_2400_647 0  0.0174842 
iB00_103_g 0 n0_1646_633  0.0174842 
iB00_104_v n1_2400_680 0  0.0174842 
iB00_104_g 0 n0_1646_666  0.0174842 
iB00_105_v n1_2400_863 0  0.0174842 
iB00_105_g 0 n0_1646_849  0.0174842 
iB00_106_v n1_2400_896 0  0.0174842 
iB00_106_g 0 n0_1646_882  0.0174842 
iB00_107_v n1_2400_1079 0  0.0174842 
iB00_107_g 0 n0_1646_1065  0.0174842 
iB00_108_v n1_2400_1112 0  0.0174842 
iB00_108_g 0 n0_1646_1098  0.0174842 
iB00_109_v n1_2400_1295 0  0.0174842 
iB00_109_g 0 n0_1646_1281  0.0174842 
iB00_110_v n1_2400_1328 0  0.0174842 
iB00_110_g 0 n0_1646_1314  0.0174842 
iB00_111_v n1_2400_1511 0  0.0174842 
iB00_111_g 0 n0_1646_1497  0.0174842 
iB00_112_v n1_2400_1544 0  0.0174842 
iB00_112_g 0 n0_1646_1530  0.0174842 
iB00_113_v n1_2400_1727 0  0.0174842 
iB00_113_g 0 n0_1554_1713  0.0174842 
iB00_114_v n1_2400_1760 0  0.0174842 
iB00_114_g 0 n0_1554_1760  0.0174842 
iB00_115_v n1_2400_1943 0  0.0174842 
iB00_115_g 0 n0_1554_1929  0.0174842 
iB00_116_v n1_2400_1976 0  0.0174842 
iB00_116_g 0 n0_2491_2793  0.0174842 
iB00_117_v n1_2400_2159 0  0.0174842 
iB00_117_g 0 n0_2491_2793  0.0174842 
iB00_118_v n1_2400_2192 0  0.0174842 
iB00_118_g 0 n0_2491_2793  0.0174842 
iB00_119_v n1_2400_2375 0  0.0174842 
iB00_119_g 0 n0_2491_2793  0.0174842 
iB00_120_v n1_2400_2408 0  0.0174842 
iB00_120_g 0 n0_2491_2793  0.0174842 
iB00_121_v n1_2400_2543 0  0.0174842 
iB00_121_g 0 n0_2491_2793  0.0174842 
iB00_122_v n1_2400_2591 0  0.0174842 
iB00_122_g 0 n0_2491_2793  0.0174842 
iB00_123_v n1_2400_2624 0  0.0174842 
iB00_123_g 0 n0_2491_2793  0.0174842 
iB00_124_v n1_2583_215 0  0.0174842 
iB00_124_g 0 n0_1646_201  0.0174842 
iB00_125_v n1_2583_248 0  0.0174842 
iB00_125_g 0 n0_1646_234  0.0174842 
iB00_126_v n1_2583_383 0  0.0174842 
iB00_126_g 0 n0_1646_417  0.0174842 
iB00_127_v n1_2771_215 0  0.0174842 
iB00_127_g 0 n0_3616_201  0.0174842 
iB00_128_v n1_2771_248 0  0.0174842 
iB00_128_g 0 n0_3616_234  0.0174842 
iB00_129_v n1_2771_383 0  0.0174842 
iB00_129_g 0 n0_3616_356  0.0174842 
iB00_130_v n1_2864_215 0  0.0174842 
iB00_130_g 0 n0_3616_201  0.0174842 
iB00_131_v n1_2864_248 0  0.0174842 
iB00_131_g 0 n0_3616_234  0.0174842 
iB00_132_v n1_2864_383 0  0.0174842 
iB00_132_g 0 n0_3616_356  0.0174842 
iB00_133_v n1_2583_431 0  0.0174842 
iB00_133_g 0 n0_1646_417  0.0174842 
iB00_134_v n1_2583_464 0  0.0174842 
iB00_134_g 0 n0_1646_450  0.0174842 
iB00_135_v n1_2583_647 0  0.0174842 
iB00_135_g 0 n0_1646_633  0.0174842 
iB00_136_v n1_2583_680 0  0.0174842 
iB00_136_g 0 n0_1646_666  0.0174842 
iB00_137_v n1_2630_431 0  0.0174842 
iB00_137_g 0 n0_3616_417  0.0174842 
iB00_138_v n1_2630_464 0  0.0174842 
iB00_138_g 0 n0_3616_450  0.0174842 
iB00_139_v n1_2771_431 0  0.0174842 
iB00_139_g 0 n0_3616_417  0.0174842 
iB00_140_v n1_2771_647 0  0.0174842 
iB00_140_g 0 n0_3616_633  0.0174842 
iB00_141_v n1_2771_680 0  0.0174842 
iB00_141_g 0 n0_3616_666  0.0174842 
iB00_142_v n1_2864_431 0  0.0174842 
iB00_142_g 0 n0_3616_417  0.0174842 
iB00_143_v n1_2864_464 0  0.0174842 
iB00_143_g 0 n0_3616_450  0.0174842 
iB00_144_v n1_2864_647 0  0.0174842 
iB00_144_g 0 n0_3616_633  0.0174842 
iB00_145_v n1_2864_680 0  0.0174842 
iB00_145_g 0 n0_3616_666  0.0174842 
iB00_146_v n1_2583_863 0  0.0174842 
iB00_146_g 0 n0_1646_849  0.0174842 
iB00_147_v n1_2583_896 0  0.0174842 
iB00_147_g 0 n0_1646_882  0.0174842 
iB00_148_v n1_2583_1079 0  0.0174842 
iB00_148_g 0 n0_1646_1065  0.0174842 
iB00_149_v n1_2583_1112 0  0.0174842 
iB00_149_g 0 n0_1646_1098  0.0174842 
iB00_150_v n1_2771_863 0  0.0174842 
iB00_150_g 0 n0_3616_849  0.0174842 
iB00_151_v n1_2771_896 0  0.0174842 
iB00_151_g 0 n0_3616_882  0.0174842 
iB00_152_v n1_2771_1079 0  0.0174842 
iB00_152_g 0 n0_3616_1065  0.0174842 
iB00_153_v n1_2771_1112 0  0.0174842 
iB00_153_g 0 n0_3616_1098  0.0174842 
iB00_154_v n1_2864_863 0  0.0174842 
iB00_154_g 0 n0_3616_849  0.0174842 
iB00_155_v n1_2864_896 0  0.0174842 
iB00_155_g 0 n0_3616_882  0.0174842 
iB00_156_v n1_2864_1079 0  0.0174842 
iB00_156_g 0 n0_3616_1065  0.0174842 
iB00_157_v n1_2864_1112 0  0.0174842 
iB00_157_g 0 n0_3616_1098  0.0174842 
iB00_158_v n1_2583_1295 0  0.0174842 
iB00_158_g 0 n0_1646_1281  0.0174842 
iB00_159_v n1_2583_1328 0  0.0174842 
iB00_159_g 0 n0_1646_1314  0.0174842 
iB00_160_v n1_2771_1295 0  0.0174842 
iB00_160_g 0 n0_3616_1281  0.0174842 
iB00_161_v n1_2771_1328 0  0.0174842 
iB00_161_g 0 n0_3616_1314  0.0174842 
iB00_162_v n1_2771_1511 0  0.0174842 
iB00_162_g 0 n0_3616_1497  0.0174842 
iB00_163_v n1_2771_1544 0  0.0174842 
iB00_163_g 0 n0_3616_1530  0.0174842 
iB00_164_v n1_2864_1295 0  0.0174842 
iB00_164_g 0 n0_3616_1281  0.0174842 
iB00_165_v n1_2864_1328 0  0.0174842 
iB00_165_g 0 n0_3616_1314  0.0174842 
iB00_166_v n1_2864_1511 0  0.0174842 
iB00_166_g 0 n0_3616_1497  0.0174842 
iB00_167_v n1_2864_1544 0  0.0174842 
iB00_167_g 0 n0_3616_1530  0.0174842 
iB00_168_v n1_2583_1727 0  0.0174842 
iB00_168_g 0 n0_1554_1713  0.0174842 
iB00_169_v n1_2583_1760 0  0.0174842 
iB00_169_g 0 n0_1554_1760  0.0174842 
iB00_170_v n1_2583_1943 0  0.0174842 
iB00_170_g 0 n0_2491_2793  0.0174842 
iB00_171_v n1_2583_1976 0  0.0174842 
iB00_171_g 0 n0_2491_2793  0.0174842 
iB00_172_v n1_2771_1727 0  0.0174842 
iB00_172_g 0 n0_3616_1713  0.0174842 
iB00_173_v n1_2771_1760 0  0.0174842 
iB00_173_g 0 n0_3616_1746  0.0174842 
iB00_174_v n1_2771_1943 0  0.0174842 
iB00_174_g 0 n0_3616_1929  0.0174842 
iB00_175_v n1_2771_1976 0  0.0174842 
iB00_175_g 0 n0_2679_2826  0.0174842 
iB00_176_v n1_2864_1727 0  0.0174842 
iB00_176_g 0 n0_3616_1713  0.0174842 
iB00_177_v n1_2864_1760 0  0.0174842 
iB00_177_g 0 n0_3616_1746  0.0174842 
iB00_178_v n1_2864_1943 0  0.0174842 
iB00_178_g 0 n0_3616_1929  0.0174842 
iB00_179_v n1_2864_1976 0  0.0174842 
iB00_179_g 0 n0_2679_2826  0.0174842 
iB00_180_v n1_2583_2159 0  0.0174842 
iB00_180_g 0 n0_2491_2793  0.0174842 
iB00_181_v n1_2583_2192 0  0.0174842 
iB00_181_g 0 n0_2491_2793  0.0174842 
iB00_182_v n1_2583_2375 0  0.0174842 
iB00_182_g 0 n0_2491_2793  0.0174842 
iB00_183_v n1_2583_2408 0  0.0174842 
iB00_183_g 0 n0_2491_2793  0.0174842 
iB00_184_v n1_2771_2159 0  0.0174842 
iB00_184_g 0 n0_2679_2826  0.0174842 
iB00_185_v n1_2771_2192 0  0.0174842 
iB00_185_g 0 n0_2679_2826  0.0174842 
iB00_186_v n1_2771_2375 0  0.0174842 
iB00_186_g 0 n0_2679_2826  0.0174842 
iB00_187_v n1_2771_2408 0  0.0174842 
iB00_187_g 0 n0_2679_2826  0.0174842 
iB00_188_v n1_2864_2159 0  0.0174842 
iB00_188_g 0 n0_2679_2826  0.0174842 
iB00_189_v n1_2864_2192 0  0.0174842 
iB00_189_g 0 n0_2679_2826  0.0174842 
iB00_190_v n1_2864_2375 0  0.0174842 
iB00_190_g 0 n0_2679_2826  0.0174842 
iB00_191_v n1_2864_2408 0  0.0174842 
iB00_191_g 0 n0_2679_2826  0.0174842 
iB00_192_v n1_2583_2543 0  0.0174842 
iB00_192_g 0 n0_2491_2793  0.0174842 
iB00_193_v n1_2583_2591 0  0.0174842 
iB00_193_g 0 n0_2491_2793  0.0174842 
iB00_194_v n1_2583_2624 0  0.0174842 
iB00_194_g 0 n0_2491_2793  0.0174842 
iB00_195_v n1_2583_2807 0  0.0174842 
iB00_195_g 0 n0_2491_2793  0.0174842 
iB00_196_v n1_2583_2840 0  0.0174842 
iB00_196_g 0 n0_2491_2826  0.0174842 
iB00_197_v n1_2771_2543 0  0.0174842 
iB00_197_g 0 n0_2679_2826  0.0174842 
iB00_198_v n1_2771_2591 0  0.0174842 
iB00_198_g 0 n0_2679_2826  0.0174842 
iB00_199_v n1_2771_2624 0  0.0174842 
iB00_199_g 0 n0_2679_2826  0.0174842 
iB00_200_v n1_2771_2807 0  0.0174842 
iB00_200_g 0 n0_2679_2826  0.0174842 
iB00_201_v n1_2771_2840 0  0.0174842 
iB00_201_g 0 n0_2679_2826  0.0174842 
iB00_202_v n1_2864_2543 0  0.0174842 
iB00_202_g 0 n0_2679_2826  0.0174842 
iB00_203_v n1_2864_2591 0  0.0174842 
iB00_203_g 0 n0_2679_2826  0.0174842 
iB00_204_v n1_2864_2624 0  0.0174842 
iB00_204_g 0 n0_2679_2826  0.0174842 
iB00_205_v n1_2583_3023 0  0.0174842 
iB00_205_g 0 n0_2491_3009  0.0174842 
iB00_206_v n1_2583_3056 0  0.0174842 
iB00_206_g 0 n0_2491_3042  0.0174842 
iB00_207_v n1_2583_3239 0  0.0174842 
iB00_207_g 0 n0_2491_3225  0.0174842 
iB00_208_v n1_2771_3023 0  0.0174842 
iB00_208_g 0 n0_2679_3009  0.0174842 
iB00_209_v n1_2771_3056 0  0.0174842 
iB00_209_g 0 n0_2679_3042  0.0174842 
iB00_210_v n1_2771_3239 0  0.0174842 
iB00_210_g 0 n0_2679_3225  0.0174842 
iB00_211_v n1_2583_3272 0  0.0174842 
iB00_211_g 0 n0_2491_3272  0.0174842 
iB00_212_v n1_2583_3428 0  0.0174842 
iB00_212_g 0 n0_2491_3441  0.0174842 
iB00_213_v n1_2583_3455 0  0.0174842 
iB00_213_g 0 n0_2491_3441  0.0174842 
iB00_214_v n1_2583_3488 0  0.0174842 
iB00_214_g 0 n0_2491_3474  0.0174842 
iB00_215_v n1_2583_3671 0  0.0174842 
iB00_215_g 0 n0_2491_3657  0.0174842 
iB00_216_v n1_2771_3272 0  0.0174842 
iB00_216_g 0 n0_2679_3272  0.0174842 
iB00_217_v n1_2771_3428 0  0.0174842 
iB00_217_g 0 n0_2679_3441  0.0174842 
iB00_218_v n1_2771_3455 0  0.0174842 
iB00_218_g 0 n0_2679_3441  0.0174842 
iB00_219_v n1_2771_3488 0  0.0174842 
iB00_219_g 0 n0_2679_3474  0.0174842 
iB00_220_v n1_2771_3671 0  0.0174842 
iB00_220_g 0 n0_2679_3657  0.0174842 
iB00_221_v n1_2583_3704 0  0.0174842 
iB00_221_g 0 n0_2491_3704  0.0174842 
iB00_222_v n1_2583_4076 0  0.0174842 
iB00_222_g 0 n0_2491_4089  0.0174842 
iB00_223_v n1_2771_3704 0  0.0174842 
iB00_223_g 0 n0_2679_3704  0.0174842 
iB00_224_v n1_2771_3860 0  0.0174842 
iB00_224_g 0 n0_2679_3873  0.0174842 
iB00_225_v n1_2771_3887 0  0.0174842 
iB00_225_g 0 n0_2679_3873  0.0174842 
iB00_226_v n1_2771_3920 0  0.0174842 
iB00_226_g 0 n0_2679_3920  0.0174842 
iB00_227_v n1_2771_4076 0  0.0174842 
iB00_227_g 0 n0_2679_4089  0.0174842 
iB00_228_v n1_2583_4103 0  0.0174842 
iB00_228_g 0 n0_2491_4089  0.0174842 
iB00_229_v n1_2583_4136 0  0.0174842 
iB00_229_g 0 n0_2491_4122  0.0174842 
iB00_230_v n1_2583_4270 0  0.0174842 
iB00_230_g 0 n0_2491_4305  0.0174842 
iB00_231_v n1_2583_4319 0  0.0174842 
iB00_231_g 0 n0_2491_4305  0.0174842 
iB00_232_v n1_2583_4352 0  0.0174842 
iB00_232_g 0 n0_2491_4352  0.0174842 
iB00_233_v n1_2771_4103 0  0.0174842 
iB00_233_g 0 n0_2679_4089  0.0174842 
iB00_234_v n1_2771_4136 0  0.0174842 
iB00_234_g 0 n0_2679_4122  0.0174842 
iB00_235_v n1_2771_4270 0  0.0174842 
iB00_235_g 0 n0_2679_4305  0.0174842 
iB00_236_v n1_2771_4319 0  0.0174842 
iB00_236_g 0 n0_2679_4305  0.0174842 
iB00_237_v n1_2771_4352 0  0.0174842 
iB00_237_g 0 n0_2679_4352  0.0174842 
iB00_238_v n1_2583_4508 0  0.0174842 
iB00_238_g 0 n0_2491_4521  0.0174842 
iB00_239_v n1_2583_4535 0  0.0174842 
iB00_239_g 0 n0_2491_4521  0.0174842 
iB00_240_v n1_2583_4568 0  0.0174842 
iB00_240_g 0 n0_2491_4554  0.0174842 
iB00_241_v n1_2583_4751 0  0.0174842 
iB00_241_g 0 n0_2491_4737  0.0174842 
iB00_242_v n1_2583_4784 0  0.0174842 
iB00_242_g 0 n0_2491_4770  0.0174842 
iB00_243_v n1_2771_4508 0  0.0174842 
iB00_243_g 0 n0_2679_4521  0.0174842 
iB00_244_v n1_2771_4535 0  0.0174842 
iB00_244_g 0 n0_2679_4521  0.0174842 
iB00_245_v n1_2771_4568 0  0.0174842 
iB00_245_g 0 n0_2679_4554  0.0174842 
iB00_246_v n1_2771_4751 0  0.0174842 
iB00_246_g 0 n0_2679_4737  0.0174842 
iB00_247_v n1_2771_4784 0  0.0174842 
iB00_247_g 0 n0_2679_4770  0.0174842 
iB00_248_v n1_2583_4967 0  0.0174842 
iB00_248_g 0 n0_2491_4953  0.0174842 
iB00_249_v n1_2583_5000 0  0.0174842 
iB00_249_g 0 n0_2491_4986  0.0174842 
iB00_250_v n1_2583_5183 0  0.0174842 
iB00_250_g 0 n0_2491_5169  0.0174842 
iB00_251_v n1_2583_5216 0  0.0174842 
iB00_251_g 0 n0_2491_5202  0.0174842 
iB00_252_v n1_2630_4967 0  0.0174842 
iB00_252_g 0 n0_2491_4953  0.0174842 
iB00_253_v n1_2630_5000 0  0.0174842 
iB00_253_g 0 n0_2491_4986  0.0174842 
iB00_254_v n1_2771_5000 0  0.0174842 
iB00_254_g 0 n0_2679_5169  0.0174842 
iB00_255_v n1_2771_5183 0  0.0174842 
iB00_255_g 0 n0_2679_5169  0.0174842 
iB00_256_v n1_2771_5216 0  0.0174842 
iB00_256_g 0 n0_2679_5202  0.0174842 
iB00_257_v n1_4650_215 0  0.0174842 
iB00_257_g 0 n0_3896_201  0.0174842 
iB00_258_v n1_4650_248 0  0.0174842 
iB00_258_g 0 n0_3896_234  0.0174842 
iB00_259_v n1_4833_215 0  0.0174842 
iB00_259_g 0 n0_3896_201  0.0174842 
iB00_260_v n1_4833_248 0  0.0174842 
iB00_260_g 0 n0_3896_234  0.0174842 
iB00_261_v n1_4650_431 0  0.0174842 
iB00_261_g 0 n0_3896_417  0.0174842 
iB00_262_v n1_4650_464 0  0.0174842 
iB00_262_g 0 n0_3896_450  0.0174842 
iB00_263_v n1_4650_513 0  0.0174842 
iB00_263_g 0 n0_3896_450  0.0174842 
iB00_264_v n1_4650_647 0  0.0174842 
iB00_264_g 0 n0_3896_633  0.0174842 
iB00_265_v n1_4650_680 0  0.0174842 
iB00_265_g 0 n0_3896_666  0.0174842 
iB00_266_v n1_4833_431 0  0.0174842 
iB00_266_g 0 n0_3896_417  0.0174842 
iB00_267_v n1_4833_464 0  0.0174842 
iB00_267_g 0 n0_3896_450  0.0174842 
iB00_268_v n1_4833_513 0  0.0174842 
iB00_268_g 0 n0_3896_450  0.0174842 
iB00_269_v n1_4833_647 0  0.0174842 
iB00_269_g 0 n0_3896_633  0.0174842 
iB00_270_v n1_4833_680 0  0.0174842 
iB00_270_g 0 n0_3896_666  0.0174842 
iB00_271_v n1_4880_431 0  0.0174842 
iB00_271_g 0 n0_3896_417  0.0174842 
iB00_272_v n1_4880_464 0  0.0174842 
iB00_272_g 0 n0_3896_450  0.0174842 
iB00_273_v n1_4880_513 0  0.0174842 
iB00_273_g 0 n0_3896_450  0.0174842 
iB00_274_v n1_4650_863 0  0.0174842 
iB00_274_g 0 n0_3896_849  0.0174842 
iB00_275_v n1_4650_896 0  0.0174842 
iB00_275_g 0 n0_3896_882  0.0174842 
iB00_276_v n1_4650_945 0  0.0174842 
iB00_276_g 0 n0_3896_882  0.0174842 
iB00_277_v n1_4650_1079 0  0.0174842 
iB00_277_g 0 n0_3896_1065  0.0174842 
iB00_278_v n1_4650_1112 0  0.0174842 
iB00_278_g 0 n0_3896_1098  0.0174842 
iB00_279_v n1_4833_863 0  0.0174842 
iB00_279_g 0 n0_3896_849  0.0174842 
iB00_280_v n1_4833_896 0  0.0174842 
iB00_280_g 0 n0_3896_882  0.0174842 
iB00_281_v n1_4833_945 0  0.0174842 
iB00_281_g 0 n0_3896_882  0.0174842 
iB00_282_v n1_4833_1079 0  0.0174842 
iB00_282_g 0 n0_3896_1065  0.0174842 
iB00_283_v n1_4833_1112 0  0.0174842 
iB00_283_g 0 n0_3896_1098  0.0174842 
iB00_284_v n1_4650_1295 0  0.0174842 
iB00_284_g 0 n0_3896_1281  0.0174842 
iB00_285_v n1_4650_1328 0  0.0174842 
iB00_285_g 0 n0_3896_1314  0.0174842 
iB00_286_v n1_4650_1511 0  0.0174842 
iB00_286_g 0 n0_3896_1497  0.0174842 
iB00_287_v n1_4650_1544 0  0.0174842 
iB00_287_g 0 n0_3896_1530  0.0174842 
iB00_288_v n1_4833_1295 0  0.0174842 
iB00_288_g 0 n0_3896_1281  0.0174842 
iB00_289_v n1_4833_1328 0  0.0174842 
iB00_289_g 0 n0_3896_1314  0.0174842 
iB00_290_v n1_4650_1727 0  0.0174842 
iB00_290_g 0 n0_3896_1713  0.0174842 
iB00_291_v n1_4650_1760 0  0.0174842 
iB00_291_g 0 n0_3896_1746  0.0174842 
iB00_292_v n1_4650_1943 0  0.0174842 
iB00_292_g 0 n0_3896_1929  0.0174842 
iB00_293_v n1_4650_1976 0  0.0174842 
iB00_293_g 0 n0_3896_1976  0.0174842 
iB00_294_v n1_4833_1727 0  0.0174842 
iB00_294_g 0 n0_3896_1713  0.0174842 
iB00_295_v n1_4833_1760 0  0.0174842 
iB00_295_g 0 n0_3896_1746  0.0174842 
iB00_296_v n1_4833_1916 0  0.0174842 
iB00_296_g 0 n0_3896_1929  0.0174842 
iB00_297_v n1_4833_1943 0  0.0174842 
iB00_297_g 0 n0_3896_1929  0.0174842 
iB00_298_v n1_4833_1976 0  0.0174842 
iB00_298_g 0 n0_3896_1976  0.0174842 
iB00_299_v n1_4650_2132 0  0.0174842 
iB00_299_g 0 n0_3896_2145  0.0174842 
iB00_300_v n1_4650_2159 0  0.0174842 
iB00_300_g 0 n0_3896_2145  0.0174842 
iB00_301_v n1_4650_2192 0  0.0174842 
iB00_301_g 0 n0_3896_2178  0.0174842 
iB00_302_v n1_4650_2375 0  0.0174842 
iB00_302_g 0 n0_3896_2361  0.0174842 
iB00_303_v n1_4650_2408 0  0.0174842 
iB00_303_g 0 n0_3896_2394  0.0174842 
iB00_304_v n1_4833_2132 0  0.0174842 
iB00_304_g 0 n0_3896_2145  0.0174842 
iB00_305_v n1_4833_2159 0  0.0174842 
iB00_305_g 0 n0_3896_2145  0.0174842 
iB00_306_v n1_4833_2192 0  0.0174842 
iB00_306_g 0 n0_3896_2178  0.0174842 
iB00_307_v n1_4833_2375 0  0.0174842 
iB00_307_g 0 n0_3896_2361  0.0174842 
iB00_308_v n1_4833_2408 0  0.0174842 
iB00_308_g 0 n0_3896_2394  0.0174842 
iB00_309_v n1_4650_2543 0  0.0174842 
iB00_309_g 0 n0_3896_2577  0.0174842 
iB00_310_v n1_4650_2591 0  0.0174842 
iB00_310_g 0 n0_3896_2577  0.0174842 
iB00_311_v n1_4650_2624 0  0.0174842 
iB00_311_g 0 n0_3896_2610  0.0174842 
iB00_312_v n1_4833_2543 0  0.0174842 
iB00_312_g 0 n0_3896_2577  0.0174842 
iB00_313_v n1_4833_2564 0  0.0174842 
iB00_313_g 0 n0_3896_2577  0.0174842 
iB00_314_v n1_4833_2591 0  0.0174842 
iB00_314_g 0 n0_3896_2577  0.0174842 
iB00_315_v n1_4833_2624 0  0.0174842 
iB00_315_g 0 n0_3896_2610  0.0174842 
iB00_316_v n1_4833_2807 0  0.0174842 
iB00_316_g 0 n0_3896_2793  0.0174842 
iB00_317_v n1_4833_2840 0  0.0174842 
iB00_317_g 0 n0_3896_2826  0.0174842 
iB00_318_v n1_4833_2996 0  0.0174842 
iB00_318_g 0 n0_3896_3009  0.0174842 
iB00_319_v n1_4833_3023 0  0.0174842 
iB00_319_g 0 n0_3896_3009  0.0174842 
iB00_320_v n1_4833_3056 0  0.0174842 
iB00_320_g 0 n0_3896_3042  0.0174842 
iB00_321_v n1_4833_3212 0  0.0174842 
iB00_321_g 0 n0_3896_3225  0.0174842 
iB00_322_v n1_4833_3239 0  0.0174842 
iB00_322_g 0 n0_3896_3225  0.0174842 
iB00_323_v n1_4833_3272 0  0.0174842 
iB00_323_g 0 n0_3896_3258  0.0174842 
iB00_324_v n1_4833_3455 0  0.0174842 
iB00_324_g 0 n0_3896_3441  0.0174842 
iB00_325_v n1_4833_3488 0  0.0174842 
iB00_325_g 0 n0_3896_3474  0.0174842 
iB00_326_v n1_4833_3644 0  0.0174842 
iB00_326_g 0 n0_3896_3657  0.0174842 
iB00_327_v n1_4833_3671 0  0.0174842 
iB00_327_g 0 n0_3896_3657  0.0174842 
iB00_328_v n1_4833_3704 0  0.0174842 
iB00_328_g 0 n0_3896_3704  0.0174842 
iB00_329_v n1_4833_4103 0  0.0174842 
iB00_329_g 0 n0_5866_4089  0.0174842 
iB00_330_v n1_4833_4136 0  0.0174842 
iB00_330_g 0 n0_5866_4136  0.0174842 
iB00_331_v n1_4833_4292 0  0.0174842 
iB00_331_g 0 n0_4741_5169  0.0174842 
iB00_332_v n1_4833_4319 0  0.0174842 
iB00_332_g 0 n0_4741_5169  0.0174842 
iB00_333_v n1_4833_4352 0  0.0174842 
iB00_333_g 0 n0_4741_5169  0.0174842 
iB00_334_v n1_4833_4486 0  0.0174842 
iB00_334_g 0 n0_4741_5169  0.0174842 
iB00_335_v n1_4833_4508 0  0.0174842 
iB00_335_g 0 n0_4741_5169  0.0174842 
iB00_336_v n1_4833_4535 0  0.0174842 
iB00_336_g 0 n0_4741_5169  0.0174842 
iB00_337_v n1_4833_4568 0  0.0174842 
iB00_337_g 0 n0_4741_5169  0.0174842 
iB00_338_v n1_4833_4751 0  0.0174842 
iB00_338_g 0 n0_4741_5169  0.0174842 
iB00_339_v n1_4833_4784 0  0.0174842 
iB00_339_g 0 n0_4741_5169  0.0174842 
iB00_340_v n1_4833_4967 0  0.0174842 
iB00_340_g 0 n0_4741_5169  0.0174842 
iB00_341_v n1_4833_5000 0  0.0174842 
iB00_341_g 0 n0_4741_5169  0.0174842 
iB00_342_v n1_4833_5183 0  0.0174842 
iB00_342_g 0 n0_4741_5169  0.0174842 
iB00_343_v n1_4833_5216 0  0.0174842 
iB00_343_g 0 n0_4741_5202  0.0174842 
iB00_344_v n1_4880_4967 0  0.0174842 
iB00_344_g 0 n0_4929_5169  0.0174842 
iB00_345_v n1_4880_5000 0  0.0174842 
iB00_345_g 0 n0_4929_5169  0.0174842 
iB00_346_v n1_5021_215 0  0.0174842 
iB00_346_g 0 n0_5866_201  0.0174842 
iB00_347_v n1_5021_248 0  0.0174842 
iB00_347_g 0 n0_5866_234  0.0174842 
iB00_348_v n1_5114_215 0  0.0174842 
iB00_348_g 0 n0_5866_201  0.0174842 
iB00_349_v n1_5114_248 0  0.0174842 
iB00_349_g 0 n0_5866_234  0.0174842 
iB00_350_v n1_5021_431 0  0.0174842 
iB00_350_g 0 n0_5866_417  0.0174842 
iB00_351_v n1_5021_513 0  0.0174842 
iB00_351_g 0 n0_5866_450  0.0174842 
iB00_352_v n1_5021_647 0  0.0174842 
iB00_352_g 0 n0_5866_633  0.0174842 
iB00_353_v n1_5021_680 0  0.0174842 
iB00_353_g 0 n0_5866_666  0.0174842 
iB00_354_v n1_5114_431 0  0.0174842 
iB00_354_g 0 n0_5866_417  0.0174842 
iB00_355_v n1_5114_464 0  0.0174842 
iB00_355_g 0 n0_5866_450  0.0174842 
iB00_356_v n1_5114_513 0  0.0174842 
iB00_356_g 0 n0_5866_450  0.0174842 
iB00_357_v n1_5114_647 0  0.0174842 
iB00_357_g 0 n0_5866_633  0.0174842 
iB00_358_v n1_5114_680 0  0.0174842 
iB00_358_g 0 n0_5866_666  0.0174842 
iB00_359_v n1_5021_863 0  0.0174842 
iB00_359_g 0 n0_5866_849  0.0174842 
iB00_360_v n1_5021_896 0  0.0174842 
iB00_360_g 0 n0_5866_882  0.0174842 
iB00_361_v n1_5021_945 0  0.0174842 
iB00_361_g 0 n0_5866_882  0.0174842 
iB00_362_v n1_5021_1079 0  0.0174842 
iB00_362_g 0 n0_5866_1065  0.0174842 
iB00_363_v n1_5021_1112 0  0.0174842 
iB00_363_g 0 n0_5866_1098  0.0174842 
iB00_364_v n1_5114_863 0  0.0174842 
iB00_364_g 0 n0_5866_849  0.0174842 
iB00_365_v n1_5114_896 0  0.0174842 
iB00_365_g 0 n0_5866_882  0.0174842 
iB00_366_v n1_5114_945 0  0.0174842 
iB00_366_g 0 n0_5866_882  0.0174842 
iB00_367_v n1_5114_1079 0  0.0174842 
iB00_367_g 0 n0_5866_1065  0.0174842 
iB00_368_v n1_5114_1112 0  0.0174842 
iB00_368_g 0 n0_5866_1098  0.0174842 
iB00_369_v n1_5021_1295 0  0.0174842 
iB00_369_g 0 n0_5866_1281  0.0174842 
iB00_370_v n1_5021_1328 0  0.0174842 
iB00_370_g 0 n0_5866_1314  0.0174842 
iB00_371_v n1_5021_1511 0  0.0174842 
iB00_371_g 0 n0_5866_1497  0.0174842 
iB00_372_v n1_5021_1544 0  0.0174842 
iB00_372_g 0 n0_5866_1530  0.0174842 
iB00_373_v n1_5114_1295 0  0.0174842 
iB00_373_g 0 n0_5866_1281  0.0174842 
iB00_374_v n1_5114_1328 0  0.0174842 
iB00_374_g 0 n0_5866_1314  0.0174842 
iB00_375_v n1_5114_1511 0  0.0174842 
iB00_375_g 0 n0_5866_1497  0.0174842 
iB00_376_v n1_5114_1544 0  0.0174842 
iB00_376_g 0 n0_5866_1530  0.0174842 
iB00_377_v n1_5021_1727 0  0.0174842 
iB00_377_g 0 n0_5866_1713  0.0174842 
iB00_378_v n1_5021_1760 0  0.0174842 
iB00_378_g 0 n0_5866_1760  0.0174842 
iB00_379_v n1_5021_1916 0  0.0174842 
iB00_379_g 0 n0_5866_1929  0.0174842 
iB00_380_v n1_5021_1943 0  0.0174842 
iB00_380_g 0 n0_5866_1929  0.0174842 
iB00_381_v n1_5021_1976 0  0.0174842 
iB00_381_g 0 n0_5866_1962  0.0174842 
iB00_382_v n1_5114_1727 0  0.0174842 
iB00_382_g 0 n0_5866_1713  0.0174842 
iB00_383_v n1_5114_1760 0  0.0174842 
iB00_383_g 0 n0_5866_1760  0.0174842 
iB00_384_v n1_5114_1916 0  0.0174842 
iB00_384_g 0 n0_5866_1929  0.0174842 
iB00_385_v n1_5114_1943 0  0.0174842 
iB00_385_g 0 n0_5866_1929  0.0174842 
iB00_386_v n1_5114_1976 0  0.0174842 
iB00_386_g 0 n0_5866_1962  0.0174842 
iB00_387_v n1_5021_2132 0  0.0174842 
iB00_387_g 0 n0_5866_2145  0.0174842 
iB00_388_v n1_5021_2159 0  0.0174842 
iB00_388_g 0 n0_5866_2145  0.0174842 
iB00_389_v n1_5021_2192 0  0.0174842 
iB00_389_g 0 n0_5866_2178  0.0174842 
iB00_390_v n1_5021_2375 0  0.0174842 
iB00_390_g 0 n0_5866_2361  0.0174842 
iB00_391_v n1_5021_2408 0  0.0174842 
iB00_391_g 0 n0_5866_2408  0.0174842 
iB00_392_v n1_5114_2159 0  0.0174842 
iB00_392_g 0 n0_5866_2145  0.0174842 
iB00_393_v n1_5114_2192 0  0.0174842 
iB00_393_g 0 n0_5866_2178  0.0174842 
iB00_394_v n1_5114_2375 0  0.0174842 
iB00_394_g 0 n0_5866_2361  0.0174842 
iB00_395_v n1_5114_2408 0  0.0174842 
iB00_395_g 0 n0_5866_2408  0.0174842 
iB00_396_v n1_5021_2543 0  0.0174842 
iB00_396_g 0 n0_5866_2577  0.0174842 
iB00_397_v n1_5021_2564 0  0.0174842 
iB00_397_g 0 n0_5866_2577  0.0174842 
iB00_398_v n1_5021_2591 0  0.0174842 
iB00_398_g 0 n0_5866_2577  0.0174842 
iB00_399_v n1_5021_2624 0  0.0174842 
iB00_399_g 0 n0_5866_2610  0.0174842 
iB00_400_v n1_5021_2807 0  0.0174842 
iB00_400_g 0 n0_5866_2793  0.0174842 
iB00_401_v n1_5021_2840 0  0.0174842 
iB00_401_g 0 n0_5866_2840  0.0174842 
iB00_402_v n1_5114_2543 0  0.0174842 
iB00_402_g 0 n0_5866_2577  0.0174842 
iB00_403_v n1_5114_2564 0  0.0174842 
iB00_403_g 0 n0_5866_2577  0.0174842 
iB00_404_v n1_5114_2591 0  0.0174842 
iB00_404_g 0 n0_5866_2577  0.0174842 
iB00_405_v n1_5114_2624 0  0.0174842 
iB00_405_g 0 n0_5866_2610  0.0174842 
iB00_406_v n1_5021_2996 0  0.0174842 
iB00_406_g 0 n0_5866_3009  0.0174842 
iB00_407_v n1_5021_3023 0  0.0174842 
iB00_407_g 0 n0_5866_3009  0.0174842 
iB00_408_v n1_5021_3056 0  0.0174842 
iB00_408_g 0 n0_5866_3056  0.0174842 
iB00_409_v n1_5021_3212 0  0.0174842 
iB00_409_g 0 n0_5866_3225  0.0174842 
iB00_410_v n1_5021_3239 0  0.0174842 
iB00_410_g 0 n0_5866_3225  0.0174842 
iB00_411_v n1_5021_3272 0  0.0174842 
iB00_411_g 0 n0_5866_3258  0.0174842 
iB00_412_v n1_5021_3455 0  0.0174842 
iB00_412_g 0 n0_5866_3441  0.0174842 
iB00_413_v n1_5021_3488 0  0.0174842 
iB00_413_g 0 n0_5866_3488  0.0174842 
iB00_414_v n1_5021_3644 0  0.0174842 
iB00_414_g 0 n0_5866_3657  0.0174842 
iB00_415_v n1_5021_3671 0  0.0174842 
iB00_415_g 0 n0_5866_3657  0.0174842 
iB00_416_v n1_5021_3704 0  0.0174842 
iB00_416_g 0 n0_5866_3690  0.0174842 
iB00_417_v n1_5021_3887 0  0.0174842 
iB00_417_g 0 n0_5866_3873  0.0174842 
iB00_418_v n1_5021_3920 0  0.0174842 
iB00_418_g 0 n0_5866_3906  0.0174842 
iB00_419_v n1_5021_4103 0  0.0174842 
iB00_419_g 0 n0_5866_4089  0.0174842 
iB00_420_v n1_5021_4136 0  0.0174842 
iB00_420_g 0 n0_5866_4136  0.0174842 
iB00_421_v n1_5021_4292 0  0.0174842 
iB00_421_g 0 n0_5866_4305  0.0174842 
iB00_422_v n1_5021_4319 0  0.0174842 
iB00_422_g 0 n0_5866_4305  0.0174842 
iB00_423_v n1_5021_4352 0  0.0174842 
iB00_423_g 0 n0_5866_4352  0.0174842 
iB00_424_v n1_5021_4486 0  0.0174842 
iB00_424_g 0 n0_4929_5169  0.0174842 
iB00_425_v n1_5021_4508 0  0.0174842 
iB00_425_g 0 n0_4929_5169  0.0174842 
iB00_426_v n1_5021_4535 0  0.0174842 
iB00_426_g 0 n0_4929_5169  0.0174842 
iB00_427_v n1_5021_4568 0  0.0174842 
iB00_427_g 0 n0_4929_5169  0.0174842 
iB00_428_v n1_5021_4751 0  0.0174842 
iB00_428_g 0 n0_4929_5169  0.0174842 
iB00_429_v n1_5021_4784 0  0.0174842 
iB00_429_g 0 n0_4929_5169  0.0174842 
iB00_430_v n1_5021_5000 0  0.0174842 
iB00_430_g 0 n0_4929_5169  0.0174842 
iB00_431_v n1_5021_5183 0  0.0174842 
iB00_431_g 0 n0_4929_5169  0.0174842 
iB00_432_v n1_5021_5216 0  0.0174842 
iB00_432_g 0 n0_4929_5202  0.0174842 
iB01_0_v n1_333_5399 0  0.0191987 
iB01_0_g 0 n0_241_5385  0.0191987 
iB01_1_v n1_333_5432 0  0.0191987 
iB01_1_g 0 n0_241_5418  0.0191987 
iB01_2_v n1_333_5615 0  0.0191987 
iB01_2_g 0 n0_241_5601  0.0191987 
iB01_3_v n1_333_5648 0  0.0191987 
iB01_3_g 0 n0_241_5634  0.0191987 
iB01_4_v n1_521_5399 0  0.0191987 
iB01_4_g 0 n0_429_5385  0.0191987 
iB01_5_v n1_521_5432 0  0.0191987 
iB01_5_g 0 n0_429_5418  0.0191987 
iB01_6_v n1_521_5615 0  0.0191987 
iB01_6_g 0 n0_429_5601  0.0191987 
iB01_7_v n1_521_5648 0  0.0191987 
iB01_7_g 0 n0_429_5634  0.0191987 
iB01_8_v n1_333_5831 0  0.0191987 
iB01_8_g 0 n0_241_5817  0.0191987 
iB01_9_v n1_333_5864 0  0.0191987 
iB01_9_g 0 n0_241_5850  0.0191987 
iB01_10_v n1_521_5831 0  0.0191987 
iB01_10_g 0 n0_429_5817  0.0191987 
iB01_11_v n1_521_5864 0  0.0191987 
iB01_11_g 0 n0_429_5850  0.0191987 
iB01_12_v n1_521_6047 0  0.0191987 
iB01_12_g 0 n0_429_6033  0.0191987 
iB01_13_v n1_521_6080 0  0.0191987 
iB01_13_g 0 n0_429_6066  0.0191987 
iB01_14_v n1_333_6263 0  0.0191987 
iB01_14_g 0 n0_241_6249  0.0191987 
iB01_15_v n1_333_6296 0  0.0191987 
iB01_15_g 0 n0_241_6282  0.0191987 
iB01_16_v n1_333_6479 0  0.0191987 
iB01_16_g 0 n0_241_6465  0.0191987 
iB01_17_v n1_333_6512 0  0.0191987 
iB01_17_g 0 n0_241_6498  0.0191987 
iB01_18_v n1_521_6263 0  0.0191987 
iB01_18_g 0 n0_429_6249  0.0191987 
iB01_19_v n1_521_6296 0  0.0191987 
iB01_19_g 0 n0_429_6282  0.0191987 
iB01_20_v n1_521_6479 0  0.0191987 
iB01_20_g 0 n0_429_6465  0.0191987 
iB01_21_v n1_521_6512 0  0.0191987 
iB01_21_g 0 n0_429_6498  0.0191987 
iB01_22_v n1_333_6695 0  0.0191987 
iB01_22_g 0 n0_241_6681  0.0191987 
iB01_23_v n1_333_6728 0  0.0191987 
iB01_23_g 0 n0_241_6714  0.0191987 
iB01_24_v n1_333_6911 0  0.0191987 
iB01_24_g 0 n0_241_6897  0.0191987 
iB01_25_v n1_521_6695 0  0.0191987 
iB01_25_g 0 n0_429_6681  0.0191987 
iB01_26_v n1_521_6728 0  0.0191987 
iB01_26_g 0 n0_429_6714  0.0191987 
iB01_27_v n1_521_6911 0  0.0191987 
iB01_27_g 0 n0_429_6897  0.0191987 
iB01_28_v n1_333_6944 0  0.0191987 
iB01_28_g 0 n0_241_6930  0.0191987 
iB01_29_v n1_333_7127 0  0.0191987 
iB01_29_g 0 n0_241_7113  0.0191987 
iB01_30_v n1_333_7160 0  0.0191987 
iB01_30_g 0 n0_241_7146  0.0191987 
iB01_31_v n1_380_7160 0  0.0191987 
iB01_31_g 0 n0_429_7113  0.0191987 
iB01_32_v n1_521_6944 0  0.0191987 
iB01_32_g 0 n0_429_6930  0.0191987 
iB01_33_v n1_521_7127 0  0.0191987 
iB01_33_g 0 n0_429_7113  0.0191987 
iB01_34_v n1_521_7160 0  0.0191987 
iB01_34_g 0 n0_429_7113  0.0191987 
iB01_35_v n1_333_7343 0  0.0191987 
iB01_35_g 0 n0_241_7329  0.0191987 
iB01_36_v n1_333_7376 0  0.0191987 
iB01_36_g 0 n0_241_7362  0.0191987 
iB01_37_v n1_333_7559 0  0.0191987 
iB01_37_g 0 n0_241_7545  0.0191987 
iB01_38_v n1_333_7592 0  0.0191987 
iB01_38_g 0 n0_241_7578  0.0191987 
iB01_39_v n1_521_7343 0  0.0191987 
iB01_39_g 0 n0_429_7329  0.0191987 
iB01_40_v n1_521_7376 0  0.0191987 
iB01_40_g 0 n0_429_7362  0.0191987 
iB01_41_v n1_521_7559 0  0.0191987 
iB01_41_g 0 n0_429_7545  0.0191987 
iB01_42_v n1_521_7592 0  0.0191987 
iB01_42_g 0 n0_429_7578  0.0191987 
iB01_43_v n1_333_7775 0  0.0191987 
iB01_43_g 0 n0_241_7761  0.0191987 
iB01_44_v n1_333_7808 0  0.0191987 
iB01_44_g 0 n0_241_7794  0.0191987 
iB01_45_v n1_333_7991 0  0.0191987 
iB01_45_g 0 n0_241_7977  0.0191987 
iB01_46_v n1_333_8024 0  0.0191987 
iB01_46_g 0 n0_241_8010  0.0191987 
iB01_47_v n1_521_7775 0  0.0191987 
iB01_47_g 0 n0_429_7761  0.0191987 
iB01_48_v n1_521_7808 0  0.0191987 
iB01_48_g 0 n0_429_7794  0.0191987 
iB01_49_v n1_521_7991 0  0.0191987 
iB01_49_g 0 n0_429_7977  0.0191987 
iB01_50_v n1_521_8024 0  0.0191987 
iB01_50_g 0 n0_429_8010  0.0191987 
iB01_51_v n1_333_8207 0  0.0191987 
iB01_51_g 0 n0_241_8193  0.0191987 
iB01_52_v n1_333_8240 0  0.0191987 
iB01_52_g 0 n0_241_8226  0.0191987 
iB01_53_v n1_333_8456 0  0.0191987 
iB01_53_g 0 n0_380_8409  0.0191987 
iB01_54_v n1_521_8207 0  0.0191987 
iB01_54_g 0 n0_429_8193  0.0191987 
iB01_55_v n1_521_8240 0  0.0191987 
iB01_55_g 0 n0_429_8226  0.0191987 
iB01_56_v n1_521_8423 0  0.0191987 
iB01_56_g 0 n0_429_8409  0.0191987 
iB01_57_v n1_521_8456 0  0.0191987 
iB01_57_g 0 n0_429_8442  0.0191987 
iB01_58_v n1_333_8639 0  0.0191987 
iB01_58_g 0 n0_241_8625  0.0191987 
iB01_59_v n1_333_8672 0  0.0191987 
iB01_59_g 0 n0_241_8658  0.0191987 
iB01_60_v n1_333_8855 0  0.0191987 
iB01_60_g 0 n0_241_8841  0.0191987 
iB01_61_v n1_333_8888 0  0.0191987 
iB01_61_g 0 n0_241_8874  0.0191987 
iB01_62_v n1_521_8639 0  0.0191987 
iB01_62_g 0 n0_429_8625  0.0191987 
iB01_63_v n1_521_8672 0  0.0191987 
iB01_63_g 0 n0_429_8658  0.0191987 
iB01_64_v n1_521_8855 0  0.0191987 
iB01_64_g 0 n0_429_8841  0.0191987 
iB01_65_v n1_521_8888 0  0.0191987 
iB01_65_g 0 n0_429_8874  0.0191987 
iB01_66_v n1_333_9071 0  0.0191987 
iB01_66_g 0 n0_241_9057  0.0191987 
iB01_67_v n1_333_9104 0  0.0191987 
iB01_67_g 0 n0_241_9090  0.0191987 
iB01_68_v n1_333_9287 0  0.0191987 
iB01_68_g 0 n0_241_9273  0.0191987 
iB01_69_v n1_333_9320 0  0.0191987 
iB01_69_g 0 n0_241_9306  0.0191987 
iB01_70_v n1_521_9071 0  0.0191987 
iB01_70_g 0 n0_429_9057  0.0191987 
iB01_71_v n1_521_9104 0  0.0191987 
iB01_71_g 0 n0_429_9090  0.0191987 
iB01_72_v n1_521_9287 0  0.0191987 
iB01_72_g 0 n0_429_9273  0.0191987 
iB01_73_v n1_521_9320 0  0.0191987 
iB01_73_g 0 n0_429_9306  0.0191987 
iB01_74_v n1_333_9503 0  0.0191987 
iB01_74_g 0 n0_241_9489  0.0191987 
iB01_75_v n1_333_9536 0  0.0191987 
iB01_75_g 0 n0_241_9522  0.0191987 
iB01_76_v n1_333_9719 0  0.0191987 
iB01_76_g 0 n0_241_9705  0.0191987 
iB01_77_v n1_333_9752 0  0.0191987 
iB01_77_g 0 n0_241_9738  0.0191987 
iB01_78_v n1_380_9503 0  0.0191987 
iB01_78_g 0 n0_241_9489  0.0191987 
iB01_79_v n1_380_9536 0  0.0191987 
iB01_79_g 0 n0_241_9522  0.0191987 
iB01_80_v n1_521_9503 0  0.0191987 
iB01_80_g 0 n0_429_9306  0.0191987 
iB01_81_v n1_521_9536 0  0.0191987 
iB01_81_g 0 n0_429_9705  0.0191987 
iB01_82_v n1_521_9719 0  0.0191987 
iB01_82_g 0 n0_429_9705  0.0191987 
iB01_83_v n1_521_9752 0  0.0191987 
iB01_83_g 0 n0_429_9738  0.0191987 
iB01_84_v n1_333_9935 0  0.0191987 
iB01_84_g 0 n0_241_9921  0.0191987 
iB01_85_v n1_333_9968 0  0.0191987 
iB01_85_g 0 n0_241_9954  0.0191987 
iB01_86_v n1_333_10151 0  0.0191987 
iB01_86_g 0 n0_241_10137  0.0191987 
iB01_87_v n1_333_10184 0  0.0191987 
iB01_87_g 0 n0_241_10170  0.0191987 
iB01_88_v n1_521_9935 0  0.0191987 
iB01_88_g 0 n0_429_9921  0.0191987 
iB01_89_v n1_521_9968 0  0.0191987 
iB01_89_g 0 n0_429_9954  0.0191987 
iB01_90_v n1_521_10151 0  0.0191987 
iB01_90_g 0 n0_429_10137  0.0191987 
iB01_91_v n1_521_10184 0  0.0191987 
iB01_91_g 0 n0_429_10170  0.0191987 
iB01_92_v n1_333_10367 0  0.0191987 
iB01_92_g 0 n0_241_10353  0.0191987 
iB01_93_v n1_333_10400 0  0.0191987 
iB01_93_g 0 n0_241_10386  0.0191987 
iB01_94_v n1_521_10367 0  0.0191987 
iB01_94_g 0 n0_429_10353  0.0191987 
iB01_95_v n1_521_10400 0  0.0191987 
iB01_95_g 0 n0_429_10386  0.0191987 
iB01_96_v n1_521_10616 0  0.0191987 
iB01_96_g 0 n0_429_10602  0.0191987 
iB01_97_v n1_2583_5399 0  0.0191987 
iB01_97_g 0 n0_2491_5385  0.0191987 
iB01_98_v n1_2583_5432 0  0.0191987 
iB01_98_g 0 n0_2491_5432  0.0191987 
iB01_99_v n1_2583_5446 0  0.0191987 
iB01_99_g 0 n0_2491_5432  0.0191987 
iB01_100_v n1_2583_5588 0  0.0191987 
iB01_100_g 0 n0_2491_5601  0.0191987 
iB01_101_v n1_2583_5615 0  0.0191987 
iB01_101_g 0 n0_2491_5601  0.0191987 
iB01_102_v n1_2583_5648 0  0.0191987 
iB01_102_g 0 n0_2491_5634  0.0191987 
iB01_103_v n1_2771_5399 0  0.0191987 
iB01_103_g 0 n0_2679_5385  0.0191987 
iB01_104_v n1_2771_5432 0  0.0191987 
iB01_104_g 0 n0_2679_5432  0.0191987 
iB01_105_v n1_2771_5446 0  0.0191987 
iB01_105_g 0 n0_2679_5432  0.0191987 
iB01_106_v n1_2771_5588 0  0.0191987 
iB01_106_g 0 n0_2679_5601  0.0191987 
iB01_107_v n1_2771_5615 0  0.0191987 
iB01_107_g 0 n0_2679_5601  0.0191987 
iB01_108_v n1_2771_5648 0  0.0191987 
iB01_108_g 0 n0_2679_5634  0.0191987 
iB01_109_v n1_2583_5831 0  0.0191987 
iB01_109_g 0 n0_2491_5817  0.0191987 
iB01_110_v n1_2583_5864 0  0.0191987 
iB01_110_g 0 n0_2491_5850  0.0191987 
iB01_111_v n1_2771_5831 0  0.0191987 
iB01_111_g 0 n0_2679_5817  0.0191987 
iB01_112_v n1_2771_5864 0  0.0191987 
iB01_112_g 0 n0_2679_5850  0.0191987 
iB01_113_v n1_2771_6047 0  0.0191987 
iB01_113_g 0 n0_2679_6033  0.0191987 
iB01_114_v n1_2771_6080 0  0.0191987 
iB01_114_g 0 n0_2679_6066  0.0191987 
iB01_115_v n1_2583_6263 0  0.0191987 
iB01_115_g 0 n0_2491_6249  0.0191987 
iB01_116_v n1_2583_6296 0  0.0191987 
iB01_116_g 0 n0_2491_6282  0.0191987 
iB01_117_v n1_2583_6479 0  0.0191987 
iB01_117_g 0 n0_2491_6465  0.0191987 
iB01_118_v n1_2583_6512 0  0.0191987 
iB01_118_g 0 n0_2491_6498  0.0191987 
iB01_119_v n1_2771_6263 0  0.0191987 
iB01_119_g 0 n0_2679_6249  0.0191987 
iB01_120_v n1_2771_6296 0  0.0191987 
iB01_120_g 0 n0_2679_6282  0.0191987 
iB01_121_v n1_2771_6479 0  0.0191987 
iB01_121_g 0 n0_2679_6465  0.0191987 
iB01_122_v n1_2771_6512 0  0.0191987 
iB01_122_g 0 n0_2679_6498  0.0191987 
iB01_123_v n1_2583_6549 0  0.0191987 
iB01_123_g 0 n0_2491_6535  0.0191987 
iB01_124_v n1_2583_6646 0  0.0191987 
iB01_124_g 0 n0_2491_6681  0.0191987 
iB01_125_v n1_2583_6695 0  0.0191987 
iB01_125_g 0 n0_2491_6681  0.0191987 
iB01_126_v n1_2583_6728 0  0.0191987 
iB01_126_g 0 n0_2491_6714  0.0191987 
iB01_127_v n1_2583_6911 0  0.0191987 
iB01_127_g 0 n0_2491_6897  0.0191987 
iB01_128_v n1_2771_6549 0  0.0191987 
iB01_128_g 0 n0_2679_6535  0.0191987 
iB01_129_v n1_2771_6646 0  0.0191987 
iB01_129_g 0 n0_2679_6681  0.0191987 
iB01_130_v n1_2771_6695 0  0.0191987 
iB01_130_g 0 n0_2679_6681  0.0191987 
iB01_131_v n1_2771_6728 0  0.0191987 
iB01_131_g 0 n0_2679_6714  0.0191987 
iB01_132_v n1_2771_6911 0  0.0191987 
iB01_132_g 0 n0_2679_6897  0.0191987 
iB01_133_v n1_2583_6944 0  0.0191987 
iB01_133_g 0 n0_2491_6930  0.0191987 
iB01_134_v n1_2583_7127 0  0.0191987 
iB01_134_g 0 n0_2491_7113  0.0191987 
iB01_135_v n1_2583_7160 0  0.0191987 
iB01_135_g 0 n0_2491_7146  0.0191987 
iB01_136_v n1_2630_7160 0  0.0191987 
iB01_136_g 0 n0_2679_7113  0.0191987 
iB01_137_v n1_2771_6944 0  0.0191987 
iB01_137_g 0 n0_2679_6930  0.0191987 
iB01_138_v n1_2771_7127 0  0.0191987 
iB01_138_g 0 n0_2679_7113  0.0191987 
iB01_139_v n1_2771_7160 0  0.0191987 
iB01_139_g 0 n0_2679_7113  0.0191987 
iB01_140_v n1_2583_7343 0  0.0191987 
iB01_140_g 0 n0_2491_7329  0.0191987 
iB01_141_v n1_2583_7376 0  0.0191987 
iB01_141_g 0 n0_2491_7362  0.0191987 
iB01_142_v n1_2583_7559 0  0.0191987 
iB01_142_g 0 n0_2491_7545  0.0191987 
iB01_143_v n1_2583_7592 0  0.0191987 
iB01_143_g 0 n0_2491_7578  0.0191987 
iB01_144_v n1_2771_7343 0  0.0191987 
iB01_144_g 0 n0_2679_7329  0.0191987 
iB01_145_v n1_2771_7376 0  0.0191987 
iB01_145_g 0 n0_2679_7362  0.0191987 
iB01_146_v n1_2771_7559 0  0.0191987 
iB01_146_g 0 n0_2679_7545  0.0191987 
iB01_147_v n1_2771_7592 0  0.0191987 
iB01_147_g 0 n0_2679_7578  0.0191987 
iB01_148_v n1_2583_7775 0  0.0191987 
iB01_148_g 0 n0_2491_7761  0.0191987 
iB01_149_v n1_2583_7808 0  0.0191987 
iB01_149_g 0 n0_2491_7808  0.0191987 
iB01_150_v n1_2583_7822 0  0.0191987 
iB01_150_g 0 n0_2491_7808  0.0191987 
iB01_151_v n1_2583_7964 0  0.0191987 
iB01_151_g 0 n0_2491_7977  0.0191987 
iB01_152_v n1_2583_7991 0  0.0191987 
iB01_152_g 0 n0_2491_7977  0.0191987 
iB01_153_v n1_2583_8024 0  0.0191987 
iB01_153_g 0 n0_2491_8010  0.0191987 
iB01_154_v n1_2771_7775 0  0.0191987 
iB01_154_g 0 n0_2679_7761  0.0191987 
iB01_155_v n1_2771_7808 0  0.0191987 
iB01_155_g 0 n0_2679_7808  0.0191987 
iB01_156_v n1_2771_7822 0  0.0191987 
iB01_156_g 0 n0_2679_7808  0.0191987 
iB01_157_v n1_2771_7964 0  0.0191987 
iB01_157_g 0 n0_2679_7977  0.0191987 
iB01_158_v n1_2771_7991 0  0.0191987 
iB01_158_g 0 n0_2679_7977  0.0191987 
iB01_159_v n1_2771_8024 0  0.0191987 
iB01_159_g 0 n0_2679_8010  0.0191987 
iB01_160_v n1_2583_8207 0  0.0191987 
iB01_160_g 0 n0_2491_8193  0.0191987 
iB01_161_v n1_2583_8240 0  0.0191987 
iB01_161_g 0 n0_2491_8226  0.0191987 
iB01_162_v n1_2583_8456 0  0.0191987 
iB01_162_g 0 n0_2630_8409  0.0191987 
iB01_163_v n1_2771_8207 0  0.0191987 
iB01_163_g 0 n0_2679_8193  0.0191987 
iB01_164_v n1_2771_8240 0  0.0191987 
iB01_164_g 0 n0_2679_8226  0.0191987 
iB01_165_v n1_2771_8423 0  0.0191987 
iB01_165_g 0 n0_2679_8409  0.0191987 
iB01_166_v n1_2771_8456 0  0.0191987 
iB01_166_g 0 n0_2679_8442  0.0191987 
iB01_167_v n1_2583_8639 0  0.0191987 
iB01_167_g 0 n0_2491_8625  0.0191987 
iB01_168_v n1_2583_8672 0  0.0191987 
iB01_168_g 0 n0_2491_8658  0.0191987 
iB01_169_v n1_2583_8855 0  0.0191987 
iB01_169_g 0 n0_2491_8841  0.0191987 
iB01_170_v n1_2583_8888 0  0.0191987 
iB01_170_g 0 n0_2491_8888  0.0191987 
iB01_171_v n1_2583_8902 0  0.0191987 
iB01_171_g 0 n0_2491_8911  0.0191987 
iB01_172_v n1_2771_8639 0  0.0191987 
iB01_172_g 0 n0_2679_8625  0.0191987 
iB01_173_v n1_2771_8672 0  0.0191987 
iB01_173_g 0 n0_2679_8658  0.0191987 
iB01_174_v n1_2771_8855 0  0.0191987 
iB01_174_g 0 n0_2679_8841  0.0191987 
iB01_175_v n1_2771_8888 0  0.0191987 
iB01_175_g 0 n0_2679_8888  0.0191987 
iB01_176_v n1_2771_8902 0  0.0191987 
iB01_176_g 0 n0_2679_8911  0.0191987 
iB01_177_v n1_2583_9022 0  0.0191987 
iB01_177_g 0 n0_2491_9057  0.0191987 
iB01_178_v n1_2583_9044 0  0.0191987 
iB01_178_g 0 n0_2491_9057  0.0191987 
iB01_179_v n1_2583_9071 0  0.0191987 
iB01_179_g 0 n0_2491_9057  0.0191987 
iB01_180_v n1_2583_9104 0  0.0191987 
iB01_180_g 0 n0_2491_9090  0.0191987 
iB01_181_v n1_2583_9287 0  0.0191987 
iB01_181_g 0 n0_2491_9273  0.0191987 
iB01_182_v n1_2583_9320 0  0.0191987 
iB01_182_g 0 n0_2491_9306  0.0191987 
iB01_183_v n1_2771_9022 0  0.0191987 
iB01_183_g 0 n0_2679_9057  0.0191987 
iB01_184_v n1_2771_9044 0  0.0191987 
iB01_184_g 0 n0_2679_9057  0.0191987 
iB01_185_v n1_2771_9071 0  0.0191987 
iB01_185_g 0 n0_2679_9057  0.0191987 
iB01_186_v n1_2771_9104 0  0.0191987 
iB01_186_g 0 n0_2679_9090  0.0191987 
iB01_187_v n1_2771_9287 0  0.0191987 
iB01_187_g 0 n0_2679_9273  0.0191987 
iB01_188_v n1_2771_9320 0  0.0191987 
iB01_188_g 0 n0_2679_9306  0.0191987 
iB01_189_v n1_2583_9503 0  0.0191987 
iB01_189_g 0 n0_2491_9489  0.0191987 
iB01_190_v n1_2583_9536 0  0.0191987 
iB01_190_g 0 n0_2491_9522  0.0191987 
iB01_191_v n1_2583_9719 0  0.0191987 
iB01_191_g 0 n0_2491_9705  0.0191987 
iB01_192_v n1_2583_9752 0  0.0191987 
iB01_192_g 0 n0_2491_9738  0.0191987 
iB01_193_v n1_2630_9503 0  0.0191987 
iB01_193_g 0 n0_2491_9489  0.0191987 
iB01_194_v n1_2630_9536 0  0.0191987 
iB01_194_g 0 n0_2491_9522  0.0191987 
iB01_195_v n1_2771_9503 0  0.0191987 
iB01_195_g 0 n0_2679_9306  0.0191987 
iB01_196_v n1_2771_9536 0  0.0191987 
iB01_196_g 0 n0_2679_9705  0.0191987 
iB01_197_v n1_2771_9719 0  0.0191987 
iB01_197_g 0 n0_2679_9705  0.0191987 
iB01_198_v n1_2771_9752 0  0.0191987 
iB01_198_g 0 n0_2679_9738  0.0191987 
iB01_199_v n1_2583_9935 0  0.0191987 
iB01_199_g 0 n0_2491_9921  0.0191987 
iB01_200_v n1_2583_9968 0  0.0191987 
iB01_200_g 0 n0_2491_9968  0.0191987 
iB01_201_v n1_2583_9982 0  0.0191987 
iB01_201_g 0 n0_2491_9968  0.0191987 
iB01_202_v n1_2583_10124 0  0.0191987 
iB01_202_g 0 n0_2491_10137  0.0191987 
iB01_203_v n1_2583_10151 0  0.0191987 
iB01_203_g 0 n0_2491_10137  0.0191987 
iB01_204_v n1_2583_10184 0  0.0191987 
iB01_204_g 0 n0_2491_10170  0.0191987 
iB01_205_v n1_2771_9935 0  0.0191987 
iB01_205_g 0 n0_2679_9921  0.0191987 
iB01_206_v n1_2771_9968 0  0.0191987 
iB01_206_g 0 n0_2679_9968  0.0191987 
iB01_207_v n1_2771_9982 0  0.0191987 
iB01_207_g 0 n0_2679_9968  0.0191987 
iB01_208_v n1_2771_10124 0  0.0191987 
iB01_208_g 0 n0_2679_10137  0.0191987 
iB01_209_v n1_2771_10151 0  0.0191987 
iB01_209_g 0 n0_2679_10137  0.0191987 
iB01_210_v n1_2771_10184 0  0.0191987 
iB01_210_g 0 n0_2679_10170  0.0191987 
iB01_211_v n1_2583_10367 0  0.0191987 
iB01_211_g 0 n0_2491_10353  0.0191987 
iB01_212_v n1_2583_10400 0  0.0191987 
iB01_212_g 0 n0_2491_10386  0.0191987 
iB01_213_v n1_2771_10367 0  0.0191987 
iB01_213_g 0 n0_2679_10353  0.0191987 
iB01_214_v n1_2771_10400 0  0.0191987 
iB01_214_g 0 n0_2679_10386  0.0191987 
iB01_215_v n1_2771_10616 0  0.0191987 
iB01_215_g 0 n0_2679_10602  0.0191987 
iB01_216_v n1_4833_5399 0  0.0191987 
iB01_216_g 0 n0_4741_5385  0.0191987 
iB01_217_v n1_4833_5432 0  0.0191987 
iB01_217_g 0 n0_4741_5432  0.0191987 
iB01_218_v n1_4833_5446 0  0.0191987 
iB01_218_g 0 n0_4741_5432  0.0191987 
iB01_219_v n1_4833_5588 0  0.0191987 
iB01_219_g 0 n0_4741_5601  0.0191987 
iB01_220_v n1_4833_5615 0  0.0191987 
iB01_220_g 0 n0_4741_5601  0.0191987 
iB01_221_v n1_4833_5648 0  0.0191987 
iB01_221_g 0 n0_4741_5634  0.0191987 
iB01_222_v n1_4833_5831 0  0.0191987 
iB01_222_g 0 n0_4741_5817  0.0191987 
iB01_223_v n1_4833_5864 0  0.0191987 
iB01_223_g 0 n0_4741_5850  0.0191987 
iB01_224_v n1_4833_6263 0  0.0191987 
iB01_224_g 0 n0_4741_6249  0.0191987 
iB01_225_v n1_4833_6296 0  0.0191987 
iB01_225_g 0 n0_4741_6282  0.0191987 
iB01_226_v n1_4833_6479 0  0.0191987 
iB01_226_g 0 n0_4741_6465  0.0191987 
iB01_227_v n1_4833_6512 0  0.0191987 
iB01_227_g 0 n0_4741_6498  0.0191987 
iB01_228_v n1_4833_6549 0  0.0191987 
iB01_228_g 0 n0_4741_6535  0.0191987 
iB01_229_v n1_4833_6646 0  0.0191987 
iB01_229_g 0 n0_4741_6681  0.0191987 
iB01_230_v n1_4833_6695 0  0.0191987 
iB01_230_g 0 n0_4741_6681  0.0191987 
iB01_231_v n1_4833_6728 0  0.0191987 
iB01_231_g 0 n0_4741_6714  0.0191987 
iB01_232_v n1_4833_6911 0  0.0191987 
iB01_232_g 0 n0_4741_6897  0.0191987 
iB01_233_v n1_4833_6944 0  0.0191987 
iB01_233_g 0 n0_4741_6930  0.0191987 
iB01_234_v n1_4833_7127 0  0.0191987 
iB01_234_g 0 n0_4741_7113  0.0191987 
iB01_235_v n1_4833_7160 0  0.0191987 
iB01_235_g 0 n0_4741_7146  0.0191987 
iB01_236_v n1_4880_7160 0  0.0191987 
iB01_236_g 0 n0_4929_7113  0.0191987 
iB01_237_v n1_4833_7343 0  0.0191987 
iB01_237_g 0 n0_4741_7329  0.0191987 
iB01_238_v n1_4833_7376 0  0.0191987 
iB01_238_g 0 n0_4741_7362  0.0191987 
iB01_239_v n1_4833_7559 0  0.0191987 
iB01_239_g 0 n0_4741_7545  0.0191987 
iB01_240_v n1_4833_7592 0  0.0191987 
iB01_240_g 0 n0_4741_7578  0.0191987 
iB01_241_v n1_4833_7775 0  0.0191987 
iB01_241_g 0 n0_4741_7761  0.0191987 
iB01_242_v n1_4833_7808 0  0.0191987 
iB01_242_g 0 n0_4741_7808  0.0191987 
iB01_243_v n1_4833_7822 0  0.0191987 
iB01_243_g 0 n0_4741_7808  0.0191987 
iB01_244_v n1_4833_7964 0  0.0191987 
iB01_244_g 0 n0_4741_7977  0.0191987 
iB01_245_v n1_4833_7991 0  0.0191987 
iB01_245_g 0 n0_4741_7977  0.0191987 
iB01_246_v n1_4833_8024 0  0.0191987 
iB01_246_g 0 n0_4741_8010  0.0191987 
iB01_247_v n1_4833_8207 0  0.0191987 
iB01_247_g 0 n0_4741_8193  0.0191987 
iB01_248_v n1_4833_8240 0  0.0191987 
iB01_248_g 0 n0_4741_8226  0.0191987 
iB01_249_v n1_4833_8456 0  0.0191987 
iB01_249_g 0 n0_4880_8409  0.0191987 
iB01_250_v n1_4833_8639 0  0.0191987 
iB01_250_g 0 n0_4741_8625  0.0191987 
iB01_251_v n1_4833_8672 0  0.0191987 
iB01_251_g 0 n0_4741_8658  0.0191987 
iB01_252_v n1_4833_8855 0  0.0191987 
iB01_252_g 0 n0_4741_8841  0.0191987 
iB01_253_v n1_4833_8888 0  0.0191987 
iB01_253_g 0 n0_4741_8888  0.0191987 
iB01_254_v n1_4833_8902 0  0.0191987 
iB01_254_g 0 n0_4741_8911  0.0191987 
iB01_255_v n1_4833_9022 0  0.0191987 
iB01_255_g 0 n0_4741_9057  0.0191987 
iB01_256_v n1_4833_9044 0  0.0191987 
iB01_256_g 0 n0_4741_9057  0.0191987 
iB01_257_v n1_4833_9071 0  0.0191987 
iB01_257_g 0 n0_4741_9057  0.0191987 
iB01_258_v n1_4833_9104 0  0.0191987 
iB01_258_g 0 n0_4741_9090  0.0191987 
iB01_259_v n1_4833_9287 0  0.0191987 
iB01_259_g 0 n0_4741_9273  0.0191987 
iB01_260_v n1_4833_9320 0  0.0191987 
iB01_260_g 0 n0_4741_9306  0.0191987 
iB01_261_v n1_4833_9503 0  0.0191987 
iB01_261_g 0 n0_4741_9489  0.0191987 
iB01_262_v n1_4833_9536 0  0.0191987 
iB01_262_g 0 n0_4741_9522  0.0191987 
iB01_263_v n1_4833_9719 0  0.0191987 
iB01_263_g 0 n0_4741_9705  0.0191987 
iB01_264_v n1_4833_9752 0  0.0191987 
iB01_264_g 0 n0_4741_9738  0.0191987 
iB01_265_v n1_4880_9503 0  0.0191987 
iB01_265_g 0 n0_4741_9489  0.0191987 
iB01_266_v n1_4880_9536 0  0.0191987 
iB01_266_g 0 n0_4741_9522  0.0191987 
iB01_267_v n1_4833_9935 0  0.0191987 
iB01_267_g 0 n0_4741_9921  0.0191987 
iB01_268_v n1_4833_9968 0  0.0191987 
iB01_268_g 0 n0_4741_9968  0.0191987 
iB01_269_v n1_4833_9982 0  0.0191987 
iB01_269_g 0 n0_4741_9968  0.0191987 
iB01_270_v n1_4833_10124 0  0.0191987 
iB01_270_g 0 n0_4741_10137  0.0191987 
iB01_271_v n1_4833_10151 0  0.0191987 
iB01_271_g 0 n0_4741_10137  0.0191987 
iB01_272_v n1_4833_10184 0  0.0191987 
iB01_272_g 0 n0_4741_10170  0.0191987 
iB01_273_v n1_4833_10367 0  0.0191987 
iB01_273_g 0 n0_4741_10353  0.0191987 
iB01_274_v n1_4833_10400 0  0.0191987 
iB01_274_g 0 n0_4741_10386  0.0191987 
iB01_275_v n1_5021_5399 0  0.0191987 
iB01_275_g 0 n0_4929_5385  0.0191987 
iB01_276_v n1_5021_5432 0  0.0191987 
iB01_276_g 0 n0_4929_5432  0.0191987 
iB01_277_v n1_5021_5446 0  0.0191987 
iB01_277_g 0 n0_4929_5432  0.0191987 
iB01_278_v n1_5021_5588 0  0.0191987 
iB01_278_g 0 n0_4929_5601  0.0191987 
iB01_279_v n1_5021_5615 0  0.0191987 
iB01_279_g 0 n0_4929_5601  0.0191987 
iB01_280_v n1_5021_5648 0  0.0191987 
iB01_280_g 0 n0_4929_5634  0.0191987 
iB01_281_v n1_5021_5831 0  0.0191987 
iB01_281_g 0 n0_4929_5817  0.0191987 
iB01_282_v n1_5021_5864 0  0.0191987 
iB01_282_g 0 n0_4929_5850  0.0191987 
iB01_283_v n1_5021_6047 0  0.0191987 
iB01_283_g 0 n0_4929_6033  0.0191987 
iB01_284_v n1_5021_6080 0  0.0191987 
iB01_284_g 0 n0_4929_6066  0.0191987 
iB01_285_v n1_5021_6263 0  0.0191987 
iB01_285_g 0 n0_4929_6249  0.0191987 
iB01_286_v n1_5021_6296 0  0.0191987 
iB01_286_g 0 n0_4929_6282  0.0191987 
iB01_287_v n1_5021_6479 0  0.0191987 
iB01_287_g 0 n0_4929_6465  0.0191987 
iB01_288_v n1_5021_6512 0  0.0191987 
iB01_288_g 0 n0_4929_6498  0.0191987 
iB01_289_v n1_5021_6549 0  0.0191987 
iB01_289_g 0 n0_4929_6535  0.0191987 
iB01_290_v n1_5021_6646 0  0.0191987 
iB01_290_g 0 n0_4929_6681  0.0191987 
iB01_291_v n1_5021_6695 0  0.0191987 
iB01_291_g 0 n0_4929_6681  0.0191987 
iB01_292_v n1_5021_6728 0  0.0191987 
iB01_292_g 0 n0_4929_6714  0.0191987 
iB01_293_v n1_5021_6911 0  0.0191987 
iB01_293_g 0 n0_4929_6897  0.0191987 
iB01_294_v n1_5021_6944 0  0.0191987 
iB01_294_g 0 n0_4929_6930  0.0191987 
iB01_295_v n1_5021_7127 0  0.0191987 
iB01_295_g 0 n0_4929_7113  0.0191987 
iB01_296_v n1_5021_7160 0  0.0191987 
iB01_296_g 0 n0_4929_7113  0.0191987 
iB01_297_v n1_5021_7343 0  0.0191987 
iB01_297_g 0 n0_4929_7329  0.0191987 
iB01_298_v n1_5021_7376 0  0.0191987 
iB01_298_g 0 n0_4929_7362  0.0191987 
iB01_299_v n1_5021_7559 0  0.0191987 
iB01_299_g 0 n0_4929_7545  0.0191987 
iB01_300_v n1_5021_7592 0  0.0191987 
iB01_300_g 0 n0_4929_7578  0.0191987 
iB01_301_v n1_5021_7775 0  0.0191987 
iB01_301_g 0 n0_4929_7761  0.0191987 
iB01_302_v n1_5021_7808 0  0.0191987 
iB01_302_g 0 n0_4929_7808  0.0191987 
iB01_303_v n1_5021_7822 0  0.0191987 
iB01_303_g 0 n0_4929_7808  0.0191987 
iB01_304_v n1_5021_7964 0  0.0191987 
iB01_304_g 0 n0_4929_7977  0.0191987 
iB01_305_v n1_5021_7991 0  0.0191987 
iB01_305_g 0 n0_4929_7977  0.0191987 
iB01_306_v n1_5021_8024 0  0.0191987 
iB01_306_g 0 n0_4929_8010  0.0191987 
iB01_307_v n1_5021_8207 0  0.0191987 
iB01_307_g 0 n0_4929_8193  0.0191987 
iB01_308_v n1_5021_8240 0  0.0191987 
iB01_308_g 0 n0_4929_8226  0.0191987 
iB01_309_v n1_5021_8423 0  0.0191987 
iB01_309_g 0 n0_4929_8409  0.0191987 
iB01_310_v n1_5021_8456 0  0.0191987 
iB01_310_g 0 n0_4929_8442  0.0191987 
iB01_311_v n1_5021_8639 0  0.0191987 
iB01_311_g 0 n0_4929_8625  0.0191987 
iB01_312_v n1_5021_8672 0  0.0191987 
iB01_312_g 0 n0_4929_8658  0.0191987 
iB01_313_v n1_5021_8855 0  0.0191987 
iB01_313_g 0 n0_4929_8841  0.0191987 
iB01_314_v n1_5021_8888 0  0.0191987 
iB01_314_g 0 n0_4929_8888  0.0191987 
iB01_315_v n1_5021_8902 0  0.0191987 
iB01_315_g 0 n0_4929_8911  0.0191987 
iB01_316_v n1_5021_9022 0  0.0191987 
iB01_316_g 0 n0_4929_9057  0.0191987 
iB01_317_v n1_5021_9044 0  0.0191987 
iB01_317_g 0 n0_4929_9057  0.0191987 
iB01_318_v n1_5021_9071 0  0.0191987 
iB01_318_g 0 n0_4929_9057  0.0191987 
iB01_319_v n1_5021_9104 0  0.0191987 
iB01_319_g 0 n0_4929_9090  0.0191987 
iB01_320_v n1_5021_9287 0  0.0191987 
iB01_320_g 0 n0_4929_9273  0.0191987 
iB01_321_v n1_5021_9320 0  0.0191987 
iB01_321_g 0 n0_4929_9306  0.0191987 
iB01_322_v n1_5021_9503 0  0.0191987 
iB01_322_g 0 n0_4929_9306  0.0191987 
iB01_323_v n1_5021_9536 0  0.0191987 
iB01_323_g 0 n0_4929_9705  0.0191987 
iB01_324_v n1_5021_9719 0  0.0191987 
iB01_324_g 0 n0_4929_9705  0.0191987 
iB01_325_v n1_5021_9752 0  0.0191987 
iB01_325_g 0 n0_4929_9738  0.0191987 
iB01_326_v n1_5021_9935 0  0.0191987 
iB01_326_g 0 n0_4929_9921  0.0191987 
iB01_327_v n1_5021_9968 0  0.0191987 
iB01_327_g 0 n0_4929_9968  0.0191987 
iB01_328_v n1_5021_9982 0  0.0191987 
iB01_328_g 0 n0_4929_9968  0.0191987 
iB01_329_v n1_5021_10124 0  0.0191987 
iB01_329_g 0 n0_4929_10137  0.0191987 
iB01_330_v n1_5021_10151 0  0.0191987 
iB01_330_g 0 n0_4929_10137  0.0191987 
iB01_331_v n1_5021_10184 0  0.0191987 
iB01_331_g 0 n0_4929_10170  0.0191987 
iB01_332_v n1_5021_10367 0  0.0191987 
iB01_332_g 0 n0_4929_10353  0.0191987 
iB01_333_v n1_5021_10400 0  0.0191987 
iB01_333_g 0 n0_4929_10386  0.0191987 
iB01_334_v n1_5021_10616 0  0.0191987 
iB01_334_g 0 n0_4929_10602  0.0191987 
iB02_0_v n1_333_10799 0  0.0191328 
iB02_0_g 0 n0_241_10785  0.0191328 
iB02_1_v n1_333_10832 0  0.0191328 
iB02_1_g 0 n0_241_10818  0.0191328 
iB02_2_v n1_521_10799 0  0.0191328 
iB02_2_g 0 n0_429_10785  0.0191328 
iB02_3_v n1_521_10832 0  0.0191328 
iB02_3_g 0 n0_429_10818  0.0191328 
iB02_4_v n1_333_11015 0  0.0191328 
iB02_4_g 0 n0_241_11001  0.0191328 
iB02_5_v n1_333_11048 0  0.0191328 
iB02_5_g 0 n0_241_11034  0.0191328 
iB02_6_v n1_333_11231 0  0.0191328 
iB02_6_g 0 n0_241_11217  0.0191328 
iB02_7_v n1_333_11264 0  0.0191328 
iB02_7_g 0 n0_241_11250  0.0191328 
iB02_8_v n1_521_11015 0  0.0191328 
iB02_8_g 0 n0_429_11001  0.0191328 
iB02_9_v n1_521_11048 0  0.0191328 
iB02_9_g 0 n0_429_11034  0.0191328 
iB02_10_v n1_521_11231 0  0.0191328 
iB02_10_g 0 n0_429_11217  0.0191328 
iB02_11_v n1_521_11264 0  0.0191328 
iB02_11_g 0 n0_429_11250  0.0191328 
iB02_12_v n1_333_11447 0  0.0191328 
iB02_12_g 0 n0_241_11433  0.0191328 
iB02_13_v n1_333_11480 0  0.0191328 
iB02_13_g 0 n0_241_11466  0.0191328 
iB02_14_v n1_333_11663 0  0.0191328 
iB02_14_g 0 n0_241_11649  0.0191328 
iB02_15_v n1_333_11696 0  0.0191328 
iB02_15_g 0 n0_241_11682  0.0191328 
iB02_16_v n1_380_11663 0  0.0191328 
iB02_16_g 0 n0_241_11649  0.0191328 
iB02_17_v n1_380_11696 0  0.0191328 
iB02_17_g 0 n0_241_11682  0.0191328 
iB02_18_v n1_521_11447 0  0.0191328 
iB02_18_g 0 n0_429_11433  0.0191328 
iB02_19_v n1_521_11480 0  0.0191328 
iB02_19_g 0 n0_429_11466  0.0191328 
iB02_20_v n1_521_11663 0  0.0191328 
iB02_20_g 0 n0_429_11466  0.0191328 
iB02_21_v n1_521_11696 0  0.0191328 
iB02_21_g 0 n0_429_11865  0.0191328 
iB02_22_v n1_333_11879 0  0.0191328 
iB02_22_g 0 n0_241_11865  0.0191328 
iB02_23_v n1_333_11912 0  0.0191328 
iB02_23_g 0 n0_241_11898  0.0191328 
iB02_24_v n1_333_12095 0  0.0191328 
iB02_24_g 0 n0_241_12081  0.0191328 
iB02_25_v n1_333_12128 0  0.0191328 
iB02_25_g 0 n0_241_12114  0.0191328 
iB02_26_v n1_521_11879 0  0.0191328 
iB02_26_g 0 n0_429_11865  0.0191328 
iB02_27_v n1_521_11912 0  0.0191328 
iB02_27_g 0 n0_429_11898  0.0191328 
iB02_28_v n1_521_12095 0  0.0191328 
iB02_28_g 0 n0_429_12081  0.0191328 
iB02_29_v n1_521_12128 0  0.0191328 
iB02_29_g 0 n0_429_12114  0.0191328 
iB02_30_v n1_333_12311 0  0.0191328 
iB02_30_g 0 n0_241_12297  0.0191328 
iB02_31_v n1_333_12344 0  0.0191328 
iB02_31_g 0 n0_241_12330  0.0191328 
iB02_32_v n1_333_12527 0  0.0191328 
iB02_32_g 0 n0_241_12513  0.0191328 
iB02_33_v n1_333_12560 0  0.0191328 
iB02_33_g 0 n0_241_12546  0.0191328 
iB02_34_v n1_521_12311 0  0.0191328 
iB02_34_g 0 n0_429_12297  0.0191328 
iB02_35_v n1_521_12344 0  0.0191328 
iB02_35_g 0 n0_429_12330  0.0191328 
iB02_36_v n1_521_12527 0  0.0191328 
iB02_36_g 0 n0_429_12513  0.0191328 
iB02_37_v n1_521_12560 0  0.0191328 
iB02_37_g 0 n0_429_12546  0.0191328 
iB02_38_v n1_333_12743 0  0.0191328 
iB02_38_g 0 n0_241_12729  0.0191328 
iB02_39_v n1_333_12959 0  0.0191328 
iB02_39_g 0 n0_241_12945  0.0191328 
iB02_40_v n1_333_12992 0  0.0191328 
iB02_40_g 0 n0_241_12978  0.0191328 
iB02_41_v n1_521_12743 0  0.0191328 
iB02_41_g 0 n0_429_12729  0.0191328 
iB02_42_v n1_521_12776 0  0.0191328 
iB02_42_g 0 n0_429_12762  0.0191328 
iB02_43_v n1_521_12959 0  0.0191328 
iB02_43_g 0 n0_429_12945  0.0191328 
iB02_44_v n1_521_12992 0  0.0191328 
iB02_44_g 0 n0_429_12978  0.0191328 
iB02_45_v n1_333_13175 0  0.0191328 
iB02_45_g 0 n0_241_13161  0.0191328 
iB02_46_v n1_333_13208 0  0.0191328 
iB02_46_g 0 n0_241_13194  0.0191328 
iB02_47_v n1_333_13391 0  0.0191328 
iB02_47_g 0 n0_241_13377  0.0191328 
iB02_48_v n1_333_13424 0  0.0191328 
iB02_48_g 0 n0_241_13410  0.0191328 
iB02_49_v n1_521_13175 0  0.0191328 
iB02_49_g 0 n0_429_13161  0.0191328 
iB02_50_v n1_521_13208 0  0.0191328 
iB02_50_g 0 n0_429_13194  0.0191328 
iB02_51_v n1_521_13391 0  0.0191328 
iB02_51_g 0 n0_429_13377  0.0191328 
iB02_52_v n1_521_13424 0  0.0191328 
iB02_52_g 0 n0_429_13410  0.0191328 
iB02_53_v n1_333_13607 0  0.0191328 
iB02_53_g 0 n0_241_13593  0.0191328 
iB02_54_v n1_333_13640 0  0.0191328 
iB02_54_g 0 n0_241_13626  0.0191328 
iB02_55_v n1_333_13774 0  0.0191328 
iB02_55_g 0 n0_241_13809  0.0191328 
iB02_56_v n1_333_13823 0  0.0191328 
iB02_56_g 0 n0_241_13809  0.0191328 
iB02_57_v n1_333_13856 0  0.0191328 
iB02_57_g 0 n0_241_13842  0.0191328 
iB02_58_v n1_521_13607 0  0.0191328 
iB02_58_g 0 n0_429_13593  0.0191328 
iB02_59_v n1_521_13640 0  0.0191328 
iB02_59_g 0 n0_429_13626  0.0191328 
iB02_60_v n1_521_13774 0  0.0191328 
iB02_60_g 0 n0_429_13809  0.0191328 
iB02_61_v n1_521_13823 0  0.0191328 
iB02_61_g 0 n0_429_13809  0.0191328 
iB02_62_v n1_521_13856 0  0.0191328 
iB02_62_g 0 n0_429_13842  0.0191328 
iB02_63_v n1_333_14039 0  0.0191328 
iB02_63_g 0 n0_241_14025  0.0191328 
iB02_64_v n1_333_14072 0  0.0191328 
iB02_64_g 0 n0_241_14058  0.0191328 
iB02_65_v n1_333_14255 0  0.0191328 
iB02_65_g 0 n0_241_14241  0.0191328 
iB02_66_v n1_380_14039 0  0.0191328 
iB02_66_g 0 n0_241_14025  0.0191328 
iB02_67_v n1_521_14039 0  0.0191328 
iB02_67_g 0 n0_429_13842  0.0191328 
iB02_68_v n1_521_14072 0  0.0191328 
iB02_68_g 0 n0_429_14241  0.0191328 
iB02_69_v n1_521_14255 0  0.0191328 
iB02_69_g 0 n0_429_14241  0.0191328 
iB02_70_v n1_333_14288 0  0.0191328 
iB02_70_g 0 n0_241_14274  0.0191328 
iB02_71_v n1_333_14471 0  0.0191328 
iB02_71_g 0 n0_241_14457  0.0191328 
iB02_72_v n1_333_14504 0  0.0191328 
iB02_72_g 0 n0_241_14490  0.0191328 
iB02_73_v n1_521_14288 0  0.0191328 
iB02_73_g 0 n0_429_14274  0.0191328 
iB02_74_v n1_521_14471 0  0.0191328 
iB02_74_g 0 n0_429_14457  0.0191328 
iB02_75_v n1_521_14504 0  0.0191328 
iB02_75_g 0 n0_429_14490  0.0191328 
iB02_76_v n1_333_14687 0  0.0191328 
iB02_76_g 0 n0_241_14673  0.0191328 
iB02_77_v n1_333_14720 0  0.0191328 
iB02_77_g 0 n0_241_14706  0.0191328 
iB02_78_v n1_333_14903 0  0.0191328 
iB02_78_g 0 n0_241_14889  0.0191328 
iB02_79_v n1_333_14936 0  0.0191328 
iB02_79_g 0 n0_241_14922  0.0191328 
iB02_80_v n1_521_14687 0  0.0191328 
iB02_80_g 0 n0_429_14673  0.0191328 
iB02_81_v n1_521_14720 0  0.0191328 
iB02_81_g 0 n0_429_14706  0.0191328 
iB02_82_v n1_521_14903 0  0.0191328 
iB02_82_g 0 n0_429_14889  0.0191328 
iB02_83_v n1_521_14936 0  0.0191328 
iB02_83_g 0 n0_429_14922  0.0191328 
iB02_84_v n1_333_15335 0  0.0191328 
iB02_84_g 0 n0_241_15321  0.0191328 
iB02_85_v n1_333_15368 0  0.0191328 
iB02_85_g 0 n0_241_15354  0.0191328 
iB02_86_v n1_521_15119 0  0.0191328 
iB02_86_g 0 n0_429_15105  0.0191328 
iB02_87_v n1_521_15152 0  0.0191328 
iB02_87_g 0 n0_429_15138  0.0191328 
iB02_88_v n1_521_15335 0  0.0191328 
iB02_88_g 0 n0_429_15321  0.0191328 
iB02_89_v n1_521_15368 0  0.0191328 
iB02_89_g 0 n0_429_15354  0.0191328 
iB02_90_v n1_333_15551 0  0.0191328 
iB02_90_g 0 n0_241_15537  0.0191328 
iB02_91_v n1_333_15584 0  0.0191328 
iB02_91_g 0 n0_241_15570  0.0191328 
iB02_92_v n1_333_15767 0  0.0191328 
iB02_92_g 0 n0_241_15753  0.0191328 
iB02_93_v n1_333_15800 0  0.0191328 
iB02_93_g 0 n0_241_15786  0.0191328 
iB02_94_v n1_521_15551 0  0.0191328 
iB02_94_g 0 n0_429_15537  0.0191328 
iB02_95_v n1_521_15584 0  0.0191328 
iB02_95_g 0 n0_429_15570  0.0191328 
iB02_96_v n1_521_15767 0  0.0191328 
iB02_96_g 0 n0_429_15753  0.0191328 
iB02_97_v n1_521_15800 0  0.0191328 
iB02_97_g 0 n0_429_15786  0.0191328 
iB02_98_v n1_2583_10799 0  0.0191328 
iB02_98_g 0 n0_2491_10785  0.0191328 
iB02_99_v n1_2583_10832 0  0.0191328 
iB02_99_g 0 n0_2491_10818  0.0191328 
iB02_100_v n1_2771_10799 0  0.0191328 
iB02_100_g 0 n0_2679_10785  0.0191328 
iB02_101_v n1_2771_10832 0  0.0191328 
iB02_101_g 0 n0_2679_10818  0.0191328 
iB02_102_v n1_2583_11015 0  0.0191328 
iB02_102_g 0 n0_2491_11001  0.0191328 
iB02_103_v n1_2583_11048 0  0.0191328 
iB02_103_g 0 n0_2491_11048  0.0191328 
iB02_104_v n1_2583_11182 0  0.0191328 
iB02_104_g 0 n0_2491_11217  0.0191328 
iB02_105_v n1_2583_11204 0  0.0191328 
iB02_105_g 0 n0_2491_11217  0.0191328 
iB02_106_v n1_2583_11231 0  0.0191328 
iB02_106_g 0 n0_2491_11217  0.0191328 
iB02_107_v n1_2583_11264 0  0.0191328 
iB02_107_g 0 n0_2491_11250  0.0191328 
iB02_108_v n1_2771_11015 0  0.0191328 
iB02_108_g 0 n0_2679_11001  0.0191328 
iB02_109_v n1_2771_11048 0  0.0191328 
iB02_109_g 0 n0_2679_11048  0.0191328 
iB02_110_v n1_2771_11182 0  0.0191328 
iB02_110_g 0 n0_2679_11217  0.0191328 
iB02_111_v n1_2771_11204 0  0.0191328 
iB02_111_g 0 n0_2679_11217  0.0191328 
iB02_112_v n1_2771_11231 0  0.0191328 
iB02_112_g 0 n0_2679_11217  0.0191328 
iB02_113_v n1_2771_11264 0  0.0191328 
iB02_113_g 0 n0_2679_11250  0.0191328 
iB02_114_v n1_2583_11447 0  0.0191328 
iB02_114_g 0 n0_2491_11433  0.0191328 
iB02_115_v n1_2583_11480 0  0.0191328 
iB02_115_g 0 n0_2491_11466  0.0191328 
iB02_116_v n1_2583_11663 0  0.0191328 
iB02_116_g 0 n0_2491_11649  0.0191328 
iB02_117_v n1_2583_11696 0  0.0191328 
iB02_117_g 0 n0_2491_11682  0.0191328 
iB02_118_v n1_2630_11663 0  0.0191328 
iB02_118_g 0 n0_2491_11649  0.0191328 
iB02_119_v n1_2630_11696 0  0.0191328 
iB02_119_g 0 n0_2491_11682  0.0191328 
iB02_120_v n1_2771_11447 0  0.0191328 
iB02_120_g 0 n0_2679_11433  0.0191328 
iB02_121_v n1_2771_11480 0  0.0191328 
iB02_121_g 0 n0_2679_11466  0.0191328 
iB02_122_v n1_2771_11663 0  0.0191328 
iB02_122_g 0 n0_2679_11466  0.0191328 
iB02_123_v n1_2771_11696 0  0.0191328 
iB02_123_g 0 n0_2679_11865  0.0191328 
iB02_124_v n1_2583_11879 0  0.0191328 
iB02_124_g 0 n0_2491_11865  0.0191328 
iB02_125_v n1_2583_11912 0  0.0191328 
iB02_125_g 0 n0_2491_11898  0.0191328 
iB02_126_v n1_2583_12095 0  0.0191328 
iB02_126_g 0 n0_2491_12081  0.0191328 
iB02_127_v n1_2583_12128 0  0.0191328 
iB02_127_g 0 n0_2491_12128  0.0191328 
iB02_128_v n1_2771_11879 0  0.0191328 
iB02_128_g 0 n0_2679_11865  0.0191328 
iB02_129_v n1_2771_11912 0  0.0191328 
iB02_129_g 0 n0_2679_11898  0.0191328 
iB02_130_v n1_2771_12095 0  0.0191328 
iB02_130_g 0 n0_2679_12081  0.0191328 
iB02_131_v n1_2771_12128 0  0.0191328 
iB02_131_g 0 n0_2679_12128  0.0191328 
iB02_132_v n1_2583_12262 0  0.0191328 
iB02_132_g 0 n0_2491_12297  0.0191328 
iB02_133_v n1_2583_12284 0  0.0191328 
iB02_133_g 0 n0_2491_12297  0.0191328 
iB02_134_v n1_2583_12311 0  0.0191328 
iB02_134_g 0 n0_2491_12297  0.0191328 
iB02_135_v n1_2583_12344 0  0.0191328 
iB02_135_g 0 n0_2491_12330  0.0191328 
iB02_136_v n1_2583_12527 0  0.0191328 
iB02_136_g 0 n0_2491_12513  0.0191328 
iB02_137_v n1_2583_12560 0  0.0191328 
iB02_137_g 0 n0_2491_12546  0.0191328 
iB02_138_v n1_2771_12262 0  0.0191328 
iB02_138_g 0 n0_2679_12297  0.0191328 
iB02_139_v n1_2771_12284 0  0.0191328 
iB02_139_g 0 n0_2679_12297  0.0191328 
iB02_140_v n1_2771_12311 0  0.0191328 
iB02_140_g 0 n0_2679_12297  0.0191328 
iB02_141_v n1_2771_12344 0  0.0191328 
iB02_141_g 0 n0_2679_12330  0.0191328 
iB02_142_v n1_2771_12527 0  0.0191328 
iB02_142_g 0 n0_2679_12513  0.0191328 
iB02_143_v n1_2771_12560 0  0.0191328 
iB02_143_g 0 n0_2679_12546  0.0191328 
iB02_144_v n1_2583_12743 0  0.0191328 
iB02_144_g 0 n0_2491_12729  0.0191328 
iB02_145_v n1_2583_12959 0  0.0191328 
iB02_145_g 0 n0_2491_12945  0.0191328 
iB02_146_v n1_2583_12992 0  0.0191328 
iB02_146_g 0 n0_2491_12978  0.0191328 
iB02_147_v n1_2771_12743 0  0.0191328 
iB02_147_g 0 n0_2679_12729  0.0191328 
iB02_148_v n1_2771_12776 0  0.0191328 
iB02_148_g 0 n0_2679_12762  0.0191328 
iB02_149_v n1_2771_12959 0  0.0191328 
iB02_149_g 0 n0_2679_12945  0.0191328 
iB02_150_v n1_2771_12992 0  0.0191328 
iB02_150_g 0 n0_2679_12978  0.0191328 
iB02_151_v n1_2583_13175 0  0.0191328 
iB02_151_g 0 n0_2491_13161  0.0191328 
iB02_152_v n1_2583_13208 0  0.0191328 
iB02_152_g 0 n0_2491_13194  0.0191328 
iB02_153_v n1_2583_13391 0  0.0191328 
iB02_153_g 0 n0_2491_13377  0.0191328 
iB02_154_v n1_2583_13424 0  0.0191328 
iB02_154_g 0 n0_2491_13424  0.0191328 
iB02_155_v n1_2771_13175 0  0.0191328 
iB02_155_g 0 n0_2679_13161  0.0191328 
iB02_156_v n1_2771_13208 0  0.0191328 
iB02_156_g 0 n0_2679_13194  0.0191328 
iB02_157_v n1_2771_13391 0  0.0191328 
iB02_157_g 0 n0_2679_13377  0.0191328 
iB02_158_v n1_2771_13424 0  0.0191328 
iB02_158_g 0 n0_2679_13424  0.0191328 
iB02_159_v n1_2583_13558 0  0.0191328 
iB02_159_g 0 n0_2491_13593  0.0191328 
iB02_160_v n1_2583_13580 0  0.0191328 
iB02_160_g 0 n0_2491_13593  0.0191328 
iB02_161_v n1_2583_13607 0  0.0191328 
iB02_161_g 0 n0_2491_13593  0.0191328 
iB02_162_v n1_2583_13640 0  0.0191328 
iB02_162_g 0 n0_2491_13640  0.0191328 
iB02_163_v n1_2583_13796 0  0.0191328 
iB02_163_g 0 n0_2491_13809  0.0191328 
iB02_164_v n1_2583_13823 0  0.0191328 
iB02_164_g 0 n0_2491_13809  0.0191328 
iB02_165_v n1_2583_13856 0  0.0191328 
iB02_165_g 0 n0_2491_13842  0.0191328 
iB02_166_v n1_2771_13558 0  0.0191328 
iB02_166_g 0 n0_2679_13593  0.0191328 
iB02_167_v n1_2771_13580 0  0.0191328 
iB02_167_g 0 n0_2679_13593  0.0191328 
iB02_168_v n1_2771_13607 0  0.0191328 
iB02_168_g 0 n0_2679_13593  0.0191328 
iB02_169_v n1_2771_13640 0  0.0191328 
iB02_169_g 0 n0_2679_13640  0.0191328 
iB02_170_v n1_2771_13796 0  0.0191328 
iB02_170_g 0 n0_2679_13809  0.0191328 
iB02_171_v n1_2771_13823 0  0.0191328 
iB02_171_g 0 n0_2679_13809  0.0191328 
iB02_172_v n1_2771_13856 0  0.0191328 
iB02_172_g 0 n0_2679_13842  0.0191328 
iB02_173_v n1_2583_13990 0  0.0191328 
iB02_173_g 0 n0_2491_14025  0.0191328 
iB02_174_v n1_2583_14039 0  0.0191328 
iB02_174_g 0 n0_2491_14025  0.0191328 
iB02_175_v n1_2583_14072 0  0.0191328 
iB02_175_g 0 n0_2491_14058  0.0191328 
iB02_176_v n1_2583_14206 0  0.0191328 
iB02_176_g 0 n0_2491_14241  0.0191328 
iB02_177_v n1_2583_14255 0  0.0191328 
iB02_177_g 0 n0_2491_14241  0.0191328 
iB02_178_v n1_2630_13990 0  0.0191328 
iB02_178_g 0 n0_2679_14100  0.0191328 
iB02_179_v n1_2630_14039 0  0.0191328 
iB02_179_g 0 n0_2679_14100  0.0191328 
iB02_180_v n1_2771_13990 0  0.0191328 
iB02_180_g 0 n0_2679_14100  0.0191328 
iB02_181_v n1_2771_14039 0  0.0191328 
iB02_181_g 0 n0_2679_14100  0.0191328 
iB02_182_v n1_2771_14072 0  0.0191328 
iB02_182_g 0 n0_2679_14100  0.0191328 
iB02_183_v n1_2771_14206 0  0.0191328 
iB02_183_g 0 n0_2679_14241  0.0191328 
iB02_184_v n1_2771_14255 0  0.0191328 
iB02_184_g 0 n0_2679_14241  0.0191328 
iB02_185_v n1_2583_14288 0  0.0191328 
iB02_185_g 0 n0_2491_14274  0.0191328 
iB02_186_v n1_2583_14471 0  0.0191328 
iB02_186_g 0 n0_2491_14457  0.0191328 
iB02_187_v n1_2583_14504 0  0.0191328 
iB02_187_g 0 n0_2491_14504  0.0191328 
iB02_188_v n1_2583_14660 0  0.0191328 
iB02_188_g 0 n0_2491_14673  0.0191328 
iB02_189_v n1_2771_14288 0  0.0191328 
iB02_189_g 0 n0_2679_14274  0.0191328 
iB02_190_v n1_2771_14471 0  0.0191328 
iB02_190_g 0 n0_2679_14457  0.0191328 
iB02_191_v n1_2771_14504 0  0.0191328 
iB02_191_g 0 n0_2679_14504  0.0191328 
iB02_192_v n1_2771_14660 0  0.0191328 
iB02_192_g 0 n0_2679_14673  0.0191328 
iB02_193_v n1_2583_14687 0  0.0191328 
iB02_193_g 0 n0_2491_14673  0.0191328 
iB02_194_v n1_2583_14720 0  0.0191328 
iB02_194_g 0 n0_2491_14706  0.0191328 
iB02_195_v n1_2583_14903 0  0.0191328 
iB02_195_g 0 n0_2491_14889  0.0191328 
iB02_196_v n1_2583_14936 0  0.0191328 
iB02_196_g 0 n0_2491_14922  0.0191328 
iB02_197_v n1_2771_14687 0  0.0191328 
iB02_197_g 0 n0_2679_14673  0.0191328 
iB02_198_v n1_2771_14720 0  0.0191328 
iB02_198_g 0 n0_2679_14706  0.0191328 
iB02_199_v n1_2771_14903 0  0.0191328 
iB02_199_g 0 n0_2679_14889  0.0191328 
iB02_200_v n1_2771_14936 0  0.0191328 
iB02_200_g 0 n0_2679_14922  0.0191328 
iB02_201_v n1_2583_15335 0  0.0191328 
iB02_201_g 0 n0_2491_15321  0.0191328 
iB02_202_v n1_2583_15368 0  0.0191328 
iB02_202_g 0 n0_2491_15368  0.0191328 
iB02_203_v n1_2771_15119 0  0.0191328 
iB02_203_g 0 n0_2679_15105  0.0191328 
iB02_204_v n1_2771_15152 0  0.0191328 
iB02_204_g 0 n0_2679_15138  0.0191328 
iB02_205_v n1_2771_15335 0  0.0191328 
iB02_205_g 0 n0_2679_15321  0.0191328 
iB02_206_v n1_2771_15368 0  0.0191328 
iB02_206_g 0 n0_2679_15368  0.0191328 
iB02_207_v n1_2583_15524 0  0.0191328 
iB02_207_g 0 n0_2491_15537  0.0191328 
iB02_208_v n1_2583_15551 0  0.0191328 
iB02_208_g 0 n0_2491_15537  0.0191328 
iB02_209_v n1_2583_15584 0  0.0191328 
iB02_209_g 0 n0_2491_15584  0.0191328 
iB02_210_v n1_2583_15740 0  0.0191328 
iB02_210_g 0 n0_2491_15753  0.0191328 
iB02_211_v n1_2583_15767 0  0.0191328 
iB02_211_g 0 n0_2491_15753  0.0191328 
iB02_212_v n1_2583_15800 0  0.0191328 
iB02_212_g 0 n0_2491_15786  0.0191328 
iB02_213_v n1_2771_15524 0  0.0191328 
iB02_213_g 0 n0_2679_15537  0.0191328 
iB02_214_v n1_2771_15551 0  0.0191328 
iB02_214_g 0 n0_2679_15537  0.0191328 
iB02_215_v n1_2771_15584 0  0.0191328 
iB02_215_g 0 n0_2679_15584  0.0191328 
iB02_216_v n1_2771_15740 0  0.0191328 
iB02_216_g 0 n0_2679_15753  0.0191328 
iB02_217_v n1_2771_15767 0  0.0191328 
iB02_217_g 0 n0_2679_15753  0.0191328 
iB02_218_v n1_2771_15800 0  0.0191328 
iB02_218_g 0 n0_2679_15786  0.0191328 
iB02_219_v n1_4833_10799 0  0.0191328 
iB02_219_g 0 n0_4741_10785  0.0191328 
iB02_220_v n1_4833_10832 0  0.0191328 
iB02_220_g 0 n0_4741_10818  0.0191328 
iB02_221_v n1_4833_11015 0  0.0191328 
iB02_221_g 0 n0_4741_11001  0.0191328 
iB02_222_v n1_4833_11048 0  0.0191328 
iB02_222_g 0 n0_4741_11048  0.0191328 
iB02_223_v n1_4833_11182 0  0.0191328 
iB02_223_g 0 n0_4741_11217  0.0191328 
iB02_224_v n1_4833_11204 0  0.0191328 
iB02_224_g 0 n0_4741_11217  0.0191328 
iB02_225_v n1_4833_11231 0  0.0191328 
iB02_225_g 0 n0_4741_11217  0.0191328 
iB02_226_v n1_4833_11264 0  0.0191328 
iB02_226_g 0 n0_4741_11250  0.0191328 
iB02_227_v n1_4833_11447 0  0.0191328 
iB02_227_g 0 n0_4741_11433  0.0191328 
iB02_228_v n1_4833_11480 0  0.0191328 
iB02_228_g 0 n0_4741_11466  0.0191328 
iB02_229_v n1_4833_11663 0  0.0191328 
iB02_229_g 0 n0_4741_11649  0.0191328 
iB02_230_v n1_4833_11696 0  0.0191328 
iB02_230_g 0 n0_4741_11682  0.0191328 
iB02_231_v n1_4880_11663 0  0.0191328 
iB02_231_g 0 n0_4741_11649  0.0191328 
iB02_232_v n1_4880_11696 0  0.0191328 
iB02_232_g 0 n0_4741_11682  0.0191328 
iB02_233_v n1_4833_11879 0  0.0191328 
iB02_233_g 0 n0_4741_11865  0.0191328 
iB02_234_v n1_4833_11912 0  0.0191328 
iB02_234_g 0 n0_4741_11898  0.0191328 
iB02_235_v n1_4833_12095 0  0.0191328 
iB02_235_g 0 n0_4741_12081  0.0191328 
iB02_236_v n1_4833_12128 0  0.0191328 
iB02_236_g 0 n0_4741_12128  0.0191328 
iB02_237_v n1_4833_12284 0  0.0191328 
iB02_237_g 0 n0_4741_12297  0.0191328 
iB02_238_v n1_4833_12311 0  0.0191328 
iB02_238_g 0 n0_4741_12297  0.0191328 
iB02_239_v n1_4833_12344 0  0.0191328 
iB02_239_g 0 n0_4741_12330  0.0191328 
iB02_240_v n1_4833_12527 0  0.0191328 
iB02_240_g 0 n0_4741_12513  0.0191328 
iB02_241_v n1_4833_12560 0  0.0191328 
iB02_241_g 0 n0_4741_12546  0.0191328 
iB02_242_v n1_4833_12743 0  0.0191328 
iB02_242_g 0 n0_4741_12729  0.0191328 
iB02_243_v n1_4833_12959 0  0.0191328 
iB02_243_g 0 n0_4741_12945  0.0191328 
iB02_244_v n1_4833_12992 0  0.0191328 
iB02_244_g 0 n0_4741_12978  0.0191328 
iB02_245_v n1_4833_13175 0  0.0191328 
iB02_245_g 0 n0_4741_13161  0.0191328 
iB02_246_v n1_4833_13208 0  0.0191328 
iB02_246_g 0 n0_4741_13194  0.0191328 
iB02_247_v n1_4833_13391 0  0.0191328 
iB02_247_g 0 n0_4741_13377  0.0191328 
iB02_248_v n1_4833_13424 0  0.0191328 
iB02_248_g 0 n0_4741_13424  0.0191328 
iB02_249_v n1_4833_13580 0  0.0191328 
iB02_249_g 0 n0_4741_13593  0.0191328 
iB02_250_v n1_4833_13607 0  0.0191328 
iB02_250_g 0 n0_4741_13593  0.0191328 
iB02_251_v n1_4833_13640 0  0.0191328 
iB02_251_g 0 n0_4741_13626  0.0191328 
iB02_252_v n1_4833_13823 0  0.0191328 
iB02_252_g 0 n0_4741_13809  0.0191328 
iB02_253_v n1_4833_13856 0  0.0191328 
iB02_253_g 0 n0_4741_13842  0.0191328 
iB02_254_v n1_4833_13990 0  0.0191328 
iB02_254_g 0 n0_4741_14025  0.0191328 
iB02_255_v n1_4833_14039 0  0.0191328 
iB02_255_g 0 n0_4741_14025  0.0191328 
iB02_256_v n1_4833_14072 0  0.0191328 
iB02_256_g 0 n0_4741_14058  0.0191328 
iB02_257_v n1_4833_14206 0  0.0191328 
iB02_257_g 0 n0_4741_14241  0.0191328 
iB02_258_v n1_4833_14255 0  0.0191328 
iB02_258_g 0 n0_4741_14241  0.0191328 
iB02_259_v n1_4880_13990 0  0.0191328 
iB02_259_g 0 n0_4929_14100  0.0191328 
iB02_260_v n1_4880_14039 0  0.0191328 
iB02_260_g 0 n0_4929_14100  0.0191328 
iB02_261_v n1_4833_14288 0  0.0191328 
iB02_261_g 0 n0_4741_14274  0.0191328 
iB02_262_v n1_4833_14471 0  0.0191328 
iB02_262_g 0 n0_4741_14457  0.0191328 
iB02_263_v n1_4833_14504 0  0.0191328 
iB02_263_g 0 n0_4741_14490  0.0191328 
iB02_264_v n1_4833_14687 0  0.0191328 
iB02_264_g 0 n0_4741_14673  0.0191328 
iB02_265_v n1_4833_14720 0  0.0191328 
iB02_265_g 0 n0_4741_14706  0.0191328 
iB02_266_v n1_4833_14903 0  0.0191328 
iB02_266_g 0 n0_4741_14889  0.0191328 
iB02_267_v n1_4833_14936 0  0.0191328 
iB02_267_g 0 n0_4741_14922  0.0191328 
iB02_268_v n1_4833_15335 0  0.0191328 
iB02_268_g 0 n0_4741_15321  0.0191328 
iB02_269_v n1_4833_15368 0  0.0191328 
iB02_269_g 0 n0_4741_15368  0.0191328 
iB02_270_v n1_4833_15524 0  0.0191328 
iB02_270_g 0 n0_4741_15537  0.0191328 
iB02_271_v n1_4833_15551 0  0.0191328 
iB02_271_g 0 n0_4741_15537  0.0191328 
iB02_272_v n1_4833_15584 0  0.0191328 
iB02_272_g 0 n0_4741_15584  0.0191328 
iB02_273_v n1_4833_15740 0  0.0191328 
iB02_273_g 0 n0_4741_15753  0.0191328 
iB02_274_v n1_4833_15767 0  0.0191328 
iB02_274_g 0 n0_4741_15753  0.0191328 
iB02_275_v n1_4833_15800 0  0.0191328 
iB02_275_g 0 n0_4741_15786  0.0191328 
iB02_276_v n1_5021_10799 0  0.0191328 
iB02_276_g 0 n0_4929_10785  0.0191328 
iB02_277_v n1_5021_10832 0  0.0191328 
iB02_277_g 0 n0_4929_10818  0.0191328 
iB02_278_v n1_5021_11015 0  0.0191328 
iB02_278_g 0 n0_4929_11001  0.0191328 
iB02_279_v n1_5021_11048 0  0.0191328 
iB02_279_g 0 n0_4929_11048  0.0191328 
iB02_280_v n1_5021_11182 0  0.0191328 
iB02_280_g 0 n0_4929_11217  0.0191328 
iB02_281_v n1_5021_11204 0  0.0191328 
iB02_281_g 0 n0_4929_11217  0.0191328 
iB02_282_v n1_5021_11231 0  0.0191328 
iB02_282_g 0 n0_4929_11217  0.0191328 
iB02_283_v n1_5021_11264 0  0.0191328 
iB02_283_g 0 n0_4929_11250  0.0191328 
iB02_284_v n1_5021_11447 0  0.0191328 
iB02_284_g 0 n0_4929_11433  0.0191328 
iB02_285_v n1_5021_11480 0  0.0191328 
iB02_285_g 0 n0_4929_11466  0.0191328 
iB02_286_v n1_5021_11663 0  0.0191328 
iB02_286_g 0 n0_4929_11466  0.0191328 
iB02_287_v n1_5021_11696 0  0.0191328 
iB02_287_g 0 n0_4929_11865  0.0191328 
iB02_288_v n1_5021_11879 0  0.0191328 
iB02_288_g 0 n0_4929_11865  0.0191328 
iB02_289_v n1_5021_11912 0  0.0191328 
iB02_289_g 0 n0_4929_11898  0.0191328 
iB02_290_v n1_5021_12095 0  0.0191328 
iB02_290_g 0 n0_4929_12081  0.0191328 
iB02_291_v n1_5021_12128 0  0.0191328 
iB02_291_g 0 n0_4929_12128  0.0191328 
iB02_292_v n1_5021_12284 0  0.0191328 
iB02_292_g 0 n0_4929_12297  0.0191328 
iB02_293_v n1_5021_12311 0  0.0191328 
iB02_293_g 0 n0_4929_12297  0.0191328 
iB02_294_v n1_5021_12344 0  0.0191328 
iB02_294_g 0 n0_4929_12330  0.0191328 
iB02_295_v n1_5021_12527 0  0.0191328 
iB02_295_g 0 n0_4929_12513  0.0191328 
iB02_296_v n1_5021_12560 0  0.0191328 
iB02_296_g 0 n0_4929_12546  0.0191328 
iB02_297_v n1_5021_12743 0  0.0191328 
iB02_297_g 0 n0_4929_12729  0.0191328 
iB02_298_v n1_5021_12776 0  0.0191328 
iB02_298_g 0 n0_4929_12762  0.0191328 
iB02_299_v n1_5021_12959 0  0.0191328 
iB02_299_g 0 n0_4929_12945  0.0191328 
iB02_300_v n1_5021_12992 0  0.0191328 
iB02_300_g 0 n0_4929_12978  0.0191328 
iB02_301_v n1_5021_13175 0  0.0191328 
iB02_301_g 0 n0_4929_13161  0.0191328 
iB02_302_v n1_5021_13208 0  0.0191328 
iB02_302_g 0 n0_4929_13194  0.0191328 
iB02_303_v n1_5021_13391 0  0.0191328 
iB02_303_g 0 n0_4929_13377  0.0191328 
iB02_304_v n1_5021_13424 0  0.0191328 
iB02_304_g 0 n0_4929_13424  0.0191328 
iB02_305_v n1_5021_13580 0  0.0191328 
iB02_305_g 0 n0_4929_13593  0.0191328 
iB02_306_v n1_5021_13607 0  0.0191328 
iB02_306_g 0 n0_4929_13593  0.0191328 
iB02_307_v n1_5021_13640 0  0.0191328 
iB02_307_g 0 n0_4929_13626  0.0191328 
iB02_308_v n1_5021_13823 0  0.0191328 
iB02_308_g 0 n0_4929_13809  0.0191328 
iB02_309_v n1_5021_13856 0  0.0191328 
iB02_309_g 0 n0_4929_13842  0.0191328 
iB02_310_v n1_5021_14039 0  0.0191328 
iB02_310_g 0 n0_4929_14100  0.0191328 
iB02_311_v n1_5021_14072 0  0.0191328 
iB02_311_g 0 n0_4929_14100  0.0191328 
iB02_312_v n1_5021_14206 0  0.0191328 
iB02_312_g 0 n0_4929_14241  0.0191328 
iB02_313_v n1_5021_14255 0  0.0191328 
iB02_313_g 0 n0_4929_14241  0.0191328 
iB02_314_v n1_5021_14288 0  0.0191328 
iB02_314_g 0 n0_4929_14274  0.0191328 
iB02_315_v n1_5021_14471 0  0.0191328 
iB02_315_g 0 n0_4929_14457  0.0191328 
iB02_316_v n1_5021_14504 0  0.0191328 
iB02_316_g 0 n0_4929_14490  0.0191328 
iB02_317_v n1_5021_14687 0  0.0191328 
iB02_317_g 0 n0_4929_14673  0.0191328 
iB02_318_v n1_5021_14720 0  0.0191328 
iB02_318_g 0 n0_4929_14706  0.0191328 
iB02_319_v n1_5021_14903 0  0.0191328 
iB02_319_g 0 n0_4929_14889  0.0191328 
iB02_320_v n1_5021_14936 0  0.0191328 
iB02_320_g 0 n0_4929_14922  0.0191328 
iB02_321_v n1_5021_15119 0  0.0191328 
iB02_321_g 0 n0_4929_15105  0.0191328 
iB02_322_v n1_5021_15152 0  0.0191328 
iB02_322_g 0 n0_4929_15138  0.0191328 
iB02_323_v n1_5021_15335 0  0.0191328 
iB02_323_g 0 n0_4929_15321  0.0191328 
iB02_324_v n1_5021_15368 0  0.0191328 
iB02_324_g 0 n0_4929_15368  0.0191328 
iB02_325_v n1_5021_15524 0  0.0191328 
iB02_325_g 0 n0_4929_15537  0.0191328 
iB02_326_v n1_5021_15551 0  0.0191328 
iB02_326_g 0 n0_4929_15537  0.0191328 
iB02_327_v n1_5021_15584 0  0.0191328 
iB02_327_g 0 n0_4929_15584  0.0191328 
iB02_328_v n1_5021_15740 0  0.0191328 
iB02_328_g 0 n0_4929_15753  0.0191328 
iB02_329_v n1_5021_15767 0  0.0191328 
iB02_329_g 0 n0_4929_15753  0.0191328 
iB02_330_v n1_5021_15800 0  0.0191328 
iB02_330_g 0 n0_4929_15786  0.0191328 
iB20_0_v n1_11400_215 0  0.0189263 
iB20_0_g 0 n0_10646_201  0.0189263 
iB20_1_v n1_11400_248 0  0.0189263 
iB20_1_g 0 n0_10646_234  0.0189263 
iB20_2_v n1_11400_383 0  0.0189263 
iB20_2_g 0 n0_10646_417  0.0189263 
iB20_3_v n1_11583_215 0  0.0189263 
iB20_3_g 0 n0_10646_201  0.0189263 
iB20_4_v n1_11583_248 0  0.0189263 
iB20_4_g 0 n0_10646_234  0.0189263 
iB20_5_v n1_11583_383 0  0.0189263 
iB20_5_g 0 n0_10646_417  0.0189263 
iB20_6_v n1_11400_431 0  0.0189263 
iB20_6_g 0 n0_10646_417  0.0189263 
iB20_7_v n1_11400_464 0  0.0189263 
iB20_7_g 0 n0_10646_450  0.0189263 
iB20_8_v n1_11400_647 0  0.0189263 
iB20_8_g 0 n0_10646_633  0.0189263 
iB20_9_v n1_11400_680 0  0.0189263 
iB20_9_g 0 n0_10646_666  0.0189263 
iB20_10_v n1_11583_431 0  0.0189263 
iB20_10_g 0 n0_10646_417  0.0189263 
iB20_11_v n1_11583_464 0  0.0189263 
iB20_11_g 0 n0_10646_450  0.0189263 
iB20_12_v n1_11583_647 0  0.0189263 
iB20_12_g 0 n0_10646_633  0.0189263 
iB20_13_v n1_11583_680 0  0.0189263 
iB20_13_g 0 n0_10646_666  0.0189263 
iB20_14_v n1_11630_431 0  0.0189263 
iB20_14_g 0 n0_10646_417  0.0189263 
iB20_15_v n1_11630_464 0  0.0189263 
iB20_15_g 0 n0_10646_450  0.0189263 
iB20_16_v n1_11400_863 0  0.0189263 
iB20_16_g 0 n0_10646_849  0.0189263 
iB20_17_v n1_11400_896 0  0.0189263 
iB20_17_g 0 n0_10646_882  0.0189263 
iB20_18_v n1_11400_1079 0  0.0189263 
iB20_18_g 0 n0_10646_1065  0.0189263 
iB20_19_v n1_11400_1112 0  0.0189263 
iB20_19_g 0 n0_10646_1098  0.0189263 
iB20_20_v n1_11583_863 0  0.0189263 
iB20_20_g 0 n0_10646_849  0.0189263 
iB20_21_v n1_11583_896 0  0.0189263 
iB20_21_g 0 n0_10646_882  0.0189263 
iB20_22_v n1_11583_1079 0  0.0189263 
iB20_22_g 0 n0_10646_1065  0.0189263 
iB20_23_v n1_11583_1112 0  0.0189263 
iB20_23_g 0 n0_10646_1098  0.0189263 
iB20_24_v n1_11400_1295 0  0.0189263 
iB20_24_g 0 n0_10646_1281  0.0189263 
iB20_25_v n1_11400_1328 0  0.0189263 
iB20_25_g 0 n0_10646_1314  0.0189263 
iB20_26_v n1_11400_1511 0  0.0189263 
iB20_26_g 0 n0_10646_1497  0.0189263 
iB20_27_v n1_11400_1544 0  0.0189263 
iB20_27_g 0 n0_10646_1530  0.0189263 
iB20_28_v n1_11583_1295 0  0.0189263 
iB20_28_g 0 n0_10646_1281  0.0189263 
iB20_29_v n1_11583_1328 0  0.0189263 
iB20_29_g 0 n0_10646_1314  0.0189263 
iB20_30_v n1_11400_1727 0  0.0189263 
iB20_30_g 0 n0_10646_1713  0.0189263 
iB20_31_v n1_11400_1760 0  0.0189263 
iB20_31_g 0 n0_10646_1760  0.0189263 
iB20_32_v n1_11400_1894 0  0.0189263 
iB20_32_g 0 n0_10646_1929  0.0189263 
iB20_33_v n1_11400_1943 0  0.0189263 
iB20_33_g 0 n0_10646_1929  0.0189263 
iB20_34_v n1_11400_1976 0  0.0189263 
iB20_34_g 0 n0_10646_1962  0.0189263 
iB20_35_v n1_11583_1727 0  0.0189263 
iB20_35_g 0 n0_10646_1713  0.0189263 
iB20_36_v n1_11583_1760 0  0.0189263 
iB20_36_g 0 n0_10646_1760  0.0189263 
iB20_37_v n1_11583_1894 0  0.0189263 
iB20_37_g 0 n0_10646_1929  0.0189263 
iB20_38_v n1_11583_1943 0  0.0189263 
iB20_38_g 0 n0_10646_1929  0.0189263 
iB20_39_v n1_11583_1976 0  0.0189263 
iB20_39_g 0 n0_10646_1962  0.0189263 
iB20_40_v n1_11400_2159 0  0.0189263 
iB20_40_g 0 n0_10646_2145  0.0189263 
iB20_41_v n1_11400_2192 0  0.0189263 
iB20_41_g 0 n0_10646_2178  0.0189263 
iB20_42_v n1_11400_2375 0  0.0189263 
iB20_42_g 0 n0_10646_2361  0.0189263 
iB20_43_v n1_11400_2408 0  0.0189263 
iB20_43_g 0 n0_10646_2408  0.0189263 
iB20_44_v n1_11583_2159 0  0.0189263 
iB20_44_g 0 n0_10646_2145  0.0189263 
iB20_45_v n1_11583_2192 0  0.0189263 
iB20_45_g 0 n0_10646_2178  0.0189263 
iB20_46_v n1_11583_2375 0  0.0189263 
iB20_46_g 0 n0_10646_2361  0.0189263 
iB20_47_v n1_11583_2408 0  0.0189263 
iB20_47_g 0 n0_10646_2408  0.0189263 
iB20_48_v n1_11400_2543 0  0.0189263 
iB20_48_g 0 n0_10646_2577  0.0189263 
iB20_49_v n1_11400_2591 0  0.0189263 
iB20_49_g 0 n0_10646_2577  0.0189263 
iB20_50_v n1_11400_2624 0  0.0189263 
iB20_50_g 0 n0_10646_2610  0.0189263 
iB20_51_v n1_11583_2542 0  0.0189263 
iB20_51_g 0 n0_10646_2577  0.0189263 
iB20_52_v n1_11583_2543 0  0.0189263 
iB20_52_g 0 n0_10646_2577  0.0189263 
iB20_53_v n1_11583_2591 0  0.0189263 
iB20_53_g 0 n0_10646_2577  0.0189263 
iB20_54_v n1_11583_2624 0  0.0189263 
iB20_54_g 0 n0_10646_2610  0.0189263 
iB20_55_v n1_11583_2760 0  0.0189263 
iB20_55_g 0 n0_10646_2793  0.0189263 
iB20_56_v n1_11583_2807 0  0.0189263 
iB20_56_g 0 n0_10646_2793  0.0189263 
iB20_57_v n1_11583_2840 0  0.0189263 
iB20_57_g 0 n0_10646_2840  0.0189263 
iB20_58_v n1_11630_2760 0  0.0189263 
iB20_58_g 0 n0_10646_2793  0.0189263 
iB20_59_v n1_11583_2974 0  0.0189263 
iB20_59_g 0 n0_10646_3009  0.0189263 
iB20_60_v n1_11583_3023 0  0.0189263 
iB20_60_g 0 n0_10646_3009  0.0189263 
iB20_61_v n1_11583_3056 0  0.0189263 
iB20_61_g 0 n0_10646_3042  0.0189263 
iB20_62_v n1_11583_3239 0  0.0189263 
iB20_62_g 0 n0_10646_3225  0.0189263 
iB20_63_v n1_11583_3272 0  0.0189263 
iB20_63_g 0 n0_10646_3258  0.0189263 
iB20_64_v n1_11583_3455 0  0.0189263 
iB20_64_g 0 n0_10646_3441  0.0189263 
iB20_65_v n1_11583_3488 0  0.0189263 
iB20_65_g 0 n0_10646_3488  0.0189263 
iB20_66_v n1_11583_3622 0  0.0189263 
iB20_66_g 0 n0_10646_3657  0.0189263 
iB20_67_v n1_11583_3671 0  0.0189263 
iB20_67_g 0 n0_10646_3657  0.0189263 
iB20_68_v n1_11583_3704 0  0.0189263 
iB20_68_g 0 n0_10646_3690  0.0189263 
iB20_69_v n1_11583_4103 0  0.0189263 
iB20_69_g 0 n0_10646_4089  0.0189263 
iB20_70_v n1_11583_4136 0  0.0189263 
iB20_70_g 0 n0_10646_4136  0.0189263 
iB20_71_v n1_11583_4270 0  0.0189263 
iB20_71_g 0 n0_10646_4305  0.0189263 
iB20_72_v n1_11583_4319 0  0.0189263 
iB20_72_g 0 n0_10646_4305  0.0189263 
iB20_73_v n1_11583_4352 0  0.0189263 
iB20_73_g 0 n0_10646_4338  0.0189263 
iB20_74_v n1_11583_4535 0  0.0189263 
iB20_74_g 0 n0_10646_4521  0.0189263 
iB20_75_v n1_11583_4568 0  0.0189263 
iB20_75_g 0 n0_10646_4568  0.0189263 
iB20_76_v n1_11583_4702 0  0.0189263 
iB20_76_g 0 n0_10646_4737  0.0189263 
iB20_77_v n1_11583_4751 0  0.0189263 
iB20_77_g 0 n0_10646_4737  0.0189263 
iB20_78_v n1_11583_4784 0  0.0189263 
iB20_78_g 0 n0_10646_4770  0.0189263 
iB20_79_v n1_11583_4967 0  0.0189263 
iB20_79_g 0 n0_10646_4953  0.0189263 
iB20_80_v n1_11583_5000 0  0.0189263 
iB20_80_g 0 n0_10646_4953  0.0189263 
iB20_81_v n1_11583_5183 0  0.0189263 
iB20_81_g 0 n0_10646_5169  0.0189263 
iB20_82_v n1_11583_5216 0  0.0189263 
iB20_82_g 0 n0_10646_5202  0.0189263 
iB20_83_v n1_11630_4967 0  0.0189263 
iB20_83_g 0 n0_10646_4953  0.0189263 
iB20_84_v n1_11630_5000 0  0.0189263 
iB20_84_g 0 n0_12616_5023  0.0189263 
iB20_85_v n1_11771_215 0  0.0189263 
iB20_85_g 0 n0_12616_201  0.0189263 
iB20_86_v n1_11771_248 0  0.0189263 
iB20_86_g 0 n0_12616_234  0.0189263 
iB20_87_v n1_11771_383 0  0.0189263 
iB20_87_g 0 n0_12616_417  0.0189263 
iB20_88_v n1_11864_215 0  0.0189263 
iB20_88_g 0 n0_12616_201  0.0189263 
iB20_89_v n1_11864_248 0  0.0189263 
iB20_89_g 0 n0_12616_234  0.0189263 
iB20_90_v n1_11864_383 0  0.0189263 
iB20_90_g 0 n0_12616_417  0.0189263 
iB20_91_v n1_11771_431 0  0.0189263 
iB20_91_g 0 n0_12616_417  0.0189263 
iB20_92_v n1_11771_647 0  0.0189263 
iB20_92_g 0 n0_12616_633  0.0189263 
iB20_93_v n1_11771_680 0  0.0189263 
iB20_93_g 0 n0_12616_666  0.0189263 
iB20_94_v n1_11864_431 0  0.0189263 
iB20_94_g 0 n0_12616_417  0.0189263 
iB20_95_v n1_11864_464 0  0.0189263 
iB20_95_g 0 n0_12616_450  0.0189263 
iB20_96_v n1_11864_647 0  0.0189263 
iB20_96_g 0 n0_12616_633  0.0189263 
iB20_97_v n1_11864_680 0  0.0189263 
iB20_97_g 0 n0_12616_666  0.0189263 
iB20_98_v n1_11771_863 0  0.0189263 
iB20_98_g 0 n0_12616_849  0.0189263 
iB20_99_v n1_11771_896 0  0.0189263 
iB20_99_g 0 n0_12616_882  0.0189263 
iB20_100_v n1_11771_1079 0  0.0189263 
iB20_100_g 0 n0_12616_1065  0.0189263 
iB20_101_v n1_11771_1112 0  0.0189263 
iB20_101_g 0 n0_12616_1098  0.0189263 
iB20_102_v n1_11864_863 0  0.0189263 
iB20_102_g 0 n0_12616_849  0.0189263 
iB20_103_v n1_11864_896 0  0.0189263 
iB20_103_g 0 n0_12616_882  0.0189263 
iB20_104_v n1_11864_1079 0  0.0189263 
iB20_104_g 0 n0_12616_1065  0.0189263 
iB20_105_v n1_11864_1112 0  0.0189263 
iB20_105_g 0 n0_12616_1098  0.0189263 
iB20_106_v n1_11771_1295 0  0.0189263 
iB20_106_g 0 n0_12616_1281  0.0189263 
iB20_107_v n1_11771_1328 0  0.0189263 
iB20_107_g 0 n0_12616_1314  0.0189263 
iB20_108_v n1_11771_1511 0  0.0189263 
iB20_108_g 0 n0_12616_1497  0.0189263 
iB20_109_v n1_11771_1544 0  0.0189263 
iB20_109_g 0 n0_12616_1530  0.0189263 
iB20_110_v n1_11864_1295 0  0.0189263 
iB20_110_g 0 n0_12616_1281  0.0189263 
iB20_111_v n1_11864_1328 0  0.0189263 
iB20_111_g 0 n0_12616_1314  0.0189263 
iB20_112_v n1_11864_1511 0  0.0189263 
iB20_112_g 0 n0_12616_1497  0.0189263 
iB20_113_v n1_11864_1544 0  0.0189263 
iB20_113_g 0 n0_12616_1530  0.0189263 
iB20_114_v n1_11771_1727 0  0.0189263 
iB20_114_g 0 n0_12616_1713  0.0189263 
iB20_115_v n1_11771_1760 0  0.0189263 
iB20_115_g 0 n0_12616_1746  0.0189263 
iB20_116_v n1_11771_1894 0  0.0189263 
iB20_116_g 0 n0_12616_1929  0.0189263 
iB20_117_v n1_11771_1943 0  0.0189263 
iB20_117_g 0 n0_12616_1929  0.0189263 
iB20_118_v n1_11771_1976 0  0.0189263 
iB20_118_g 0 n0_12616_1962  0.0189263 
iB20_119_v n1_11864_1727 0  0.0189263 
iB20_119_g 0 n0_12616_1713  0.0189263 
iB20_120_v n1_11864_1760 0  0.0189263 
iB20_120_g 0 n0_12616_1746  0.0189263 
iB20_121_v n1_11864_1894 0  0.0189263 
iB20_121_g 0 n0_12616_1929  0.0189263 
iB20_122_v n1_11864_1943 0  0.0189263 
iB20_122_g 0 n0_12616_1929  0.0189263 
iB20_123_v n1_11864_1976 0  0.0189263 
iB20_123_g 0 n0_12616_1962  0.0189263 
iB20_124_v n1_11771_2159 0  0.0189263 
iB20_124_g 0 n0_12616_2145  0.0189263 
iB20_125_v n1_11771_2192 0  0.0189263 
iB20_125_g 0 n0_12616_2178  0.0189263 
iB20_126_v n1_11771_2375 0  0.0189263 
iB20_126_g 0 n0_12616_2361  0.0189263 
iB20_127_v n1_11771_2408 0  0.0189263 
iB20_127_g 0 n0_12616_2394  0.0189263 
iB20_128_v n1_11864_2159 0  0.0189263 
iB20_128_g 0 n0_12616_2145  0.0189263 
iB20_129_v n1_11864_2192 0  0.0189263 
iB20_129_g 0 n0_12616_2178  0.0189263 
iB20_130_v n1_11864_2375 0  0.0189263 
iB20_130_g 0 n0_12616_2361  0.0189263 
iB20_131_v n1_11864_2408 0  0.0189263 
iB20_131_g 0 n0_12616_2394  0.0189263 
iB20_132_v n1_11771_2542 0  0.0189263 
iB20_132_g 0 n0_12616_2577  0.0189263 
iB20_133_v n1_11771_2543 0  0.0189263 
iB20_133_g 0 n0_12616_2577  0.0189263 
iB20_134_v n1_11771_2591 0  0.0189263 
iB20_134_g 0 n0_12616_2577  0.0189263 
iB20_135_v n1_11771_2624 0  0.0189263 
iB20_135_g 0 n0_12616_2610  0.0189263 
iB20_136_v n1_11771_2760 0  0.0189263 
iB20_136_g 0 n0_12616_2793  0.0189263 
iB20_137_v n1_11771_2807 0  0.0189263 
iB20_137_g 0 n0_12616_2793  0.0189263 
iB20_138_v n1_11771_2840 0  0.0189263 
iB20_138_g 0 n0_12616_2826  0.0189263 
iB20_139_v n1_11864_2542 0  0.0189263 
iB20_139_g 0 n0_12616_2577  0.0189263 
iB20_140_v n1_11864_2543 0  0.0189263 
iB20_140_g 0 n0_12616_2577  0.0189263 
iB20_141_v n1_11864_2591 0  0.0189263 
iB20_141_g 0 n0_12616_2577  0.0189263 
iB20_142_v n1_11864_2624 0  0.0189263 
iB20_142_g 0 n0_12616_2610  0.0189263 
iB20_143_v n1_11771_2974 0  0.0189263 
iB20_143_g 0 n0_12616_3009  0.0189263 
iB20_144_v n1_11771_3023 0  0.0189263 
iB20_144_g 0 n0_12616_3009  0.0189263 
iB20_145_v n1_11771_3056 0  0.0189263 
iB20_145_g 0 n0_12616_3042  0.0189263 
iB20_146_v n1_11771_3239 0  0.0189263 
iB20_146_g 0 n0_12616_3225  0.0189263 
iB20_147_v n1_11771_3272 0  0.0189263 
iB20_147_g 0 n0_12616_3258  0.0189263 
iB20_148_v n1_11771_3455 0  0.0189263 
iB20_148_g 0 n0_12616_3441  0.0189263 
iB20_149_v n1_11771_3488 0  0.0189263 
iB20_149_g 0 n0_12616_3474  0.0189263 
iB20_150_v n1_11771_3622 0  0.0189263 
iB20_150_g 0 n0_12616_3657  0.0189263 
iB20_151_v n1_11771_3671 0  0.0189263 
iB20_151_g 0 n0_12616_3657  0.0189263 
iB20_152_v n1_11771_3704 0  0.0189263 
iB20_152_g 0 n0_12616_3690  0.0189263 
iB20_153_v n1_11771_3887 0  0.0189263 
iB20_153_g 0 n0_12616_3873  0.0189263 
iB20_154_v n1_11771_3920 0  0.0189263 
iB20_154_g 0 n0_12616_3906  0.0189263 
iB20_155_v n1_11771_4103 0  0.0189263 
iB20_155_g 0 n0_12616_4089  0.0189263 
iB20_156_v n1_11771_4136 0  0.0189263 
iB20_156_g 0 n0_12616_4122  0.0189263 
iB20_157_v n1_11771_4270 0  0.0189263 
iB20_157_g 0 n0_12616_4305  0.0189263 
iB20_158_v n1_11771_4319 0  0.0189263 
iB20_158_g 0 n0_12616_4305  0.0189263 
iB20_159_v n1_11771_4352 0  0.0189263 
iB20_159_g 0 n0_12616_4338  0.0189263 
iB20_160_v n1_11771_4535 0  0.0189263 
iB20_160_g 0 n0_12616_4521  0.0189263 
iB20_161_v n1_11771_4568 0  0.0189263 
iB20_161_g 0 n0_12616_4554  0.0189263 
iB20_162_v n1_11771_4702 0  0.0189263 
iB20_162_g 0 n0_12616_4737  0.0189263 
iB20_163_v n1_11771_4751 0  0.0189263 
iB20_163_g 0 n0_12616_4737  0.0189263 
iB20_164_v n1_11771_4784 0  0.0189263 
iB20_164_g 0 n0_12616_4770  0.0189263 
iB20_165_v n1_11771_5000 0  0.0189263 
iB20_165_g 0 n0_12616_5023  0.0189263 
iB20_166_v n1_11771_5183 0  0.0189263 
iB20_166_g 0 n0_12616_5169  0.0189263 
iB20_167_v n1_11771_5216 0  0.0189263 
iB20_167_g 0 n0_12616_5202  0.0189263 
iB20_168_v n1_13650_215 0  0.0189263 
iB20_168_g 0 n0_12896_201  0.0189263 
iB20_169_v n1_13650_248 0  0.0189263 
iB20_169_g 0 n0_12896_234  0.0189263 
iB20_170_v n1_13650_383 0  0.0189263 
iB20_170_g 0 n0_12896_417  0.0189263 
iB20_171_v n1_13650_431 0  0.0189263 
iB20_171_g 0 n0_12896_417  0.0189263 
iB20_172_v n1_13650_464 0  0.0189263 
iB20_172_g 0 n0_12896_450  0.0189263 
iB20_173_v n1_13650_647 0  0.0189263 
iB20_173_g 0 n0_12896_633  0.0189263 
iB20_174_v n1_13650_680 0  0.0189263 
iB20_174_g 0 n0_12896_666  0.0189263 
iB20_175_v n1_13650_863 0  0.0189263 
iB20_175_g 0 n0_12896_849  0.0189263 
iB20_176_v n1_13650_896 0  0.0189263 
iB20_176_g 0 n0_12896_882  0.0189263 
iB20_177_v n1_13650_1079 0  0.0189263 
iB20_177_g 0 n0_12896_1065  0.0189263 
iB20_178_v n1_13650_1112 0  0.0189263 
iB20_178_g 0 n0_12896_1098  0.0189263 
iB20_179_v n1_13650_1295 0  0.0189263 
iB20_179_g 0 n0_12896_1281  0.0189263 
iB20_180_v n1_13650_1328 0  0.0189263 
iB20_180_g 0 n0_12896_1314  0.0189263 
iB20_181_v n1_13650_1511 0  0.0189263 
iB20_181_g 0 n0_12896_1497  0.0189263 
iB20_182_v n1_13650_1544 0  0.0189263 
iB20_182_g 0 n0_12896_1530  0.0189263 
iB20_183_v n1_13650_1727 0  0.0189263 
iB20_183_g 0 n0_12896_1713  0.0189263 
iB20_184_v n1_13650_1760 0  0.0189263 
iB20_184_g 0 n0_12896_1746  0.0189263 
iB20_185_v n1_13650_1894 0  0.0189263 
iB20_185_g 0 n0_12896_1929  0.0189263 
iB20_186_v n1_13650_1943 0  0.0189263 
iB20_186_g 0 n0_12896_1929  0.0189263 
iB20_187_v n1_13650_1976 0  0.0189263 
iB20_187_g 0 n0_12896_1962  0.0189263 
iB20_188_v n1_13650_2159 0  0.0189263 
iB20_188_g 0 n0_12896_2145  0.0189263 
iB20_189_v n1_13650_2192 0  0.0189263 
iB20_189_g 0 n0_12896_2178  0.0189263 
iB20_190_v n1_13650_2375 0  0.0189263 
iB20_190_g 0 n0_12896_2361  0.0189263 
iB20_191_v n1_13650_2408 0  0.0189263 
iB20_191_g 0 n0_12896_2394  0.0189263 
iB20_192_v n1_13650_2445 0  0.0189263 
iB20_192_g 0 n0_12896_2431  0.0189263 
iB20_193_v n1_13650_2542 0  0.0189263 
iB20_193_g 0 n0_12896_2577  0.0189263 
iB20_194_v n1_13650_2543 0  0.0189263 
iB20_194_g 0 n0_12896_2577  0.0189263 
iB20_195_v n1_13650_2591 0  0.0189263 
iB20_195_g 0 n0_12896_2577  0.0189263 
iB20_196_v n1_13650_2624 0  0.0189263 
iB20_196_g 0 n0_12896_2610  0.0189263 
iB20_197_v n1_13833_215 0  0.0189263 
iB20_197_g 0 n0_12896_201  0.0189263 
iB20_198_v n1_13833_248 0  0.0189263 
iB20_198_g 0 n0_12896_234  0.0189263 
iB20_199_v n1_13833_383 0  0.0189263 
iB20_199_g 0 n0_12896_417  0.0189263 
iB20_200_v n1_14021_215 0  0.0189263 
iB20_200_g 0 n0_14866_201  0.0189263 
iB20_201_v n1_14021_248 0  0.0189263 
iB20_201_g 0 n0_14866_234  0.0189263 
iB20_202_v n1_14021_383 0  0.0189263 
iB20_202_g 0 n0_14866_417  0.0189263 
iB20_203_v n1_14114_215 0  0.0189263 
iB20_203_g 0 n0_14866_201  0.0189263 
iB20_204_v n1_14114_248 0  0.0189263 
iB20_204_g 0 n0_14866_234  0.0189263 
iB20_205_v n1_14114_383 0  0.0189263 
iB20_205_g 0 n0_14866_417  0.0189263 
iB20_206_v n1_13833_431 0  0.0189263 
iB20_206_g 0 n0_12896_417  0.0189263 
iB20_207_v n1_13833_464 0  0.0189263 
iB20_207_g 0 n0_12896_450  0.0189263 
iB20_208_v n1_13833_647 0  0.0189263 
iB20_208_g 0 n0_12896_633  0.0189263 
iB20_209_v n1_13833_680 0  0.0189263 
iB20_209_g 0 n0_12896_666  0.0189263 
iB20_210_v n1_13880_431 0  0.0189263 
iB20_210_g 0 n0_12896_417  0.0189263 
iB20_211_v n1_13880_464 0  0.0189263 
iB20_211_g 0 n0_12896_450  0.0189263 
iB20_212_v n1_14021_431 0  0.0189263 
iB20_212_g 0 n0_14866_417  0.0189263 
iB20_213_v n1_14021_647 0  0.0189263 
iB20_213_g 0 n0_14866_633  0.0189263 
iB20_214_v n1_14021_680 0  0.0189263 
iB20_214_g 0 n0_14866_666  0.0189263 
iB20_215_v n1_14114_431 0  0.0189263 
iB20_215_g 0 n0_14866_417  0.0189263 
iB20_216_v n1_14114_464 0  0.0189263 
iB20_216_g 0 n0_14866_450  0.0189263 
iB20_217_v n1_14114_647 0  0.0189263 
iB20_217_g 0 n0_14866_633  0.0189263 
iB20_218_v n1_14114_680 0  0.0189263 
iB20_218_g 0 n0_14866_666  0.0189263 
iB20_219_v n1_13833_863 0  0.0189263 
iB20_219_g 0 n0_12896_849  0.0189263 
iB20_220_v n1_13833_896 0  0.0189263 
iB20_220_g 0 n0_12896_882  0.0189263 
iB20_221_v n1_13833_1079 0  0.0189263 
iB20_221_g 0 n0_12896_1065  0.0189263 
iB20_222_v n1_13833_1112 0  0.0189263 
iB20_222_g 0 n0_12896_1098  0.0189263 
iB20_223_v n1_14021_863 0  0.0189263 
iB20_223_g 0 n0_14866_849  0.0189263 
iB20_224_v n1_14021_896 0  0.0189263 
iB20_224_g 0 n0_14866_882  0.0189263 
iB20_225_v n1_14021_1079 0  0.0189263 
iB20_225_g 0 n0_14866_1065  0.0189263 
iB20_226_v n1_14021_1112 0  0.0189263 
iB20_226_g 0 n0_14866_1098  0.0189263 
iB20_227_v n1_14114_863 0  0.0189263 
iB20_227_g 0 n0_14866_849  0.0189263 
iB20_228_v n1_14114_896 0  0.0189263 
iB20_228_g 0 n0_14866_882  0.0189263 
iB20_229_v n1_14114_1079 0  0.0189263 
iB20_229_g 0 n0_14866_1065  0.0189263 
iB20_230_v n1_14114_1112 0  0.0189263 
iB20_230_g 0 n0_14866_1098  0.0189263 
iB20_231_v n1_13833_1295 0  0.0189263 
iB20_231_g 0 n0_12896_1281  0.0189263 
iB20_232_v n1_13833_1328 0  0.0189263 
iB20_232_g 0 n0_12896_1314  0.0189263 
iB20_233_v n1_14021_1295 0  0.0189263 
iB20_233_g 0 n0_14866_1281  0.0189263 
iB20_234_v n1_14021_1328 0  0.0189263 
iB20_234_g 0 n0_14866_1314  0.0189263 
iB20_235_v n1_14021_1511 0  0.0189263 
iB20_235_g 0 n0_14866_1497  0.0189263 
iB20_236_v n1_14021_1544 0  0.0189263 
iB20_236_g 0 n0_14866_1530  0.0189263 
iB20_237_v n1_14114_1295 0  0.0189263 
iB20_237_g 0 n0_14866_1281  0.0189263 
iB20_238_v n1_14114_1328 0  0.0189263 
iB20_238_g 0 n0_14866_1314  0.0189263 
iB20_239_v n1_14114_1511 0  0.0189263 
iB20_239_g 0 n0_14866_1497  0.0189263 
iB20_240_v n1_14114_1544 0  0.0189263 
iB20_240_g 0 n0_14866_1530  0.0189263 
iB20_241_v n1_13833_1727 0  0.0189263 
iB20_241_g 0 n0_12896_1713  0.0189263 
iB20_242_v n1_13833_1760 0  0.0189263 
iB20_242_g 0 n0_12896_1746  0.0189263 
iB20_243_v n1_13833_1894 0  0.0189263 
iB20_243_g 0 n0_12896_1929  0.0189263 
iB20_244_v n1_13833_1943 0  0.0189263 
iB20_244_g 0 n0_12896_1929  0.0189263 
iB20_245_v n1_13833_1976 0  0.0189263 
iB20_245_g 0 n0_12896_1962  0.0189263 
iB20_246_v n1_14021_1727 0  0.0189263 
iB20_246_g 0 n0_14866_1713  0.0189263 
iB20_247_v n1_14021_1760 0  0.0189263 
iB20_247_g 0 n0_14866_1746  0.0189263 
iB20_248_v n1_14021_1894 0  0.0189263 
iB20_248_g 0 n0_14866_1929  0.0189263 
iB20_249_v n1_14021_1943 0  0.0189263 
iB20_249_g 0 n0_14866_1929  0.0189263 
iB20_250_v n1_14021_1976 0  0.0189263 
iB20_250_g 0 n0_14866_1962  0.0189263 
iB20_251_v n1_14114_1727 0  0.0189263 
iB20_251_g 0 n0_14866_1713  0.0189263 
iB20_252_v n1_14114_1760 0  0.0189263 
iB20_252_g 0 n0_14866_1746  0.0189263 
iB20_253_v n1_14114_1894 0  0.0189263 
iB20_253_g 0 n0_14866_1929  0.0189263 
iB20_254_v n1_14114_1943 0  0.0189263 
iB20_254_g 0 n0_14866_1929  0.0189263 
iB20_255_v n1_14114_1976 0  0.0189263 
iB20_255_g 0 n0_14866_1962  0.0189263 
iB20_256_v n1_13833_2159 0  0.0189263 
iB20_256_g 0 n0_12896_2145  0.0189263 
iB20_257_v n1_13833_2192 0  0.0189263 
iB20_257_g 0 n0_12896_2178  0.0189263 
iB20_258_v n1_13833_2375 0  0.0189263 
iB20_258_g 0 n0_12896_2361  0.0189263 
iB20_259_v n1_13833_2408 0  0.0189263 
iB20_259_g 0 n0_12896_2394  0.0189263 
iB20_260_v n1_13833_2445 0  0.0189263 
iB20_260_g 0 n0_12896_2431  0.0189263 
iB20_261_v n1_14021_2159 0  0.0189263 
iB20_261_g 0 n0_14866_2145  0.0189263 
iB20_262_v n1_14021_2192 0  0.0189263 
iB20_262_g 0 n0_14866_2178  0.0189263 
iB20_263_v n1_14021_2375 0  0.0189263 
iB20_263_g 0 n0_14866_2361  0.0189263 
iB20_264_v n1_14021_2408 0  0.0189263 
iB20_264_g 0 n0_14866_2394  0.0189263 
iB20_265_v n1_14021_2445 0  0.0189263 
iB20_265_g 0 n0_14866_2431  0.0189263 
iB20_266_v n1_14114_2159 0  0.0189263 
iB20_266_g 0 n0_14866_2145  0.0189263 
iB20_267_v n1_14114_2192 0  0.0189263 
iB20_267_g 0 n0_14866_2178  0.0189263 
iB20_268_v n1_14114_2375 0  0.0189263 
iB20_268_g 0 n0_14866_2361  0.0189263 
iB20_269_v n1_14114_2408 0  0.0189263 
iB20_269_g 0 n0_14866_2394  0.0189263 
iB20_270_v n1_14114_2445 0  0.0189263 
iB20_270_g 0 n0_14866_2431  0.0189263 
iB20_271_v n1_13833_2542 0  0.0189263 
iB20_271_g 0 n0_12896_2577  0.0189263 
iB20_272_v n1_13833_2543 0  0.0189263 
iB20_272_g 0 n0_12896_2577  0.0189263 
iB20_273_v n1_13833_2591 0  0.0189263 
iB20_273_g 0 n0_12896_2577  0.0189263 
iB20_274_v n1_13833_2624 0  0.0189263 
iB20_274_g 0 n0_12896_2610  0.0189263 
iB20_275_v n1_13833_2807 0  0.0189263 
iB20_275_g 0 n0_12896_2793  0.0189263 
iB20_276_v n1_13833_2840 0  0.0189263 
iB20_276_g 0 n0_12896_2826  0.0189263 
iB20_277_v n1_14021_2542 0  0.0189263 
iB20_277_g 0 n0_14866_2577  0.0189263 
iB20_278_v n1_14021_2543 0  0.0189263 
iB20_278_g 0 n0_14866_2577  0.0189263 
iB20_279_v n1_14021_2591 0  0.0189263 
iB20_279_g 0 n0_14866_2577  0.0189263 
iB20_280_v n1_14021_2624 0  0.0189263 
iB20_280_g 0 n0_14866_2610  0.0189263 
iB20_281_v n1_14021_2807 0  0.0189263 
iB20_281_g 0 n0_14866_2793  0.0189263 
iB20_282_v n1_14021_2840 0  0.0189263 
iB20_282_g 0 n0_14866_2826  0.0189263 
iB20_283_v n1_14114_2542 0  0.0189263 
iB20_283_g 0 n0_14866_2577  0.0189263 
iB20_284_v n1_14114_2543 0  0.0189263 
iB20_284_g 0 n0_14866_2577  0.0189263 
iB20_285_v n1_14114_2591 0  0.0189263 
iB20_285_g 0 n0_14866_2577  0.0189263 
iB20_286_v n1_14114_2624 0  0.0189263 
iB20_286_g 0 n0_14866_2610  0.0189263 
iB20_287_v n1_13833_2877 0  0.0189263 
iB20_287_g 0 n0_12896_2863  0.0189263 
iB20_288_v n1_13833_2974 0  0.0189263 
iB20_288_g 0 n0_12896_3009  0.0189263 
iB20_289_v n1_13833_3023 0  0.0189263 
iB20_289_g 0 n0_12896_3009  0.0189263 
iB20_290_v n1_13833_3056 0  0.0189263 
iB20_290_g 0 n0_12896_3042  0.0189263 
iB20_291_v n1_13833_3239 0  0.0189263 
iB20_291_g 0 n0_12896_3225  0.0189263 
iB20_292_v n1_14021_2877 0  0.0189263 
iB20_292_g 0 n0_14866_2863  0.0189263 
iB20_293_v n1_14021_2974 0  0.0189263 
iB20_293_g 0 n0_14866_3009  0.0189263 
iB20_294_v n1_14021_3023 0  0.0189263 
iB20_294_g 0 n0_14866_3009  0.0189263 
iB20_295_v n1_14021_3056 0  0.0189263 
iB20_295_g 0 n0_14866_3042  0.0189263 
iB20_296_v n1_14021_3239 0  0.0189263 
iB20_296_g 0 n0_14866_3225  0.0189263 
iB20_297_v n1_13833_3272 0  0.0189263 
iB20_297_g 0 n0_12896_3258  0.0189263 
iB20_298_v n1_13833_3455 0  0.0189263 
iB20_298_g 0 n0_12896_3441  0.0189263 
iB20_299_v n1_13833_3488 0  0.0189263 
iB20_299_g 0 n0_12896_3474  0.0189263 
iB20_300_v n1_13833_3622 0  0.0189263 
iB20_300_g 0 n0_12896_3657  0.0189263 
iB20_301_v n1_13833_3671 0  0.0189263 
iB20_301_g 0 n0_12896_3657  0.0189263 
iB20_302_v n1_14021_3272 0  0.0189263 
iB20_302_g 0 n0_14866_3258  0.0189263 
iB20_303_v n1_14021_3455 0  0.0189263 
iB20_303_g 0 n0_14866_3441  0.0189263 
iB20_304_v n1_14021_3488 0  0.0189263 
iB20_304_g 0 n0_14866_3474  0.0189263 
iB20_305_v n1_14021_3622 0  0.0189263 
iB20_305_g 0 n0_14866_3657  0.0189263 
iB20_306_v n1_14021_3671 0  0.0189263 
iB20_306_g 0 n0_14866_3657  0.0189263 
iB20_307_v n1_13833_3704 0  0.0189263 
iB20_307_g 0 n0_12896_3690  0.0189263 
iB20_308_v n1_13833_4054 0  0.0189263 
iB20_308_g 0 n0_12896_4089  0.0189263 
iB20_309_v n1_14021_3704 0  0.0189263 
iB20_309_g 0 n0_14866_3690  0.0189263 
iB20_310_v n1_14021_3887 0  0.0189263 
iB20_310_g 0 n0_14866_3873  0.0189263 
iB20_311_v n1_14021_3920 0  0.0189263 
iB20_311_g 0 n0_14866_3906  0.0189263 
iB20_312_v n1_14021_4054 0  0.0189263 
iB20_312_g 0 n0_14866_4089  0.0189263 
iB20_313_v n1_13833_4103 0  0.0189263 
iB20_313_g 0 n0_12896_4089  0.0189263 
iB20_314_v n1_13833_4136 0  0.0189263 
iB20_314_g 0 n0_12896_4122  0.0189263 
iB20_315_v n1_13833_4270 0  0.0189263 
iB20_315_g 0 n0_12896_4305  0.0189263 
iB20_316_v n1_13833_4319 0  0.0189263 
iB20_316_g 0 n0_12896_4305  0.0189263 
iB20_317_v n1_13833_4352 0  0.0189263 
iB20_317_g 0 n0_12896_4338  0.0189263 
iB20_318_v n1_14021_4103 0  0.0189263 
iB20_318_g 0 n0_14866_4089  0.0189263 
iB20_319_v n1_14021_4136 0  0.0189263 
iB20_319_g 0 n0_14866_4122  0.0189263 
iB20_320_v n1_14021_4270 0  0.0189263 
iB20_320_g 0 n0_14866_4305  0.0189263 
iB20_321_v n1_14021_4319 0  0.0189263 
iB20_321_g 0 n0_14866_4305  0.0189263 
iB20_322_v n1_14021_4352 0  0.0189263 
iB20_322_g 0 n0_14866_4338  0.0189263 
iB20_323_v n1_13833_4535 0  0.0189263 
iB20_323_g 0 n0_12896_4521  0.0189263 
iB20_324_v n1_13833_4568 0  0.0189263 
iB20_324_g 0 n0_12896_4554  0.0189263 
iB20_325_v n1_13833_4702 0  0.0189263 
iB20_325_g 0 n0_12896_4737  0.0189263 
iB20_326_v n1_13833_4751 0  0.0189263 
iB20_326_g 0 n0_12896_4737  0.0189263 
iB20_327_v n1_13833_4784 0  0.0189263 
iB20_327_g 0 n0_12896_4770  0.0189263 
iB20_328_v n1_14021_4535 0  0.0189263 
iB20_328_g 0 n0_14866_4521  0.0189263 
iB20_329_v n1_14021_4568 0  0.0189263 
iB20_329_g 0 n0_14866_4554  0.0189263 
iB20_330_v n1_14021_4702 0  0.0189263 
iB20_330_g 0 n0_14866_4737  0.0189263 
iB20_331_v n1_14021_4751 0  0.0189263 
iB20_331_g 0 n0_14866_4737  0.0189263 
iB20_332_v n1_14021_4784 0  0.0189263 
iB20_332_g 0 n0_14866_4770  0.0189263 
iB20_333_v n1_13833_4967 0  0.0189263 
iB20_333_g 0 n0_12896_4953  0.0189263 
iB20_334_v n1_13833_5000 0  0.0189263 
iB20_334_g 0 n0_12896_5023  0.0189263 
iB20_335_v n1_13833_5134 0  0.0189263 
iB20_335_g 0 n0_12896_5169  0.0189263 
iB20_336_v n1_13833_5183 0  0.0189263 
iB20_336_g 0 n0_12896_5169  0.0189263 
iB20_337_v n1_13833_5216 0  0.0189263 
iB20_337_g 0 n0_12896_5202  0.0189263 
iB20_338_v n1_13880_4967 0  0.0189263 
iB20_338_g 0 n0_12896_4953  0.0189263 
iB20_339_v n1_13880_5000 0  0.0189263 
iB20_339_g 0 n0_12896_5023  0.0189263 
iB20_340_v n1_14021_5000 0  0.0189263 
iB20_340_g 0 n0_14866_4953  0.0189263 
iB20_341_v n1_14021_5134 0  0.0189263 
iB20_341_g 0 n0_14866_5169  0.0189263 
iB20_342_v n1_14021_5183 0  0.0189263 
iB20_342_g 0 n0_14866_5169  0.0189263 
iB20_343_v n1_14021_5216 0  0.0189263 
iB20_343_g 0 n0_14866_5202  0.0189263 
iB20_344_v n1_15900_215 0  0.0189263 
iB20_344_g 0 n0_15146_201  0.0189263 
iB20_345_v n1_15900_248 0  0.0189263 
iB20_345_g 0 n0_15146_234  0.0189263 
iB20_346_v n1_15900_383 0  0.0189263 
iB20_346_g 0 n0_15146_417  0.0189263 
iB20_347_v n1_15900_431 0  0.0189263 
iB20_347_g 0 n0_15146_417  0.0189263 
iB20_348_v n1_15900_464 0  0.0189263 
iB20_348_g 0 n0_15146_450  0.0189263 
iB20_349_v n1_15900_647 0  0.0189263 
iB20_349_g 0 n0_15146_633  0.0189263 
iB20_350_v n1_15900_680 0  0.0189263 
iB20_350_g 0 n0_15146_666  0.0189263 
iB20_351_v n1_15900_863 0  0.0189263 
iB20_351_g 0 n0_15146_849  0.0189263 
iB20_352_v n1_15900_896 0  0.0189263 
iB20_352_g 0 n0_15146_882  0.0189263 
iB20_353_v n1_15900_1079 0  0.0189263 
iB20_353_g 0 n0_15146_1065  0.0189263 
iB20_354_v n1_15900_1112 0  0.0189263 
iB20_354_g 0 n0_15146_1098  0.0189263 
iB20_355_v n1_15900_1295 0  0.0189263 
iB20_355_g 0 n0_15146_1281  0.0189263 
iB20_356_v n1_15900_1328 0  0.0189263 
iB20_356_g 0 n0_15146_1314  0.0189263 
iB20_357_v n1_15900_1511 0  0.0189263 
iB20_357_g 0 n0_15146_1497  0.0189263 
iB20_358_v n1_15900_1544 0  0.0189263 
iB20_358_g 0 n0_15146_1530  0.0189263 
iB20_359_v n1_15900_1727 0  0.0189263 
iB20_359_g 0 n0_15146_1713  0.0189263 
iB20_360_v n1_15900_1760 0  0.0189263 
iB20_360_g 0 n0_15146_1746  0.0189263 
iB20_361_v n1_15900_1894 0  0.0189263 
iB20_361_g 0 n0_15146_1929  0.0189263 
iB20_362_v n1_15900_1943 0  0.0189263 
iB20_362_g 0 n0_15146_1929  0.0189263 
iB20_363_v n1_15900_1976 0  0.0189263 
iB20_363_g 0 n0_15146_1962  0.0189263 
iB20_364_v n1_15900_2159 0  0.0189263 
iB20_364_g 0 n0_15146_2145  0.0189263 
iB20_365_v n1_15900_2192 0  0.0189263 
iB20_365_g 0 n0_15146_2178  0.0189263 
iB20_366_v n1_15900_2375 0  0.0189263 
iB20_366_g 0 n0_15146_2361  0.0189263 
iB20_367_v n1_15900_2408 0  0.0189263 
iB20_367_g 0 n0_15146_2394  0.0189263 
iB20_368_v n1_15900_2445 0  0.0189263 
iB20_368_g 0 n0_15146_2431  0.0189263 
iB20_369_v n1_15900_2542 0  0.0189263 
iB20_369_g 0 n0_15146_2577  0.0189263 
iB20_370_v n1_15900_2543 0  0.0189263 
iB20_370_g 0 n0_15146_2577  0.0189263 
iB20_371_v n1_15900_2591 0  0.0189263 
iB20_371_g 0 n0_15146_2577  0.0189263 
iB20_372_v n1_15900_2624 0  0.0189263 
iB20_372_g 0 n0_15146_2610  0.0189263 
iB03_0_v n1_333_15983 0  0.021569 
iB03_0_g 0 n0_241_15969  0.021569 
iB03_1_v n1_333_16016 0  0.021569 
iB03_1_g 0 n0_241_16002  0.021569 
iB03_2_v n1_333_16199 0  0.021569 
iB03_2_g 0 n0_241_16185  0.021569 
iB03_3_v n1_333_16232 0  0.021569 
iB03_3_g 0 n0_241_16218  0.021569 
iB03_4_v n1_380_16199 0  0.021569 
iB03_4_g 0 n0_241_16185  0.021569 
iB03_5_v n1_380_16232 0  0.021569 
iB03_5_g 0 n0_241_16218  0.021569 
iB03_6_v n1_521_15983 0  0.021569 
iB03_6_g 0 n0_429_15969  0.021569 
iB03_7_v n1_521_16016 0  0.021569 
iB03_7_g 0 n0_429_16002  0.021569 
iB03_8_v n1_521_16199 0  0.021569 
iB03_8_g 0 n0_429_16002  0.021569 
iB03_9_v n1_333_16415 0  0.021569 
iB03_9_g 0 n0_241_16401  0.021569 
iB03_10_v n1_333_16448 0  0.021569 
iB03_10_g 0 n0_241_16434  0.021569 
iB03_11_v n1_333_16631 0  0.021569 
iB03_11_g 0 n0_241_16617  0.021569 
iB03_12_v n1_333_16664 0  0.021569 
iB03_12_g 0 n0_241_16650  0.021569 
iB03_13_v n1_521_16415 0  0.021569 
iB03_13_g 0 n0_429_16401  0.021569 
iB03_14_v n1_521_16448 0  0.021569 
iB03_14_g 0 n0_429_16434  0.021569 
iB03_15_v n1_521_16631 0  0.021569 
iB03_15_g 0 n0_429_16617  0.021569 
iB03_16_v n1_521_16664 0  0.021569 
iB03_16_g 0 n0_429_16650  0.021569 
iB03_17_v n1_333_16847 0  0.021569 
iB03_17_g 0 n0_241_16833  0.021569 
iB03_18_v n1_333_16880 0  0.021569 
iB03_18_g 0 n0_241_16866  0.021569 
iB03_19_v n1_333_17063 0  0.021569 
iB03_19_g 0 n0_241_17049  0.021569 
iB03_20_v n1_333_17096 0  0.021569 
iB03_20_g 0 n0_241_17082  0.021569 
iB03_21_v n1_521_16847 0  0.021569 
iB03_21_g 0 n0_429_16833  0.021569 
iB03_22_v n1_521_16880 0  0.021569 
iB03_22_g 0 n0_429_16866  0.021569 
iB03_23_v n1_521_17063 0  0.021569 
iB03_23_g 0 n0_429_17049  0.021569 
iB03_24_v n1_521_17096 0  0.021569 
iB03_24_g 0 n0_429_17082  0.021569 
iB03_25_v n1_333_17495 0  0.021569 
iB03_25_g 0 n0_241_17481  0.021569 
iB03_26_v n1_521_17279 0  0.021569 
iB03_26_g 0 n0_429_17265  0.021569 
iB03_27_v n1_521_17312 0  0.021569 
iB03_27_g 0 n0_429_17298  0.021569 
iB03_28_v n1_521_17495 0  0.021569 
iB03_28_g 0 n0_429_17481  0.021569 
iB03_29_v n1_333_17528 0  0.021569 
iB03_29_g 0 n0_241_17514  0.021569 
iB03_30_v n1_333_17711 0  0.021569 
iB03_30_g 0 n0_241_17697  0.021569 
iB03_31_v n1_333_17744 0  0.021569 
iB03_31_g 0 n0_241_17730  0.021569 
iB03_32_v n1_333_17927 0  0.021569 
iB03_32_g 0 n0_241_17913  0.021569 
iB03_33_v n1_521_17528 0  0.021569 
iB03_33_g 0 n0_429_17514  0.021569 
iB03_34_v n1_521_17711 0  0.021569 
iB03_34_g 0 n0_429_17697  0.021569 
iB03_35_v n1_521_17744 0  0.021569 
iB03_35_g 0 n0_429_17730  0.021569 
iB03_36_v n1_521_17927 0  0.021569 
iB03_36_g 0 n0_429_17913  0.021569 
iB03_37_v n1_333_17960 0  0.021569 
iB03_37_g 0 n0_241_17960  0.021569 
iB03_38_v n1_333_18116 0  0.021569 
iB03_38_g 0 n0_241_18129  0.021569 
iB03_39_v n1_333_18143 0  0.021569 
iB03_39_g 0 n0_241_18129  0.021569 
iB03_40_v n1_333_18176 0  0.021569 
iB03_40_g 0 n0_241_18162  0.021569 
iB03_41_v n1_521_17960 0  0.021569 
iB03_41_g 0 n0_429_17960  0.021569 
iB03_42_v n1_521_18116 0  0.021569 
iB03_42_g 0 n0_429_18129  0.021569 
iB03_43_v n1_521_18143 0  0.021569 
iB03_43_g 0 n0_429_18129  0.021569 
iB03_44_v n1_521_18176 0  0.021569 
iB03_44_g 0 n0_429_18162  0.021569 
iB03_45_v n1_333_18359 0  0.021569 
iB03_45_g 0 n0_241_18345  0.021569 
iB03_46_v n1_333_18392 0  0.021569 
iB03_46_g 0 n0_241_18378  0.021569 
iB03_47_v n1_333_18527 0  0.021569 
iB03_47_g 0 n0_241_18561  0.021569 
iB03_48_v n1_333_18575 0  0.021569 
iB03_48_g 0 n0_241_18561  0.021569 
iB03_49_v n1_333_18608 0  0.021569 
iB03_49_g 0 n0_241_18594  0.021569 
iB03_50_v n1_380_18392 0  0.021569 
iB03_50_g 0 n0_429_18345  0.021569 
iB03_51_v n1_380_18527 0  0.021569 
iB03_51_g 0 n0_429_18594  0.021569 
iB03_52_v n1_521_18359 0  0.021569 
iB03_52_g 0 n0_429_18345  0.021569 
iB03_53_v n1_521_18392 0  0.021569 
iB03_53_g 0 n0_429_18345  0.021569 
iB03_54_v n1_521_18527 0  0.021569 
iB03_54_g 0 n0_429_18594  0.021569 
iB03_55_v n1_521_18575 0  0.021569 
iB03_55_g 0 n0_429_18594  0.021569 
iB03_56_v n1_521_18608 0  0.021569 
iB03_56_g 0 n0_429_18594  0.021569 
iB03_57_v n1_333_18791 0  0.021569 
iB03_57_g 0 n0_241_18777  0.021569 
iB03_58_v n1_333_18824 0  0.021569 
iB03_58_g 0 n0_241_18810  0.021569 
iB03_59_v n1_333_19007 0  0.021569 
iB03_59_g 0 n0_241_18993  0.021569 
iB03_60_v n1_333_19040 0  0.021569 
iB03_60_g 0 n0_241_19040  0.021569 
iB03_61_v n1_521_18791 0  0.021569 
iB03_61_g 0 n0_429_18777  0.021569 
iB03_62_v n1_521_18824 0  0.021569 
iB03_62_g 0 n0_429_18810  0.021569 
iB03_63_v n1_521_19007 0  0.021569 
iB03_63_g 0 n0_429_18993  0.021569 
iB03_64_v n1_521_19040 0  0.021569 
iB03_64_g 0 n0_429_19040  0.021569 
iB03_65_v n1_333_19196 0  0.021569 
iB03_65_g 0 n0_241_19209  0.021569 
iB03_66_v n1_333_19223 0  0.021569 
iB03_66_g 0 n0_241_19209  0.021569 
iB03_67_v n1_333_19256 0  0.021569 
iB03_67_g 0 n0_241_19256  0.021569 
iB03_68_v n1_333_19412 0  0.021569 
iB03_68_g 0 n0_241_19425  0.021569 
iB03_69_v n1_333_19439 0  0.021569 
iB03_69_g 0 n0_241_19425  0.021569 
iB03_70_v n1_333_19472 0  0.021569 
iB03_70_g 0 n0_241_19472  0.021569 
iB03_71_v n1_521_19196 0  0.021569 
iB03_71_g 0 n0_429_19209  0.021569 
iB03_72_v n1_521_19223 0  0.021569 
iB03_72_g 0 n0_429_19209  0.021569 
iB03_73_v n1_521_19256 0  0.021569 
iB03_73_g 0 n0_429_19256  0.021569 
iB03_74_v n1_521_19412 0  0.021569 
iB03_74_g 0 n0_429_19425  0.021569 
iB03_75_v n1_521_19439 0  0.021569 
iB03_75_g 0 n0_429_19425  0.021569 
iB03_76_v n1_521_19472 0  0.021569 
iB03_76_g 0 n0_429_19472  0.021569 
iB03_77_v n1_333_19871 0  0.021569 
iB03_77_g 0 n0_241_19857  0.021569 
iB03_78_v n1_333_19904 0  0.021569 
iB03_78_g 0 n0_241_19890  0.021569 
iB03_79_v n1_521_19655 0  0.021569 
iB03_79_g 0 n0_429_19641  0.021569 
iB03_80_v n1_521_19688 0  0.021569 
iB03_80_g 0 n0_429_19674  0.021569 
iB03_81_v n1_521_19871 0  0.021569 
iB03_81_g 0 n0_429_19857  0.021569 
iB03_82_v n1_521_19904 0  0.021569 
iB03_82_g 0 n0_429_19890  0.021569 
iB03_83_v n1_333_20087 0  0.021569 
iB03_83_g 0 n0_241_20073  0.021569 
iB03_84_v n1_333_20120 0  0.021569 
iB03_84_g 0 n0_241_20106  0.021569 
iB03_85_v n1_333_20303 0  0.021569 
iB03_85_g 0 n0_241_20289  0.021569 
iB03_86_v n1_333_20336 0  0.021569 
iB03_86_g 0 n0_241_20322  0.021569 
iB03_87_v n1_521_20087 0  0.021569 
iB03_87_g 0 n0_429_20073  0.021569 
iB03_88_v n1_521_20120 0  0.021569 
iB03_88_g 0 n0_429_20106  0.021569 
iB03_89_v n1_521_20303 0  0.021569 
iB03_89_g 0 n0_429_20289  0.021569 
iB03_90_v n1_521_20336 0  0.021569 
iB03_90_g 0 n0_429_20322  0.021569 
iB03_91_v n1_333_20519 0  0.021569 
iB03_91_g 0 n0_241_20505  0.021569 
iB03_92_v n1_333_20552 0  0.021569 
iB03_92_g 0 n0_241_20538  0.021569 
iB03_93_v n1_333_20687 0  0.021569 
iB03_93_g 0 n0_241_20538  0.021569 
iB03_94_v n1_333_20735 0  0.021569 
iB03_94_g 0 n0_241_20538  0.021569 
iB03_95_v n1_333_20768 0  0.021569 
iB03_95_g 0 n0_241_20538  0.021569 
iB03_96_v n1_380_20687 0  0.021569 
iB03_96_g 0 n0_429_20538  0.021569 
iB03_97_v n1_380_20735 0  0.021569 
iB03_97_g 0 n0_429_20538  0.021569 
iB03_98_v n1_380_20768 0  0.021569 
iB03_98_g 0 n0_429_20538  0.021569 
iB03_99_v n1_521_20519 0  0.021569 
iB03_99_g 0 n0_429_20505  0.021569 
iB03_100_v n1_521_20552 0  0.021569 
iB03_100_g 0 n0_429_20538  0.021569 
iB03_101_v n1_521_20687 0  0.021569 
iB03_101_g 0 n0_429_20538  0.021569 
iB03_102_v n1_521_20768 0  0.021569 
iB03_102_g 0 n0_429_20538  0.021569 
iB03_103_v n1_521_20951 0  0.021569 
iB03_103_g 0 n0_429_20538  0.021569 
iB03_104_v n1_521_20984 0  0.021569 
iB03_104_g 0 n0_429_20538  0.021569 
iB03_105_v n1_2400_18527 0  0.021569 
iB03_105_g 0 n0_2491_18378  0.021569 
iB03_106_v n1_2400_18575 0  0.021569 
iB03_106_g 0 n0_2491_18378  0.021569 
iB03_107_v n1_2400_18608 0  0.021569 
iB03_107_g 0 n0_2491_18378  0.021569 
iB03_108_v n1_2400_18791 0  0.021569 
iB03_108_g 0 n0_2491_18378  0.021569 
iB03_109_v n1_2400_18824 0  0.021569 
iB03_109_g 0 n0_2491_18378  0.021569 
iB03_110_v n1_2400_19007 0  0.021569 
iB03_110_g 0 n0_2491_18378  0.021569 
iB03_111_v n1_2400_19040 0  0.021569 
iB03_111_g 0 n0_2491_18378  0.021569 
iB03_112_v n1_2400_19223 0  0.021569 
iB03_112_g 0 n0_1554_19209  0.021569 
iB03_113_v n1_2400_19256 0  0.021569 
iB03_113_g 0 n0_1554_19256  0.021569 
iB03_114_v n1_2400_19439 0  0.021569 
iB03_114_g 0 n0_1554_19425  0.021569 
iB03_115_v n1_2400_19472 0  0.021569 
iB03_115_g 0 n0_1554_19472  0.021569 
iB03_116_v n1_2400_19655 0  0.021569 
iB03_116_g 0 n0_1646_19641  0.021569 
iB03_117_v n1_2400_19688 0  0.021569 
iB03_117_g 0 n0_1646_19674  0.021569 
iB03_118_v n1_2400_19871 0  0.021569 
iB03_118_g 0 n0_1646_19857  0.021569 
iB03_119_v n1_2400_19904 0  0.021569 
iB03_119_g 0 n0_1646_19890  0.021569 
iB03_120_v n1_2400_20087 0  0.021569 
iB03_120_g 0 n0_1646_20073  0.021569 
iB03_121_v n1_2400_20120 0  0.021569 
iB03_121_g 0 n0_1646_20106  0.021569 
iB03_122_v n1_2400_20303 0  0.021569 
iB03_122_g 0 n0_1646_20289  0.021569 
iB03_123_v n1_2400_20336 0  0.021569 
iB03_123_g 0 n0_1646_20322  0.021569 
iB03_124_v n1_2400_20519 0  0.021569 
iB03_124_g 0 n0_1646_20505  0.021569 
iB03_125_v n1_2400_20552 0  0.021569 
iB03_125_g 0 n0_1646_20538  0.021569 
iB03_126_v n1_2400_20687 0  0.021569 
iB03_126_g 0 n0_1646_20754  0.021569 
iB03_127_v n1_2400_20735 0  0.021569 
iB03_127_g 0 n0_1646_20754  0.021569 
iB03_128_v n1_2400_20768 0  0.021569 
iB03_128_g 0 n0_1646_20754  0.021569 
iB03_129_v n1_2400_20951 0  0.021569 
iB03_129_g 0 n0_1646_20937  0.021569 
iB03_130_v n1_2400_20984 0  0.021569 
iB03_130_g 0 n0_1646_20970  0.021569 
iB03_131_v n1_2583_15983 0  0.021569 
iB03_131_g 0 n0_2491_15969  0.021569 
iB03_132_v n1_2583_16016 0  0.021569 
iB03_132_g 0 n0_2491_16002  0.021569 
iB03_133_v n1_2583_16199 0  0.021569 
iB03_133_g 0 n0_2491_16185  0.021569 
iB03_134_v n1_2583_16232 0  0.021569 
iB03_134_g 0 n0_2491_16218  0.021569 
iB03_135_v n1_2630_16199 0  0.021569 
iB03_135_g 0 n0_2491_16185  0.021569 
iB03_136_v n1_2630_16232 0  0.021569 
iB03_136_g 0 n0_2491_16218  0.021569 
iB03_137_v n1_2771_15983 0  0.021569 
iB03_137_g 0 n0_2679_15969  0.021569 
iB03_138_v n1_2771_16016 0  0.021569 
iB03_138_g 0 n0_2679_16002  0.021569 
iB03_139_v n1_2771_16199 0  0.021569 
iB03_139_g 0 n0_2679_16002  0.021569 
iB03_140_v n1_2583_16415 0  0.021569 
iB03_140_g 0 n0_2491_16401  0.021569 
iB03_141_v n1_2583_16448 0  0.021569 
iB03_141_g 0 n0_2491_16434  0.021569 
iB03_142_v n1_2583_16582 0  0.021569 
iB03_142_g 0 n0_2491_16617  0.021569 
iB03_143_v n1_2583_16631 0  0.021569 
iB03_143_g 0 n0_2491_16617  0.021569 
iB03_144_v n1_2583_16664 0  0.021569 
iB03_144_g 0 n0_2491_16664  0.021569 
iB03_145_v n1_2771_16415 0  0.021569 
iB03_145_g 0 n0_2679_16401  0.021569 
iB03_146_v n1_2771_16448 0  0.021569 
iB03_146_g 0 n0_2679_16434  0.021569 
iB03_147_v n1_2771_16582 0  0.021569 
iB03_147_g 0 n0_2679_16617  0.021569 
iB03_148_v n1_2771_16631 0  0.021569 
iB03_148_g 0 n0_2679_16617  0.021569 
iB03_149_v n1_2771_16664 0  0.021569 
iB03_149_g 0 n0_2679_16664  0.021569 
iB03_150_v n1_2583_16798 0  0.021569 
iB03_150_g 0 n0_2491_16833  0.021569 
iB03_151_v n1_2583_16820 0  0.021569 
iB03_151_g 0 n0_2491_16833  0.021569 
iB03_152_v n1_2583_16847 0  0.021569 
iB03_152_g 0 n0_2491_16833  0.021569 
iB03_153_v n1_2583_16880 0  0.021569 
iB03_153_g 0 n0_2491_16880  0.021569 
iB03_154_v n1_2583_17036 0  0.021569 
iB03_154_g 0 n0_2491_17049  0.021569 
iB03_155_v n1_2583_17063 0  0.021569 
iB03_155_g 0 n0_2491_17049  0.021569 
iB03_156_v n1_2583_17096 0  0.021569 
iB03_156_g 0 n0_2491_17082  0.021569 
iB03_157_v n1_2771_16798 0  0.021569 
iB03_157_g 0 n0_2679_16833  0.021569 
iB03_158_v n1_2771_16820 0  0.021569 
iB03_158_g 0 n0_2679_16833  0.021569 
iB03_159_v n1_2771_16847 0  0.021569 
iB03_159_g 0 n0_2679_16833  0.021569 
iB03_160_v n1_2771_16880 0  0.021569 
iB03_160_g 0 n0_2679_16880  0.021569 
iB03_161_v n1_2771_17036 0  0.021569 
iB03_161_g 0 n0_2679_17049  0.021569 
iB03_162_v n1_2771_17063 0  0.021569 
iB03_162_g 0 n0_2679_17049  0.021569 
iB03_163_v n1_2771_17096 0  0.021569 
iB03_163_g 0 n0_2679_17082  0.021569 
iB03_164_v n1_2583_17495 0  0.021569 
iB03_164_g 0 n0_2491_17481  0.021569 
iB03_165_v n1_2771_17279 0  0.021569 
iB03_165_g 0 n0_2679_17265  0.021569 
iB03_166_v n1_2771_17312 0  0.021569 
iB03_166_g 0 n0_2679_17298  0.021569 
iB03_167_v n1_2771_17495 0  0.021569 
iB03_167_g 0 n0_2679_17481  0.021569 
iB03_168_v n1_2583_17528 0  0.021569 
iB03_168_g 0 n0_2491_17528  0.021569 
iB03_169_v n1_2583_17662 0  0.021569 
iB03_169_g 0 n0_2491_17697  0.021569 
iB03_170_v n1_2583_17684 0  0.021569 
iB03_170_g 0 n0_2491_17697  0.021569 
iB03_171_v n1_2583_17711 0  0.021569 
iB03_171_g 0 n0_2491_17697  0.021569 
iB03_172_v n1_2583_17744 0  0.021569 
iB03_172_g 0 n0_2491_17730  0.021569 
iB03_173_v n1_2583_17927 0  0.021569 
iB03_173_g 0 n0_2491_17913  0.021569 
iB03_174_v n1_2771_17528 0  0.021569 
iB03_174_g 0 n0_2679_17528  0.021569 
iB03_175_v n1_2771_17662 0  0.021569 
iB03_175_g 0 n0_2679_17697  0.021569 
iB03_176_v n1_2771_17684 0  0.021569 
iB03_176_g 0 n0_2679_17697  0.021569 
iB03_177_v n1_2771_17711 0  0.021569 
iB03_177_g 0 n0_2679_17697  0.021569 
iB03_178_v n1_2771_17744 0  0.021569 
iB03_178_g 0 n0_2679_17730  0.021569 
iB03_179_v n1_2771_17927 0  0.021569 
iB03_179_g 0 n0_2679_17913  0.021569 
iB03_180_v n1_2583_17960 0  0.021569 
iB03_180_g 0 n0_2491_17960  0.021569 
iB03_181_v n1_2583_18143 0  0.021569 
iB03_181_g 0 n0_2491_18129  0.021569 
iB03_182_v n1_2583_18176 0  0.021569 
iB03_182_g 0 n0_2491_18162  0.021569 
iB03_183_v n1_2771_17960 0  0.021569 
iB03_183_g 0 n0_2679_17960  0.021569 
iB03_184_v n1_2771_18143 0  0.021569 
iB03_184_g 0 n0_2679_18129  0.021569 
iB03_185_v n1_2771_18176 0  0.021569 
iB03_185_g 0 n0_2679_18162  0.021569 
iB03_186_v n1_2583_18359 0  0.021569 
iB03_186_g 0 n0_2491_18345  0.021569 
iB03_187_v n1_2583_18392 0  0.021569 
iB03_187_g 0 n0_2491_18378  0.021569 
iB03_188_v n1_2583_18527 0  0.021569 
iB03_188_g 0 n0_2491_18378  0.021569 
iB03_189_v n1_2583_18575 0  0.021569 
iB03_189_g 0 n0_2491_18378  0.021569 
iB03_190_v n1_2583_18608 0  0.021569 
iB03_190_g 0 n0_2491_18378  0.021569 
iB03_191_v n1_2630_18392 0  0.021569 
iB03_191_g 0 n0_2679_18345  0.021569 
iB03_192_v n1_2630_18527 0  0.021569 
iB03_192_g 0 n0_2679_18345  0.021569 
iB03_193_v n1_2771_18359 0  0.021569 
iB03_193_g 0 n0_2679_18345  0.021569 
iB03_194_v n1_2771_18392 0  0.021569 
iB03_194_g 0 n0_2679_18345  0.021569 
iB03_195_v n1_2771_18527 0  0.021569 
iB03_195_g 0 n0_2679_18345  0.021569 
iB03_196_v n1_2771_18575 0  0.021569 
iB03_196_g 0 n0_2679_18345  0.021569 
iB03_197_v n1_2771_18608 0  0.021569 
iB03_197_g 0 n0_2679_18345  0.021569 
iB03_198_v n1_2864_18527 0  0.021569 
iB03_198_g 0 n0_2679_18345  0.021569 
iB03_199_v n1_2864_18575 0  0.021569 
iB03_199_g 0 n0_2679_18345  0.021569 
iB03_200_v n1_2864_18608 0  0.021569 
iB03_200_g 0 n0_2679_18345  0.021569 
iB03_201_v n1_2583_18791 0  0.021569 
iB03_201_g 0 n0_2491_18378  0.021569 
iB03_202_v n1_2583_18824 0  0.021569 
iB03_202_g 0 n0_2491_18378  0.021569 
iB03_203_v n1_2583_19007 0  0.021569 
iB03_203_g 0 n0_2491_18378  0.021569 
iB03_204_v n1_2583_19040 0  0.021569 
iB03_204_g 0 n0_2491_18378  0.021569 
iB03_205_v n1_2771_18791 0  0.021569 
iB03_205_g 0 n0_2679_18345  0.021569 
iB03_206_v n1_2771_18824 0  0.021569 
iB03_206_g 0 n0_2679_18345  0.021569 
iB03_207_v n1_2771_19007 0  0.021569 
iB03_207_g 0 n0_2679_18345  0.021569 
iB03_208_v n1_2771_19040 0  0.021569 
iB03_208_g 0 n0_2679_18345  0.021569 
iB03_209_v n1_2864_18791 0  0.021569 
iB03_209_g 0 n0_2679_18345  0.021569 
iB03_210_v n1_2864_18824 0  0.021569 
iB03_210_g 0 n0_2679_18345  0.021569 
iB03_211_v n1_2864_19007 0  0.021569 
iB03_211_g 0 n0_2679_18345  0.021569 
iB03_212_v n1_2864_19040 0  0.021569 
iB03_212_g 0 n0_2679_18345  0.021569 
iB03_213_v n1_2583_19223 0  0.021569 
iB03_213_g 0 n0_2491_18378  0.021569 
iB03_214_v n1_2583_19256 0  0.021569 
iB03_214_g 0 n0_2491_18378  0.021569 
iB03_215_v n1_2583_19439 0  0.021569 
iB03_215_g 0 n0_1554_19425  0.021569 
iB03_216_v n1_2583_19472 0  0.021569 
iB03_216_g 0 n0_1554_19472  0.021569 
iB03_217_v n1_2771_19223 0  0.021569 
iB03_217_g 0 n0_3616_19209  0.021569 
iB03_218_v n1_2771_19256 0  0.021569 
iB03_218_g 0 n0_3616_19242  0.021569 
iB03_219_v n1_2771_19439 0  0.021569 
iB03_219_g 0 n0_3616_19425  0.021569 
iB03_220_v n1_2771_19472 0  0.021569 
iB03_220_g 0 n0_3616_19458  0.021569 
iB03_221_v n1_2864_19223 0  0.021569 
iB03_221_g 0 n0_3616_19209  0.021569 
iB03_222_v n1_2864_19256 0  0.021569 
iB03_222_g 0 n0_3616_19242  0.021569 
iB03_223_v n1_2864_19439 0  0.021569 
iB03_223_g 0 n0_3616_19425  0.021569 
iB03_224_v n1_2864_19472 0  0.021569 
iB03_224_g 0 n0_3616_19458  0.021569 
iB03_225_v n1_2583_19871 0  0.021569 
iB03_225_g 0 n0_1646_19857  0.021569 
iB03_226_v n1_2583_19904 0  0.021569 
iB03_226_g 0 n0_1646_19890  0.021569 
iB03_227_v n1_2771_19655 0  0.021569 
iB03_227_g 0 n0_3616_19641  0.021569 
iB03_228_v n1_2771_19688 0  0.021569 
iB03_228_g 0 n0_3616_19674  0.021569 
iB03_229_v n1_2771_19871 0  0.021569 
iB03_229_g 0 n0_3616_19857  0.021569 
iB03_230_v n1_2771_19904 0  0.021569 
iB03_230_g 0 n0_3616_19890  0.021569 
iB03_231_v n1_2864_19655 0  0.021569 
iB03_231_g 0 n0_3616_19641  0.021569 
iB03_232_v n1_2864_19688 0  0.021569 
iB03_232_g 0 n0_3616_19674  0.021569 
iB03_233_v n1_2864_19871 0  0.021569 
iB03_233_g 0 n0_3616_19857  0.021569 
iB03_234_v n1_2864_19904 0  0.021569 
iB03_234_g 0 n0_3616_19890  0.021569 
iB03_235_v n1_2583_20087 0  0.021569 
iB03_235_g 0 n0_1646_20073  0.021569 
iB03_236_v n1_2583_20120 0  0.021569 
iB03_236_g 0 n0_1646_20106  0.021569 
iB03_237_v n1_2583_20303 0  0.021569 
iB03_237_g 0 n0_1646_20289  0.021569 
iB03_238_v n1_2583_20336 0  0.021569 
iB03_238_g 0 n0_1646_20322  0.021569 
iB03_239_v n1_2771_20087 0  0.021569 
iB03_239_g 0 n0_3616_20073  0.021569 
iB03_240_v n1_2771_20120 0  0.021569 
iB03_240_g 0 n0_3616_20106  0.021569 
iB03_241_v n1_2771_20303 0  0.021569 
iB03_241_g 0 n0_3616_20289  0.021569 
iB03_242_v n1_2771_20336 0  0.021569 
iB03_242_g 0 n0_3616_20322  0.021569 
iB03_243_v n1_2864_20087 0  0.021569 
iB03_243_g 0 n0_3616_20073  0.021569 
iB03_244_v n1_2864_20120 0  0.021569 
iB03_244_g 0 n0_3616_20106  0.021569 
iB03_245_v n1_2864_20303 0  0.021569 
iB03_245_g 0 n0_3616_20289  0.021569 
iB03_246_v n1_2864_20336 0  0.021569 
iB03_246_g 0 n0_3616_20322  0.021569 
iB03_247_v n1_2583_20519 0  0.021569 
iB03_247_g 0 n0_1646_20505  0.021569 
iB03_248_v n1_2583_20552 0  0.021569 
iB03_248_g 0 n0_1646_20538  0.021569 
iB03_249_v n1_2583_20687 0  0.021569 
iB03_249_g 0 n0_1646_20754  0.021569 
iB03_250_v n1_2583_20735 0  0.021569 
iB03_250_g 0 n0_1646_20754  0.021569 
iB03_251_v n1_2583_20768 0  0.021569 
iB03_251_g 0 n0_1646_20754  0.021569 
iB03_252_v n1_2630_20687 0  0.021569 
iB03_252_g 0 n0_3616_20754  0.021569 
iB03_253_v n1_2630_20735 0  0.021569 
iB03_253_g 0 n0_3616_20754  0.021569 
iB03_254_v n1_2630_20768 0  0.021569 
iB03_254_g 0 n0_3616_20754  0.021569 
iB03_255_v n1_2771_20519 0  0.021569 
iB03_255_g 0 n0_3616_20505  0.021569 
iB03_256_v n1_2771_20552 0  0.021569 
iB03_256_g 0 n0_3616_20538  0.021569 
iB03_257_v n1_2771_20687 0  0.021569 
iB03_257_g 0 n0_3616_20754  0.021569 
iB03_258_v n1_2771_20768 0  0.021569 
iB03_258_g 0 n0_3616_20754  0.021569 
iB03_259_v n1_2864_20519 0  0.021569 
iB03_259_g 0 n0_3616_20505  0.021569 
iB03_260_v n1_2864_20552 0  0.021569 
iB03_260_g 0 n0_3616_20538  0.021569 
iB03_261_v n1_2864_20687 0  0.021569 
iB03_261_g 0 n0_3616_20754  0.021569 
iB03_262_v n1_2864_20735 0  0.021569 
iB03_262_g 0 n0_3616_20754  0.021569 
iB03_263_v n1_2864_20768 0  0.021569 
iB03_263_g 0 n0_3616_20754  0.021569 
iB03_264_v n1_2583_20951 0  0.021569 
iB03_264_g 0 n0_1646_20937  0.021569 
iB03_265_v n1_2583_20984 0  0.021569 
iB03_265_g 0 n0_1646_20970  0.021569 
iB03_266_v n1_2771_20951 0  0.021569 
iB03_266_g 0 n0_3616_20937  0.021569 
iB03_267_v n1_2771_20984 0  0.021569 
iB03_267_g 0 n0_3616_20970  0.021569 
iB03_268_v n1_2864_20951 0  0.021569 
iB03_268_g 0 n0_3616_20937  0.021569 
iB03_269_v n1_2864_20984 0  0.021569 
iB03_269_g 0 n0_3616_20970  0.021569 
iB03_270_v n1_4833_15983 0  0.021569 
iB03_270_g 0 n0_4741_15969  0.021569 
iB03_271_v n1_4833_16016 0  0.021569 
iB03_271_g 0 n0_4741_16016  0.021569 
iB03_272_v n1_4833_16172 0  0.021569 
iB03_272_g 0 n0_4741_16185  0.021569 
iB03_273_v n1_4833_16199 0  0.021569 
iB03_273_g 0 n0_4741_16185  0.021569 
iB03_274_v n1_4833_16232 0  0.021569 
iB03_274_g 0 n0_4741_16185  0.021569 
iB03_275_v n1_4880_16172 0  0.021569 
iB03_275_g 0 n0_4741_16185  0.021569 
iB03_276_v n1_4880_16199 0  0.021569 
iB03_276_g 0 n0_4741_16185  0.021569 
iB03_277_v n1_4880_16232 0  0.021569 
iB03_277_g 0 n0_4741_16185  0.021569 
iB03_278_v n1_4833_16415 0  0.021569 
iB03_278_g 0 n0_4741_16185  0.021569 
iB03_279_v n1_4833_16448 0  0.021569 
iB03_279_g 0 n0_4741_16185  0.021569 
iB03_280_v n1_4833_16631 0  0.021569 
iB03_280_g 0 n0_4741_16185  0.021569 
iB03_281_v n1_4833_16664 0  0.021569 
iB03_281_g 0 n0_4741_16185  0.021569 
iB03_282_v n1_4833_16847 0  0.021569 
iB03_282_g 0 n0_4741_16185  0.021569 
iB03_283_v n1_4833_16880 0  0.021569 
iB03_283_g 0 n0_4741_16185  0.021569 
iB03_284_v n1_4833_17036 0  0.021569 
iB03_284_g 0 n0_4741_16185  0.021569 
iB03_285_v n1_4833_17063 0  0.021569 
iB03_285_g 0 n0_4741_16185  0.021569 
iB03_286_v n1_4833_17096 0  0.021569 
iB03_286_g 0 n0_4741_16185  0.021569 
iB03_287_v n1_4833_17468 0  0.021569 
iB03_287_g 0 n0_3896_17481  0.021569 
iB03_288_v n1_4833_17495 0  0.021569 
iB03_288_g 0 n0_3896_17481  0.021569 
iB03_289_v n1_4833_17528 0  0.021569 
iB03_289_g 0 n0_3896_17528  0.021569 
iB03_290_v n1_4833_17684 0  0.021569 
iB03_290_g 0 n0_3896_17697  0.021569 
iB03_291_v n1_4833_17711 0  0.021569 
iB03_291_g 0 n0_3896_17697  0.021569 
iB03_292_v n1_4833_17744 0  0.021569 
iB03_292_g 0 n0_3896_17730  0.021569 
iB03_293_v n1_4833_17927 0  0.021569 
iB03_293_g 0 n0_3896_17913  0.021569 
iB03_294_v n1_4833_17960 0  0.021569 
iB03_294_g 0 n0_3896_17946  0.021569 
iB03_295_v n1_4833_18143 0  0.021569 
iB03_295_g 0 n0_3896_18129  0.021569 
iB03_296_v n1_4833_18176 0  0.021569 
iB03_296_g 0 n0_3896_18162  0.021569 
iB03_297_v n1_4650_18527 0  0.021569 
iB03_297_g 0 n0_3896_18561  0.021569 
iB03_298_v n1_4650_18575 0  0.021569 
iB03_298_g 0 n0_3896_18561  0.021569 
iB03_299_v n1_4650_18608 0  0.021569 
iB03_299_g 0 n0_3896_18594  0.021569 
iB03_300_v n1_4833_18359 0  0.021569 
iB03_300_g 0 n0_3896_18345  0.021569 
iB03_301_v n1_4833_18392 0  0.021569 
iB03_301_g 0 n0_3896_18378  0.021569 
iB03_302_v n1_4833_18527 0  0.021569 
iB03_302_g 0 n0_3896_18561  0.021569 
iB03_303_v n1_4833_18548 0  0.021569 
iB03_303_g 0 n0_3896_18561  0.021569 
iB03_304_v n1_4833_18575 0  0.021569 
iB03_304_g 0 n0_3896_18561  0.021569 
iB03_305_v n1_4833_18608 0  0.021569 
iB03_305_g 0 n0_3896_18594  0.021569 
iB03_306_v n1_4880_18392 0  0.021569 
iB03_306_g 0 n0_5866_18392  0.021569 
iB03_307_v n1_4880_18527 0  0.021569 
iB03_307_g 0 n0_3896_18561  0.021569 
iB03_308_v n1_4880_18548 0  0.021569 
iB03_308_g 0 n0_3896_18561  0.021569 
iB03_309_v n1_4650_18791 0  0.021569 
iB03_309_g 0 n0_3896_18777  0.021569 
iB03_310_v n1_4650_18824 0  0.021569 
iB03_310_g 0 n0_3896_18810  0.021569 
iB03_311_v n1_4650_19007 0  0.021569 
iB03_311_g 0 n0_3896_18993  0.021569 
iB03_312_v n1_4650_19040 0  0.021569 
iB03_312_g 0 n0_3896_19026  0.021569 
iB03_313_v n1_4833_18764 0  0.021569 
iB03_313_g 0 n0_3896_18777  0.021569 
iB03_314_v n1_4833_18791 0  0.021569 
iB03_314_g 0 n0_3896_18777  0.021569 
iB03_315_v n1_4833_18824 0  0.021569 
iB03_315_g 0 n0_3896_18810  0.021569 
iB03_316_v n1_4833_18980 0  0.021569 
iB03_316_g 0 n0_3896_18993  0.021569 
iB03_317_v n1_4833_19007 0  0.021569 
iB03_317_g 0 n0_3896_18993  0.021569 
iB03_318_v n1_4833_19040 0  0.021569 
iB03_318_g 0 n0_3896_19026  0.021569 
iB03_319_v n1_4650_19223 0  0.021569 
iB03_319_g 0 n0_3896_19209  0.021569 
iB03_320_v n1_4650_19256 0  0.021569 
iB03_320_g 0 n0_3896_19242  0.021569 
iB03_321_v n1_4650_19439 0  0.021569 
iB03_321_g 0 n0_3896_19425  0.021569 
iB03_322_v n1_4650_19472 0  0.021569 
iB03_322_g 0 n0_3896_19458  0.021569 
iB03_323_v n1_4833_19196 0  0.021569 
iB03_323_g 0 n0_3896_19209  0.021569 
iB03_324_v n1_4833_19223 0  0.021569 
iB03_324_g 0 n0_3896_19209  0.021569 
iB03_325_v n1_4833_19256 0  0.021569 
iB03_325_g 0 n0_3896_19242  0.021569 
iB03_326_v n1_4833_19439 0  0.021569 
iB03_326_g 0 n0_3896_19425  0.021569 
iB03_327_v n1_4833_19472 0  0.021569 
iB03_327_g 0 n0_3896_19458  0.021569 
iB03_328_v n1_4650_19655 0  0.021569 
iB03_328_g 0 n0_3896_19641  0.021569 
iB03_329_v n1_4650_19688 0  0.021569 
iB03_329_g 0 n0_3896_19674  0.021569 
iB03_330_v n1_4650_19871 0  0.021569 
iB03_330_g 0 n0_3896_19857  0.021569 
iB03_331_v n1_4650_19904 0  0.021569 
iB03_331_g 0 n0_3896_19890  0.021569 
iB03_332_v n1_4833_19871 0  0.021569 
iB03_332_g 0 n0_3896_19857  0.021569 
iB03_333_v n1_4833_19904 0  0.021569 
iB03_333_g 0 n0_3896_19890  0.021569 
iB03_334_v n1_4650_20087 0  0.021569 
iB03_334_g 0 n0_3896_20073  0.021569 
iB03_335_v n1_4650_20120 0  0.021569 
iB03_335_g 0 n0_3896_20106  0.021569 
iB03_336_v n1_4650_20303 0  0.021569 
iB03_336_g 0 n0_3896_20289  0.021569 
iB03_337_v n1_4650_20336 0  0.021569 
iB03_337_g 0 n0_3896_20322  0.021569 
iB03_338_v n1_4833_20087 0  0.021569 
iB03_338_g 0 n0_3896_20073  0.021569 
iB03_339_v n1_4833_20120 0  0.021569 
iB03_339_g 0 n0_3896_20106  0.021569 
iB03_340_v n1_4833_20303 0  0.021569 
iB03_340_g 0 n0_3896_20289  0.021569 
iB03_341_v n1_4833_20336 0  0.021569 
iB03_341_g 0 n0_3896_20322  0.021569 
iB03_342_v n1_4650_20519 0  0.021569 
iB03_342_g 0 n0_3896_20505  0.021569 
iB03_343_v n1_4650_20552 0  0.021569 
iB03_343_g 0 n0_3896_20538  0.021569 
iB03_344_v n1_4650_20687 0  0.021569 
iB03_344_g 0 n0_3896_20754  0.021569 
iB03_345_v n1_4650_20735 0  0.021569 
iB03_345_g 0 n0_3896_20754  0.021569 
iB03_346_v n1_4650_20768 0  0.021569 
iB03_346_g 0 n0_3896_20754  0.021569 
iB03_347_v n1_4833_20519 0  0.021569 
iB03_347_g 0 n0_3896_20505  0.021569 
iB03_348_v n1_4833_20552 0  0.021569 
iB03_348_g 0 n0_3896_20538  0.021569 
iB03_349_v n1_4833_20687 0  0.021569 
iB03_349_g 0 n0_3896_20754  0.021569 
iB03_350_v n1_4833_20735 0  0.021569 
iB03_350_g 0 n0_3896_20754  0.021569 
iB03_351_v n1_4833_20768 0  0.021569 
iB03_351_g 0 n0_3896_20754  0.021569 
iB03_352_v n1_4880_20687 0  0.021569 
iB03_352_g 0 n0_3896_20754  0.021569 
iB03_353_v n1_4880_20735 0  0.021569 
iB03_353_g 0 n0_3896_20754  0.021569 
iB03_354_v n1_4880_20768 0  0.021569 
iB03_354_g 0 n0_3896_20754  0.021569 
iB03_355_v n1_4650_20951 0  0.021569 
iB03_355_g 0 n0_3896_20937  0.021569 
iB03_356_v n1_4650_20984 0  0.021569 
iB03_356_g 0 n0_3896_20970  0.021569 
iB03_357_v n1_4833_20951 0  0.021569 
iB03_357_g 0 n0_3896_20937  0.021569 
iB03_358_v n1_4833_20984 0  0.021569 
iB03_358_g 0 n0_3896_20970  0.021569 
iB03_359_v n1_5021_15983 0  0.021569 
iB03_359_g 0 n0_4929_15969  0.021569 
iB03_360_v n1_5021_16016 0  0.021569 
iB03_360_g 0 n0_4929_16016  0.021569 
iB03_361_v n1_5021_16172 0  0.021569 
iB03_361_g 0 n0_4929_16016  0.021569 
iB03_362_v n1_5021_16199 0  0.021569 
iB03_362_g 0 n0_4929_16016  0.021569 
iB03_363_v n1_5021_16415 0  0.021569 
iB03_363_g 0 n0_4741_16185  0.021569 
iB03_364_v n1_5021_16448 0  0.021569 
iB03_364_g 0 n0_4741_16185  0.021569 
iB03_365_v n1_5021_16631 0  0.021569 
iB03_365_g 0 n0_4741_16185  0.021569 
iB03_366_v n1_5021_16664 0  0.021569 
iB03_366_g 0 n0_4741_16185  0.021569 
iB03_367_v n1_5021_16847 0  0.021569 
iB03_367_g 0 n0_4741_16185  0.021569 
iB03_368_v n1_5021_16880 0  0.021569 
iB03_368_g 0 n0_4741_16185  0.021569 
iB03_369_v n1_5021_17036 0  0.021569 
iB03_369_g 0 n0_5866_17049  0.021569 
iB03_370_v n1_5021_17063 0  0.021569 
iB03_370_g 0 n0_5866_17049  0.021569 
iB03_371_v n1_5021_17096 0  0.021569 
iB03_371_g 0 n0_5866_17096  0.021569 
iB03_372_v n1_5021_17252 0  0.021569 
iB03_372_g 0 n0_5866_17265  0.021569 
iB03_373_v n1_5021_17279 0  0.021569 
iB03_373_g 0 n0_5866_17265  0.021569 
iB03_374_v n1_5021_17312 0  0.021569 
iB03_374_g 0 n0_5866_17312  0.021569 
iB03_375_v n1_5021_17446 0  0.021569 
iB03_375_g 0 n0_5866_17481  0.021569 
iB03_376_v n1_5021_17468 0  0.021569 
iB03_376_g 0 n0_5866_17481  0.021569 
iB03_377_v n1_5021_17495 0  0.021569 
iB03_377_g 0 n0_5866_17481  0.021569 
iB03_378_v n1_5021_17528 0  0.021569 
iB03_378_g 0 n0_5866_17528  0.021569 
iB03_379_v n1_5021_17684 0  0.021569 
iB03_379_g 0 n0_5866_17697  0.021569 
iB03_380_v n1_5021_17711 0  0.021569 
iB03_380_g 0 n0_5866_17697  0.021569 
iB03_381_v n1_5021_17744 0  0.021569 
iB03_381_g 0 n0_5866_17730  0.021569 
iB03_382_v n1_5021_17927 0  0.021569 
iB03_382_g 0 n0_5866_17913  0.021569 
iB03_383_v n1_5021_17960 0  0.021569 
iB03_383_g 0 n0_5866_17946  0.021569 
iB03_384_v n1_5021_18143 0  0.021569 
iB03_384_g 0 n0_5866_18129  0.021569 
iB03_385_v n1_5021_18176 0  0.021569 
iB03_385_g 0 n0_5866_18162  0.021569 
iB03_386_v n1_5021_18359 0  0.021569 
iB03_386_g 0 n0_5866_18345  0.021569 
iB03_387_v n1_5021_18392 0  0.021569 
iB03_387_g 0 n0_5866_18392  0.021569 
iB03_388_v n1_5021_18527 0  0.021569 
iB03_388_g 0 n0_5866_18561  0.021569 
iB03_389_v n1_5021_18548 0  0.021569 
iB03_389_g 0 n0_5866_18561  0.021569 
iB03_390_v n1_5021_18575 0  0.021569 
iB03_390_g 0 n0_5866_18561  0.021569 
iB03_391_v n1_5021_18608 0  0.021569 
iB03_391_g 0 n0_5866_18608  0.021569 
iB03_392_v n1_5114_18527 0  0.021569 
iB03_392_g 0 n0_5866_18561  0.021569 
iB03_393_v n1_5114_18548 0  0.021569 
iB03_393_g 0 n0_5866_18561  0.021569 
iB03_394_v n1_5114_18575 0  0.021569 
iB03_394_g 0 n0_5866_18561  0.021569 
iB03_395_v n1_5114_18608 0  0.021569 
iB03_395_g 0 n0_5866_18608  0.021569 
iB03_396_v n1_5021_18764 0  0.021569 
iB03_396_g 0 n0_5866_18777  0.021569 
iB03_397_v n1_5021_18791 0  0.021569 
iB03_397_g 0 n0_5866_18777  0.021569 
iB03_398_v n1_5021_18824 0  0.021569 
iB03_398_g 0 n0_5866_18824  0.021569 
iB03_399_v n1_5021_18980 0  0.021569 
iB03_399_g 0 n0_5866_18993  0.021569 
iB03_400_v n1_5021_19007 0  0.021569 
iB03_400_g 0 n0_5866_18993  0.021569 
iB03_401_v n1_5021_19040 0  0.021569 
iB03_401_g 0 n0_5866_19040  0.021569 
iB03_402_v n1_5114_18764 0  0.021569 
iB03_402_g 0 n0_5866_18777  0.021569 
iB03_403_v n1_5114_18791 0  0.021569 
iB03_403_g 0 n0_5866_18777  0.021569 
iB03_404_v n1_5114_18824 0  0.021569 
iB03_404_g 0 n0_5866_18824  0.021569 
iB03_405_v n1_5114_18980 0  0.021569 
iB03_405_g 0 n0_5866_18993  0.021569 
iB03_406_v n1_5114_19007 0  0.021569 
iB03_406_g 0 n0_5866_18993  0.021569 
iB03_407_v n1_5114_19040 0  0.021569 
iB03_407_g 0 n0_5866_19040  0.021569 
iB03_408_v n1_5021_19196 0  0.021569 
iB03_408_g 0 n0_5866_19209  0.021569 
iB03_409_v n1_5021_19223 0  0.021569 
iB03_409_g 0 n0_5866_19209  0.021569 
iB03_410_v n1_5021_19256 0  0.021569 
iB03_410_g 0 n0_5866_19242  0.021569 
iB03_411_v n1_5021_19439 0  0.021569 
iB03_411_g 0 n0_5866_19425  0.021569 
iB03_412_v n1_5021_19472 0  0.021569 
iB03_412_g 0 n0_5866_19472  0.021569 
iB03_413_v n1_5114_19196 0  0.021569 
iB03_413_g 0 n0_5866_19209  0.021569 
iB03_414_v n1_5114_19223 0  0.021569 
iB03_414_g 0 n0_5866_19209  0.021569 
iB03_415_v n1_5114_19256 0  0.021569 
iB03_415_g 0 n0_5866_19242  0.021569 
iB03_416_v n1_5114_19439 0  0.021569 
iB03_416_g 0 n0_5866_19425  0.021569 
iB03_417_v n1_5114_19472 0  0.021569 
iB03_417_g 0 n0_5866_19472  0.021569 
iB03_418_v n1_5021_19628 0  0.021569 
iB03_418_g 0 n0_5866_19641  0.021569 
iB03_419_v n1_5021_19655 0  0.021569 
iB03_419_g 0 n0_5866_19641  0.021569 
iB03_420_v n1_5021_19688 0  0.021569 
iB03_420_g 0 n0_5866_19674  0.021569 
iB03_421_v n1_5021_19871 0  0.021569 
iB03_421_g 0 n0_5866_19857  0.021569 
iB03_422_v n1_5021_19904 0  0.021569 
iB03_422_g 0 n0_5866_19890  0.021569 
iB03_423_v n1_5114_19628 0  0.021569 
iB03_423_g 0 n0_5866_19641  0.021569 
iB03_424_v n1_5114_19655 0  0.021569 
iB03_424_g 0 n0_5866_19641  0.021569 
iB03_425_v n1_5114_19688 0  0.021569 
iB03_425_g 0 n0_5866_19674  0.021569 
iB03_426_v n1_5114_19871 0  0.021569 
iB03_426_g 0 n0_5866_19857  0.021569 
iB03_427_v n1_5114_19904 0  0.021569 
iB03_427_g 0 n0_5866_19890  0.021569 
iB03_428_v n1_5021_20087 0  0.021569 
iB03_428_g 0 n0_5866_20073  0.021569 
iB03_429_v n1_5021_20120 0  0.021569 
iB03_429_g 0 n0_5866_20106  0.021569 
iB03_430_v n1_5021_20303 0  0.021569 
iB03_430_g 0 n0_5866_20289  0.021569 
iB03_431_v n1_5021_20336 0  0.021569 
iB03_431_g 0 n0_5866_20322  0.021569 
iB03_432_v n1_5114_20087 0  0.021569 
iB03_432_g 0 n0_5866_20073  0.021569 
iB03_433_v n1_5114_20120 0  0.021569 
iB03_433_g 0 n0_5866_20106  0.021569 
iB03_434_v n1_5114_20303 0  0.021569 
iB03_434_g 0 n0_5866_20289  0.021569 
iB03_435_v n1_5114_20336 0  0.021569 
iB03_435_g 0 n0_5866_20322  0.021569 
iB03_436_v n1_5021_20519 0  0.021569 
iB03_436_g 0 n0_5866_20505  0.021569 
iB03_437_v n1_5021_20552 0  0.021569 
iB03_437_g 0 n0_5866_20538  0.021569 
iB03_438_v n1_5021_20687 0  0.021569 
iB03_438_g 0 n0_5866_20754  0.021569 
iB03_439_v n1_5021_20768 0  0.021569 
iB03_439_g 0 n0_5866_20754  0.021569 
iB03_440_v n1_5114_20519 0  0.021569 
iB03_440_g 0 n0_5866_20505  0.021569 
iB03_441_v n1_5114_20552 0  0.021569 
iB03_441_g 0 n0_5866_20538  0.021569 
iB03_442_v n1_5114_20687 0  0.021569 
iB03_442_g 0 n0_5866_20754  0.021569 
iB03_443_v n1_5114_20735 0  0.021569 
iB03_443_g 0 n0_5866_20754  0.021569 
iB03_444_v n1_5114_20768 0  0.021569 
iB03_444_g 0 n0_5866_20754  0.021569 
iB03_445_v n1_5021_20951 0  0.021569 
iB03_445_g 0 n0_5866_20937  0.021569 
iB03_446_v n1_5021_20984 0  0.021569 
iB03_446_g 0 n0_5866_20970  0.021569 
iB03_447_v n1_5114_20951 0  0.021569 
iB03_447_g 0 n0_5866_20937  0.021569 
iB03_448_v n1_5114_20984 0  0.021569 
iB03_448_g 0 n0_5866_20970  0.021569 
iB21_0_v n1_11583_5350 0  0.0413994 
iB21_0_g 0 n0_10646_5385  0.0413994 
iB21_1_v n1_11583_5399 0  0.0413994 
iB21_1_g 0 n0_10646_5385  0.0413994 
iB21_2_v n1_11583_5432 0  0.0413994 
iB21_2_g 0 n0_10646_5432  0.0413994 
iB21_3_v n1_11583_5566 0  0.0413994 
iB21_3_g 0 n0_10646_5601  0.0413994 
iB21_4_v n1_11583_5615 0  0.0413994 
iB21_4_g 0 n0_10646_5601  0.0413994 
iB21_5_v n1_11583_5648 0  0.0413994 
iB21_5_g 0 n0_10646_5634  0.0413994 
iB21_6_v n1_11583_5782 0  0.0413994 
iB21_6_g 0 n0_10646_5817  0.0413994 
iB21_7_v n1_11583_5831 0  0.0413994 
iB21_7_g 0 n0_10646_5817  0.0413994 
iB21_8_v n1_11583_5864 0  0.0413994 
iB21_8_g 0 n0_10646_5850  0.0413994 
iB21_9_v n1_11583_6263 0  0.0413994 
iB21_9_g 0 n0_10646_6249  0.0413994 
iB21_10_v n1_11583_6296 0  0.0413994 
iB21_10_g 0 n0_10646_6282  0.0413994 
iB21_11_v n1_11583_6430 0  0.0413994 
iB21_11_g 0 n0_10646_6465  0.0413994 
iB21_12_v n1_11583_6479 0  0.0413994 
iB21_12_g 0 n0_10646_6465  0.0413994 
iB21_13_v n1_11583_6512 0  0.0413994 
iB21_13_g 0 n0_10646_6512  0.0413994 
iB21_14_v n1_11583_6646 0  0.0413994 
iB21_14_g 0 n0_10646_6681  0.0413994 
iB21_15_v n1_11583_6695 0  0.0413994 
iB21_15_g 0 n0_10646_6681  0.0413994 
iB21_16_v n1_11583_6728 0  0.0413994 
iB21_16_g 0 n0_10646_6714  0.0413994 
iB21_17_v n1_11583_6862 0  0.0413994 
iB21_17_g 0 n0_10646_6897  0.0413994 
iB21_18_v n1_11583_6911 0  0.0413994 
iB21_18_g 0 n0_10646_6897  0.0413994 
iB21_19_v n1_11583_6944 0  0.0413994 
iB21_19_g 0 n0_10646_6944  0.0413994 
iB21_20_v n1_11583_7078 0  0.0413994 
iB21_20_g 0 n0_10646_7113  0.0413994 
iB21_21_v n1_11583_7127 0  0.0413994 
iB21_21_g 0 n0_10646_7113  0.0413994 
iB21_22_v n1_11583_7160 0  0.0413994 
iB21_22_g 0 n0_10646_7160  0.0413994 
iB21_23_v n1_11583_7294 0  0.0413994 
iB21_23_g 0 n0_10646_7329  0.0413994 
iB21_24_v n1_11630_7160 0  0.0413994 
iB21_24_g 0 n0_10646_7160  0.0413994 
iB21_25_v n1_11630_7294 0  0.0413994 
iB21_25_g 0 n0_10646_7329  0.0413994 
iB21_26_v n1_11583_7343 0  0.0413994 
iB21_26_g 0 n0_10646_7329  0.0413994 
iB21_27_v n1_11583_7376 0  0.0413994 
iB21_27_g 0 n0_10646_7376  0.0413994 
iB21_28_v n1_11583_7510 0  0.0413994 
iB21_28_g 0 n0_10646_7545  0.0413994 
iB21_29_v n1_11583_7559 0  0.0413994 
iB21_29_g 0 n0_10646_7545  0.0413994 
iB21_30_v n1_11583_7592 0  0.0413994 
iB21_30_g 0 n0_10646_7578  0.0413994 
iB21_31_v n1_11583_7775 0  0.0413994 
iB21_31_g 0 n0_10646_7761  0.0413994 
iB21_32_v n1_11583_7808 0  0.0413994 
iB21_32_g 0 n0_10646_7794  0.0413994 
iB21_33_v n1_11583_7991 0  0.0413994 
iB21_33_g 0 n0_10646_7977  0.0413994 
iB21_34_v n1_11583_8024 0  0.0413994 
iB21_34_g 0 n0_10646_8010  0.0413994 
iB21_35_v n1_11583_8207 0  0.0413994 
iB21_35_g 0 n0_10646_8193  0.0413994 
iB21_36_v n1_11583_8240 0  0.0413994 
iB21_36_g 0 n0_10646_8226  0.0413994 
iB21_37_v n1_11583_8456 0  0.0413994 
iB21_37_g 0 n0_10646_8442  0.0413994 
iB21_38_v n1_11583_8639 0  0.0413994 
iB21_38_g 0 n0_11491_9489  0.0413994 
iB21_39_v n1_11583_8672 0  0.0413994 
iB21_39_g 0 n0_11491_9489  0.0413994 
iB21_40_v n1_11583_8855 0  0.0413994 
iB21_40_g 0 n0_11491_9489  0.0413994 
iB21_41_v n1_11583_8888 0  0.0413994 
iB21_41_g 0 n0_11491_9489  0.0413994 
iB21_42_v n1_11583_9071 0  0.0413994 
iB21_42_g 0 n0_11491_9489  0.0413994 
iB21_43_v n1_11583_9104 0  0.0413994 
iB21_43_g 0 n0_11491_9489  0.0413994 
iB21_44_v n1_11583_9287 0  0.0413994 
iB21_44_g 0 n0_11491_9489  0.0413994 
iB21_45_v n1_11583_9320 0  0.0413994 
iB21_45_g 0 n0_11491_9489  0.0413994 
iB21_46_v n1_11583_9503 0  0.0413994 
iB21_46_g 0 n0_11491_9489  0.0413994 
iB21_47_v n1_11583_9536 0  0.0413994 
iB21_47_g 0 n0_11491_9522  0.0413994 
iB21_48_v n1_11583_9719 0  0.0413994 
iB21_48_g 0 n0_11491_9705  0.0413994 
iB21_49_v n1_11583_9752 0  0.0413994 
iB21_49_g 0 n0_11491_9738  0.0413994 
iB21_50_v n1_11630_9503 0  0.0413994 
iB21_50_g 0 n0_11491_9489  0.0413994 
iB21_51_v n1_11630_9536 0  0.0413994 
iB21_51_g 0 n0_11491_9522  0.0413994 
iB21_52_v n1_11583_9935 0  0.0413994 
iB21_52_g 0 n0_11491_9921  0.0413994 
iB21_53_v n1_11583_9968 0  0.0413994 
iB21_53_g 0 n0_11491_9954  0.0413994 
iB21_54_v n1_11583_10151 0  0.0413994 
iB21_54_g 0 n0_11491_10137  0.0413994 
iB21_55_v n1_11583_10184 0  0.0413994 
iB21_55_g 0 n0_11491_10170  0.0413994 
iB21_56_v n1_11583_10367 0  0.0413994 
iB21_56_g 0 n0_11491_10353  0.0413994 
iB21_57_v n1_11583_10400 0  0.0413994 
iB21_57_g 0 n0_11491_10386  0.0413994 
iB21_58_v n1_11771_5350 0  0.0413994 
iB21_58_g 0 n0_12616_5385  0.0413994 
iB21_59_v n1_11771_5399 0  0.0413994 
iB21_59_g 0 n0_12616_5385  0.0413994 
iB21_60_v n1_11771_5432 0  0.0413994 
iB21_60_g 0 n0_12616_5418  0.0413994 
iB21_61_v n1_11771_5566 0  0.0413994 
iB21_61_g 0 n0_12616_5601  0.0413994 
iB21_62_v n1_11771_5615 0  0.0413994 
iB21_62_g 0 n0_12616_5601  0.0413994 
iB21_63_v n1_11771_5648 0  0.0413994 
iB21_63_g 0 n0_12616_5634  0.0413994 
iB21_64_v n1_11771_5782 0  0.0413994 
iB21_64_g 0 n0_12616_5817  0.0413994 
iB21_65_v n1_11771_5831 0  0.0413994 
iB21_65_g 0 n0_12616_5817  0.0413994 
iB21_66_v n1_11771_5864 0  0.0413994 
iB21_66_g 0 n0_12616_5850  0.0413994 
iB21_67_v n1_11771_6047 0  0.0413994 
iB21_67_g 0 n0_12616_6033  0.0413994 
iB21_68_v n1_11771_6080 0  0.0413994 
iB21_68_g 0 n0_12616_6066  0.0413994 
iB21_69_v n1_11771_6263 0  0.0413994 
iB21_69_g 0 n0_12616_6249  0.0413994 
iB21_70_v n1_11771_6296 0  0.0413994 
iB21_70_g 0 n0_12616_6282  0.0413994 
iB21_71_v n1_11771_6430 0  0.0413994 
iB21_71_g 0 n0_12616_6465  0.0413994 
iB21_72_v n1_11771_6479 0  0.0413994 
iB21_72_g 0 n0_12616_6465  0.0413994 
iB21_73_v n1_11771_6512 0  0.0413994 
iB21_73_g 0 n0_12616_6498  0.0413994 
iB21_74_v n1_11771_6646 0  0.0413994 
iB21_74_g 0 n0_12616_6681  0.0413994 
iB21_75_v n1_11771_6695 0  0.0413994 
iB21_75_g 0 n0_12616_6681  0.0413994 
iB21_76_v n1_11771_6728 0  0.0413994 
iB21_76_g 0 n0_12616_6714  0.0413994 
iB21_77_v n1_11771_6862 0  0.0413994 
iB21_77_g 0 n0_12616_6897  0.0413994 
iB21_78_v n1_11771_6911 0  0.0413994 
iB21_78_g 0 n0_12616_6897  0.0413994 
iB21_79_v n1_11771_6944 0  0.0413994 
iB21_79_g 0 n0_12616_6930  0.0413994 
iB21_80_v n1_11771_7078 0  0.0413994 
iB21_80_g 0 n0_12616_7113  0.0413994 
iB21_81_v n1_11771_7127 0  0.0413994 
iB21_81_g 0 n0_12616_7113  0.0413994 
iB21_82_v n1_11771_7160 0  0.0413994 
iB21_82_g 0 n0_12616_7146  0.0413994 
iB21_83_v n1_11771_7294 0  0.0413994 
iB21_83_g 0 n0_12616_7329  0.0413994 
iB21_84_v n1_11771_7343 0  0.0413994 
iB21_84_g 0 n0_12616_7329  0.0413994 
iB21_85_v n1_11771_7376 0  0.0413994 
iB21_85_g 0 n0_12616_7362  0.0413994 
iB21_86_v n1_11771_7510 0  0.0413994 
iB21_86_g 0 n0_12616_7545  0.0413994 
iB21_87_v n1_11771_7559 0  0.0413994 
iB21_87_g 0 n0_12616_7545  0.0413994 
iB21_88_v n1_11771_7592 0  0.0413994 
iB21_88_g 0 n0_12616_7578  0.0413994 
iB21_89_v n1_11771_7775 0  0.0413994 
iB21_89_g 0 n0_12616_7761  0.0413994 
iB21_90_v n1_11771_7808 0  0.0413994 
iB21_90_g 0 n0_12616_7794  0.0413994 
iB21_91_v n1_11771_7991 0  0.0413994 
iB21_91_g 0 n0_12616_7977  0.0413994 
iB21_92_v n1_11771_8024 0  0.0413994 
iB21_92_g 0 n0_12616_8010  0.0413994 
iB21_93_v n1_11771_8207 0  0.0413994 
iB21_93_g 0 n0_12616_8193  0.0413994 
iB21_94_v n1_11771_8240 0  0.0413994 
iB21_94_g 0 n0_12616_8226  0.0413994 
iB21_95_v n1_11771_8423 0  0.0413994 
iB21_95_g 0 n0_12616_8409  0.0413994 
iB21_96_v n1_11771_8456 0  0.0413994 
iB21_96_g 0 n0_12616_8442  0.0413994 
iB21_97_v n1_11771_8639 0  0.0413994 
iB21_97_g 0 n0_12616_8625  0.0413994 
iB21_98_v n1_11771_8672 0  0.0413994 
iB21_98_g 0 n0_12616_8658  0.0413994 
iB21_99_v n1_11771_8855 0  0.0413994 
iB21_99_g 0 n0_12616_8841  0.0413994 
iB21_100_v n1_11771_8888 0  0.0413994 
iB21_100_g 0 n0_12616_8874  0.0413994 
iB21_101_v n1_11771_9071 0  0.0413994 
iB21_101_g 0 n0_11491_9489  0.0413994 
iB21_102_v n1_11771_9104 0  0.0413994 
iB21_102_g 0 n0_11491_9489  0.0413994 
iB21_103_v n1_11771_9287 0  0.0413994 
iB21_103_g 0 n0_11491_9489  0.0413994 
iB21_104_v n1_11771_9320 0  0.0413994 
iB21_104_g 0 n0_11491_9489  0.0413994 
iB21_105_v n1_11771_9503 0  0.0413994 
iB21_105_g 0 n0_11491_9489  0.0413994 
iB21_106_v n1_11771_9536 0  0.0413994 
iB21_106_g 0 n0_11679_9705  0.0413994 
iB21_107_v n1_11771_9719 0  0.0413994 
iB21_107_g 0 n0_11679_9705  0.0413994 
iB21_108_v n1_11771_9752 0  0.0413994 
iB21_108_g 0 n0_11679_9738  0.0413994 
iB21_109_v n1_11771_9935 0  0.0413994 
iB21_109_g 0 n0_11679_9921  0.0413994 
iB21_110_v n1_11771_9968 0  0.0413994 
iB21_110_g 0 n0_11679_9954  0.0413994 
iB21_111_v n1_11771_10151 0  0.0413994 
iB21_111_g 0 n0_11679_10137  0.0413994 
iB21_112_v n1_11771_10184 0  0.0413994 
iB21_112_g 0 n0_11679_10170  0.0413994 
iB21_113_v n1_11771_10367 0  0.0413994 
iB21_113_g 0 n0_11679_10353  0.0413994 
iB21_114_v n1_11771_10400 0  0.0413994 
iB21_114_g 0 n0_11679_10386  0.0413994 
iB21_115_v n1_11771_10616 0  0.0413994 
iB21_115_g 0 n0_11679_10602  0.0413994 
iB21_116_v n1_13833_5350 0  0.0413994 
iB21_116_g 0 n0_12896_5385  0.0413994 
iB21_117_v n1_13833_5399 0  0.0413994 
iB21_117_g 0 n0_12896_5385  0.0413994 
iB21_118_v n1_13833_5432 0  0.0413994 
iB21_118_g 0 n0_12896_5418  0.0413994 
iB21_119_v n1_13833_5615 0  0.0413994 
iB21_119_g 0 n0_12896_5601  0.0413994 
iB21_120_v n1_13833_5648 0  0.0413994 
iB21_120_g 0 n0_12896_5634  0.0413994 
iB21_121_v n1_14021_5350 0  0.0413994 
iB21_121_g 0 n0_14866_5385  0.0413994 
iB21_122_v n1_14021_5399 0  0.0413994 
iB21_122_g 0 n0_14866_5385  0.0413994 
iB21_123_v n1_14021_5432 0  0.0413994 
iB21_123_g 0 n0_14866_5418  0.0413994 
iB21_124_v n1_14021_5615 0  0.0413994 
iB21_124_g 0 n0_14866_5601  0.0413994 
iB21_125_v n1_14021_5648 0  0.0413994 
iB21_125_g 0 n0_14866_5634  0.0413994 
iB21_126_v n1_13833_5782 0  0.0413994 
iB21_126_g 0 n0_12896_5817  0.0413994 
iB21_127_v n1_13833_5831 0  0.0413994 
iB21_127_g 0 n0_12896_5817  0.0413994 
iB21_128_v n1_13833_5864 0  0.0413994 
iB21_128_g 0 n0_12896_5850  0.0413994 
iB21_129_v n1_14021_5782 0  0.0413994 
iB21_129_g 0 n0_14866_5817  0.0413994 
iB21_130_v n1_14021_5831 0  0.0413994 
iB21_130_g 0 n0_14866_5817  0.0413994 
iB21_131_v n1_14021_5864 0  0.0413994 
iB21_131_g 0 n0_14866_5850  0.0413994 
iB21_132_v n1_14021_6047 0  0.0413994 
iB21_132_g 0 n0_14866_6033  0.0413994 
iB21_133_v n1_14021_6080 0  0.0413994 
iB21_133_g 0 n0_14866_6066  0.0413994 
iB21_134_v n1_13833_6263 0  0.0413994 
iB21_134_g 0 n0_12896_6249  0.0413994 
iB21_135_v n1_13833_6296 0  0.0413994 
iB21_135_g 0 n0_12896_6282  0.0413994 
iB21_136_v n1_13833_6430 0  0.0413994 
iB21_136_g 0 n0_12896_6465  0.0413994 
iB21_137_v n1_13833_6479 0  0.0413994 
iB21_137_g 0 n0_13741_7329  0.0413994 
iB21_138_v n1_13833_6512 0  0.0413994 
iB21_138_g 0 n0_13741_7329  0.0413994 
iB21_139_v n1_14021_6263 0  0.0413994 
iB21_139_g 0 n0_14866_6249  0.0413994 
iB21_140_v n1_14021_6296 0  0.0413994 
iB21_140_g 0 n0_14866_6282  0.0413994 
iB21_141_v n1_14021_6430 0  0.0413994 
iB21_141_g 0 n0_14866_6465  0.0413994 
iB21_142_v n1_14021_6479 0  0.0413994 
iB21_142_g 0 n0_13929_7329  0.0413994 
iB21_143_v n1_14021_6512 0  0.0413994 
iB21_143_g 0 n0_13929_7329  0.0413994 
iB21_144_v n1_13833_6646 0  0.0413994 
iB21_144_g 0 n0_13741_7329  0.0413994 
iB21_145_v n1_13833_6695 0  0.0413994 
iB21_145_g 0 n0_13741_7329  0.0413994 
iB21_146_v n1_13833_6728 0  0.0413994 
iB21_146_g 0 n0_13741_7329  0.0413994 
iB21_147_v n1_13833_6911 0  0.0413994 
iB21_147_g 0 n0_13741_7329  0.0413994 
iB21_148_v n1_14021_6646 0  0.0413994 
iB21_148_g 0 n0_13929_7329  0.0413994 
iB21_149_v n1_14021_6695 0  0.0413994 
iB21_149_g 0 n0_13929_7329  0.0413994 
iB21_150_v n1_14021_6728 0  0.0413994 
iB21_150_g 0 n0_13929_7329  0.0413994 
iB21_151_v n1_14021_6911 0  0.0413994 
iB21_151_g 0 n0_13929_7329  0.0413994 
iB21_152_v n1_13833_6944 0  0.0413994 
iB21_152_g 0 n0_13741_7329  0.0413994 
iB21_153_v n1_13833_7127 0  0.0413994 
iB21_153_g 0 n0_13741_7329  0.0413994 
iB21_154_v n1_13833_7160 0  0.0413994 
iB21_154_g 0 n0_13741_7329  0.0413994 
iB21_155_v n1_13880_7160 0  0.0413994 
iB21_155_g 0 n0_13929_7329  0.0413994 
iB21_156_v n1_14021_6944 0  0.0413994 
iB21_156_g 0 n0_13929_7329  0.0413994 
iB21_157_v n1_14021_7127 0  0.0413994 
iB21_157_g 0 n0_13929_7329  0.0413994 
iB21_158_v n1_14021_7160 0  0.0413994 
iB21_158_g 0 n0_13929_7329  0.0413994 
iB21_159_v n1_13833_7343 0  0.0413994 
iB21_159_g 0 n0_13741_7329  0.0413994 
iB21_160_v n1_13833_7376 0  0.0413994 
iB21_160_g 0 n0_13741_7362  0.0413994 
iB21_161_v n1_13833_7559 0  0.0413994 
iB21_161_g 0 n0_13741_7545  0.0413994 
iB21_162_v n1_13833_7592 0  0.0413994 
iB21_162_g 0 n0_13741_7578  0.0413994 
iB21_163_v n1_14021_7343 0  0.0413994 
iB21_163_g 0 n0_13929_7329  0.0413994 
iB21_164_v n1_14021_7376 0  0.0413994 
iB21_164_g 0 n0_13929_7362  0.0413994 
iB21_165_v n1_14021_7559 0  0.0413994 
iB21_165_g 0 n0_13929_7545  0.0413994 
iB21_166_v n1_14021_7592 0  0.0413994 
iB21_166_g 0 n0_13929_7578  0.0413994 
iB21_167_v n1_13833_7775 0  0.0413994 
iB21_167_g 0 n0_13741_7761  0.0413994 
iB21_168_v n1_13833_7808 0  0.0413994 
iB21_168_g 0 n0_13741_7794  0.0413994 
iB21_169_v n1_13833_7845 0  0.0413994 
iB21_169_g 0 n0_13741_7831  0.0413994 
iB21_170_v n1_13833_7942 0  0.0413994 
iB21_170_g 0 n0_13741_7977  0.0413994 
iB21_171_v n1_13833_7991 0  0.0413994 
iB21_171_g 0 n0_13741_7977  0.0413994 
iB21_172_v n1_13833_8024 0  0.0413994 
iB21_172_g 0 n0_13741_8010  0.0413994 
iB21_173_v n1_14021_7775 0  0.0413994 
iB21_173_g 0 n0_13929_7761  0.0413994 
iB21_174_v n1_14021_7808 0  0.0413994 
iB21_174_g 0 n0_13929_7794  0.0413994 
iB21_175_v n1_14021_7845 0  0.0413994 
iB21_175_g 0 n0_13929_7831  0.0413994 
iB21_176_v n1_14021_7942 0  0.0413994 
iB21_176_g 0 n0_13929_7977  0.0413994 
iB21_177_v n1_14021_7991 0  0.0413994 
iB21_177_g 0 n0_13929_7977  0.0413994 
iB21_178_v n1_14021_8024 0  0.0413994 
iB21_178_g 0 n0_13929_8010  0.0413994 
iB21_179_v n1_13833_8207 0  0.0413994 
iB21_179_g 0 n0_13741_8193  0.0413994 
iB21_180_v n1_13833_8240 0  0.0413994 
iB21_180_g 0 n0_13741_8226  0.0413994 
iB21_181_v n1_13833_8456 0  0.0413994 
iB21_181_g 0 n0_13880_8409  0.0413994 
iB21_182_v n1_14021_8207 0  0.0413994 
iB21_182_g 0 n0_13929_8193  0.0413994 
iB21_183_v n1_14021_8240 0  0.0413994 
iB21_183_g 0 n0_13929_8226  0.0413994 
iB21_184_v n1_14021_8423 0  0.0413994 
iB21_184_g 0 n0_13929_8409  0.0413994 
iB21_185_v n1_14021_8456 0  0.0413994 
iB21_185_g 0 n0_13929_8442  0.0413994 
iB21_186_v n1_13833_8639 0  0.0413994 
iB21_186_g 0 n0_13741_8625  0.0413994 
iB21_187_v n1_13833_8672 0  0.0413994 
iB21_187_g 0 n0_13741_8658  0.0413994 
iB21_188_v n1_13833_8806 0  0.0413994 
iB21_188_g 0 n0_13741_8841  0.0413994 
iB21_189_v n1_13833_8855 0  0.0413994 
iB21_189_g 0 n0_13741_8841  0.0413994 
iB21_190_v n1_13833_8888 0  0.0413994 
iB21_190_g 0 n0_13741_8874  0.0413994 
iB21_191_v n1_13833_8925 0  0.0413994 
iB21_191_g 0 n0_13741_8911  0.0413994 
iB21_192_v n1_14021_8639 0  0.0413994 
iB21_192_g 0 n0_13929_8625  0.0413994 
iB21_193_v n1_14021_8672 0  0.0413994 
iB21_193_g 0 n0_13929_8658  0.0413994 
iB21_194_v n1_14021_8806 0  0.0413994 
iB21_194_g 0 n0_13929_8841  0.0413994 
iB21_195_v n1_14021_8855 0  0.0413994 
iB21_195_g 0 n0_13929_8841  0.0413994 
iB21_196_v n1_14021_8888 0  0.0413994 
iB21_196_g 0 n0_13929_8874  0.0413994 
iB21_197_v n1_14021_8925 0  0.0413994 
iB21_197_g 0 n0_13929_8911  0.0413994 
iB21_198_v n1_13833_9022 0  0.0413994 
iB21_198_g 0 n0_13741_9057  0.0413994 
iB21_199_v n1_13833_9071 0  0.0413994 
iB21_199_g 0 n0_13741_9057  0.0413994 
iB21_200_v n1_13833_9104 0  0.0413994 
iB21_200_g 0 n0_13741_9090  0.0413994 
iB21_201_v n1_13833_9287 0  0.0413994 
iB21_201_g 0 n0_13741_9273  0.0413994 
iB21_202_v n1_13833_9320 0  0.0413994 
iB21_202_g 0 n0_13741_9306  0.0413994 
iB21_203_v n1_14021_9022 0  0.0413994 
iB21_203_g 0 n0_13929_9057  0.0413994 
iB21_204_v n1_14021_9071 0  0.0413994 
iB21_204_g 0 n0_13929_9057  0.0413994 
iB21_205_v n1_14021_9104 0  0.0413994 
iB21_205_g 0 n0_13929_9090  0.0413994 
iB21_206_v n1_14021_9287 0  0.0413994 
iB21_206_g 0 n0_13929_9273  0.0413994 
iB21_207_v n1_14021_9320 0  0.0413994 
iB21_207_g 0 n0_13929_9306  0.0413994 
iB21_208_v n1_13833_9503 0  0.0413994 
iB21_208_g 0 n0_13741_9489  0.0413994 
iB21_209_v n1_13833_9536 0  0.0413994 
iB21_209_g 0 n0_13741_9522  0.0413994 
iB21_210_v n1_13833_9719 0  0.0413994 
iB21_210_g 0 n0_13741_9705  0.0413994 
iB21_211_v n1_13833_9752 0  0.0413994 
iB21_211_g 0 n0_13741_9738  0.0413994 
iB21_212_v n1_13880_9503 0  0.0413994 
iB21_212_g 0 n0_13741_9489  0.0413994 
iB21_213_v n1_13880_9536 0  0.0413994 
iB21_213_g 0 n0_13741_9522  0.0413994 
iB21_214_v n1_14021_9503 0  0.0413994 
iB21_214_g 0 n0_13929_9306  0.0413994 
iB21_215_v n1_14021_9536 0  0.0413994 
iB21_215_g 0 n0_13929_9705  0.0413994 
iB21_216_v n1_14021_9719 0  0.0413994 
iB21_216_g 0 n0_13929_9705  0.0413994 
iB21_217_v n1_14021_9752 0  0.0413994 
iB21_217_g 0 n0_13929_9738  0.0413994 
iB21_218_v n1_13833_9886 0  0.0413994 
iB21_218_g 0 n0_13741_9921  0.0413994 
iB21_219_v n1_13833_9935 0  0.0413994 
iB21_219_g 0 n0_13741_9921  0.0413994 
iB21_220_v n1_13833_9968 0  0.0413994 
iB21_220_g 0 n0_13741_9954  0.0413994 
iB21_221_v n1_13833_10005 0  0.0413994 
iB21_221_g 0 n0_13741_9991  0.0413994 
iB21_222_v n1_13833_10102 0  0.0413994 
iB21_222_g 0 n0_13741_10137  0.0413994 
iB21_223_v n1_13833_10151 0  0.0413994 
iB21_223_g 0 n0_13741_10137  0.0413994 
iB21_224_v n1_13833_10184 0  0.0413994 
iB21_224_g 0 n0_13741_10170  0.0413994 
iB21_225_v n1_14021_9886 0  0.0413994 
iB21_225_g 0 n0_13929_9921  0.0413994 
iB21_226_v n1_14021_9935 0  0.0413994 
iB21_226_g 0 n0_13929_9921  0.0413994 
iB21_227_v n1_14021_9968 0  0.0413994 
iB21_227_g 0 n0_13929_9954  0.0413994 
iB21_228_v n1_14021_10005 0  0.0413994 
iB21_228_g 0 n0_13929_9991  0.0413994 
iB21_229_v n1_14021_10102 0  0.0413994 
iB21_229_g 0 n0_13929_10137  0.0413994 
iB21_230_v n1_14021_10151 0  0.0413994 
iB21_230_g 0 n0_13929_10137  0.0413994 
iB21_231_v n1_14021_10184 0  0.0413994 
iB21_231_g 0 n0_13929_10170  0.0413994 
iB21_232_v n1_13833_10367 0  0.0413994 
iB21_232_g 0 n0_13741_10353  0.0413994 
iB21_233_v n1_13833_10400 0  0.0413994 
iB21_233_g 0 n0_13741_10386  0.0413994 
iB21_234_v n1_14021_10367 0  0.0413994 
iB21_234_g 0 n0_13929_10353  0.0413994 
iB21_235_v n1_14021_10400 0  0.0413994 
iB21_235_g 0 n0_13929_10386  0.0413994 
iB21_236_v n1_14021_10616 0  0.0413994 
iB21_236_g 0 n0_13929_10602  0.0413994 
iB22_0_v n1_11583_10799 0  0.0480157 
iB22_0_g 0 n0_11491_10785  0.0480157 
iB22_1_v n1_11583_10832 0  0.0480157 
iB22_1_g 0 n0_11491_10818  0.0480157 
iB22_2_v n1_11583_11015 0  0.0480157 
iB22_2_g 0 n0_11491_11001  0.0480157 
iB22_3_v n1_11583_11048 0  0.0480157 
iB22_3_g 0 n0_11491_11034  0.0480157 
iB22_4_v n1_11583_11231 0  0.0480157 
iB22_4_g 0 n0_11491_11217  0.0480157 
iB22_5_v n1_11583_11264 0  0.0480157 
iB22_5_g 0 n0_11491_11250  0.0480157 
iB22_6_v n1_11583_11447 0  0.0480157 
iB22_6_g 0 n0_11491_11433  0.0480157 
iB22_7_v n1_11583_11480 0  0.0480157 
iB22_7_g 0 n0_11491_11466  0.0480157 
iB22_8_v n1_11583_11663 0  0.0480157 
iB22_8_g 0 n0_11491_11649  0.0480157 
iB22_9_v n1_11583_11696 0  0.0480157 
iB22_9_g 0 n0_11491_11682  0.0480157 
iB22_10_v n1_11630_11663 0  0.0480157 
iB22_10_g 0 n0_11491_11649  0.0480157 
iB22_11_v n1_11630_11696 0  0.0480157 
iB22_11_g 0 n0_11491_11682  0.0480157 
iB22_12_v n1_11583_11879 0  0.0480157 
iB22_12_g 0 n0_11491_11682  0.0480157 
iB22_13_v n1_11583_11912 0  0.0480157 
iB22_13_g 0 n0_11491_11682  0.0480157 
iB22_14_v n1_11583_12095 0  0.0480157 
iB22_14_g 0 n0_11491_11682  0.0480157 
iB22_15_v n1_11583_12128 0  0.0480157 
iB22_15_g 0 n0_11491_11682  0.0480157 
iB22_16_v n1_11583_12311 0  0.0480157 
iB22_16_g 0 n0_11491_11682  0.0480157 
iB22_17_v n1_11583_12344 0  0.0480157 
iB22_17_g 0 n0_11491_11682  0.0480157 
iB22_18_v n1_11583_12527 0  0.0480157 
iB22_18_g 0 n0_11491_11682  0.0480157 
iB22_19_v n1_11583_12560 0  0.0480157 
iB22_19_g 0 n0_10646_12566  0.0480157 
iB22_20_v n1_11583_12743 0  0.0480157 
iB22_20_g 0 n0_10646_12729  0.0480157 
iB22_21_v n1_11583_12959 0  0.0480157 
iB22_21_g 0 n0_10646_12945  0.0480157 
iB22_22_v n1_11583_12992 0  0.0480157 
iB22_22_g 0 n0_10646_12978  0.0480157 
iB22_23_v n1_11583_13175 0  0.0480157 
iB22_23_g 0 n0_10646_13161  0.0480157 
iB22_24_v n1_11583_13208 0  0.0480157 
iB22_24_g 0 n0_10646_13194  0.0480157 
iB22_25_v n1_11583_13391 0  0.0480157 
iB22_25_g 0 n0_10646_13377  0.0480157 
iB22_26_v n1_11583_13424 0  0.0480157 
iB22_26_g 0 n0_10646_13410  0.0480157 
iB22_27_v n1_11583_13607 0  0.0480157 
iB22_27_g 0 n0_10646_13593  0.0480157 
iB22_28_v n1_11583_13640 0  0.0480157 
iB22_28_g 0 n0_10646_13640  0.0480157 
iB22_29_v n1_11583_13774 0  0.0480157 
iB22_29_g 0 n0_10646_13809  0.0480157 
iB22_30_v n1_11583_13823 0  0.0480157 
iB22_30_g 0 n0_10646_13809  0.0480157 
iB22_31_v n1_11583_13856 0  0.0480157 
iB22_31_g 0 n0_10646_13856  0.0480157 
iB22_32_v n1_11583_14012 0  0.0480157 
iB22_32_g 0 n0_10646_14025  0.0480157 
iB22_33_v n1_11583_14039 0  0.0480157 
iB22_33_g 0 n0_10646_14025  0.0480157 
iB22_34_v n1_11583_14072 0  0.0480157 
iB22_34_g 0 n0_10646_14072  0.0480157 
iB22_35_v n1_11583_14220 0  0.0480157 
iB22_35_g 0 n0_10646_14241  0.0480157 
iB22_36_v n1_11583_14255 0  0.0480157 
iB22_36_g 0 n0_10646_14241  0.0480157 
iB22_37_v n1_11630_14012 0  0.0480157 
iB22_37_g 0 n0_10646_14025  0.0480157 
iB22_38_v n1_11630_14039 0  0.0480157 
iB22_38_g 0 n0_10646_14025  0.0480157 
iB22_39_v n1_11583_14288 0  0.0480157 
iB22_39_g 0 n0_10646_14274  0.0480157 
iB22_40_v n1_11583_14471 0  0.0480157 
iB22_40_g 0 n0_10646_14457  0.0480157 
iB22_41_v n1_11583_14504 0  0.0480157 
iB22_41_g 0 n0_10646_14504  0.0480157 
iB22_42_v n1_11583_14660 0  0.0480157 
iB22_42_g 0 n0_10646_14673  0.0480157 
iB22_43_v n1_11583_14687 0  0.0480157 
iB22_43_g 0 n0_10646_14673  0.0480157 
iB22_44_v n1_11583_14720 0  0.0480157 
iB22_44_g 0 n0_10646_14706  0.0480157 
iB22_45_v n1_11583_14903 0  0.0480157 
iB22_45_g 0 n0_10646_14889  0.0480157 
iB22_46_v n1_11583_14936 0  0.0480157 
iB22_46_g 0 n0_10646_14922  0.0480157 
iB22_47_v n1_11583_15335 0  0.0480157 
iB22_47_g 0 n0_10646_15321  0.0480157 
iB22_48_v n1_11583_15368 0  0.0480157 
iB22_48_g 0 n0_10646_15354  0.0480157 
iB22_49_v n1_11583_15551 0  0.0480157 
iB22_49_g 0 n0_10646_15537  0.0480157 
iB22_50_v n1_11583_15584 0  0.0480157 
iB22_50_g 0 n0_10646_15584  0.0480157 
iB22_51_v n1_11583_15740 0  0.0480157 
iB22_51_g 0 n0_10646_15753  0.0480157 
iB22_52_v n1_11583_15767 0  0.0480157 
iB22_52_g 0 n0_10646_15753  0.0480157 
iB22_53_v n1_11583_15800 0  0.0480157 
iB22_53_g 0 n0_10646_15800  0.0480157 
iB22_54_v n1_11771_10799 0  0.0480157 
iB22_54_g 0 n0_11679_10785  0.0480157 
iB22_55_v n1_11771_10832 0  0.0480157 
iB22_55_g 0 n0_11679_10818  0.0480157 
iB22_56_v n1_11771_11015 0  0.0480157 
iB22_56_g 0 n0_11679_11001  0.0480157 
iB22_57_v n1_11771_11048 0  0.0480157 
iB22_57_g 0 n0_11679_11034  0.0480157 
iB22_58_v n1_11771_11231 0  0.0480157 
iB22_58_g 0 n0_11679_11217  0.0480157 
iB22_59_v n1_11771_11264 0  0.0480157 
iB22_59_g 0 n0_11679_11250  0.0480157 
iB22_60_v n1_11771_11447 0  0.0480157 
iB22_60_g 0 n0_11679_11433  0.0480157 
iB22_61_v n1_11771_11480 0  0.0480157 
iB22_61_g 0 n0_11679_11466  0.0480157 
iB22_62_v n1_11771_11663 0  0.0480157 
iB22_62_g 0 n0_11679_11466  0.0480157 
iB22_63_v n1_11771_11696 0  0.0480157 
iB22_63_g 0 n0_11491_11682  0.0480157 
iB22_64_v n1_11771_11879 0  0.0480157 
iB22_64_g 0 n0_11491_11682  0.0480157 
iB22_65_v n1_11771_11912 0  0.0480157 
iB22_65_g 0 n0_11491_11682  0.0480157 
iB22_66_v n1_11771_12095 0  0.0480157 
iB22_66_g 0 n0_11491_11682  0.0480157 
iB22_67_v n1_11771_12128 0  0.0480157 
iB22_67_g 0 n0_11491_11682  0.0480157 
iB22_68_v n1_11771_12311 0  0.0480157 
iB22_68_g 0 n0_12616_12297  0.0480157 
iB22_69_v n1_11771_12344 0  0.0480157 
iB22_69_g 0 n0_12616_12330  0.0480157 
iB22_70_v n1_11771_12527 0  0.0480157 
iB22_70_g 0 n0_12616_12513  0.0480157 
iB22_71_v n1_11771_12560 0  0.0480157 
iB22_71_g 0 n0_12616_12546  0.0480157 
iB22_72_v n1_11771_12743 0  0.0480157 
iB22_72_g 0 n0_12616_12729  0.0480157 
iB22_73_v n1_11771_12776 0  0.0480157 
iB22_73_g 0 n0_12616_12762  0.0480157 
iB22_74_v n1_11771_12959 0  0.0480157 
iB22_74_g 0 n0_12616_12945  0.0480157 
iB22_75_v n1_11771_12992 0  0.0480157 
iB22_75_g 0 n0_12616_12978  0.0480157 
iB22_76_v n1_11771_13175 0  0.0480157 
iB22_76_g 0 n0_12616_13161  0.0480157 
iB22_77_v n1_11771_13208 0  0.0480157 
iB22_77_g 0 n0_12616_13194  0.0480157 
iB22_78_v n1_11771_13391 0  0.0480157 
iB22_78_g 0 n0_12616_13377  0.0480157 
iB22_79_v n1_11771_13424 0  0.0480157 
iB22_79_g 0 n0_12616_13410  0.0480157 
iB22_80_v n1_11771_13607 0  0.0480157 
iB22_80_g 0 n0_12616_13593  0.0480157 
iB22_81_v n1_11771_13640 0  0.0480157 
iB22_81_g 0 n0_12616_13626  0.0480157 
iB22_82_v n1_11771_13774 0  0.0480157 
iB22_82_g 0 n0_12616_13809  0.0480157 
iB22_83_v n1_11771_13823 0  0.0480157 
iB22_83_g 0 n0_12616_13809  0.0480157 
iB22_84_v n1_11771_13856 0  0.0480157 
iB22_84_g 0 n0_12616_13842  0.0480157 
iB22_85_v n1_11771_14012 0  0.0480157 
iB22_85_g 0 n0_12616_14025  0.0480157 
iB22_86_v n1_11771_14039 0  0.0480157 
iB22_86_g 0 n0_12616_14025  0.0480157 
iB22_87_v n1_11771_14072 0  0.0480157 
iB22_87_g 0 n0_12616_14079  0.0480157 
iB22_88_v n1_11771_14220 0  0.0480157 
iB22_88_g 0 n0_12616_14229  0.0480157 
iB22_89_v n1_11771_14255 0  0.0480157 
iB22_89_g 0 n0_12616_14241  0.0480157 
iB22_90_v n1_11771_14288 0  0.0480157 
iB22_90_g 0 n0_12616_14274  0.0480157 
iB22_91_v n1_11771_14471 0  0.0480157 
iB22_91_g 0 n0_12616_14457  0.0480157 
iB22_92_v n1_11771_14504 0  0.0480157 
iB22_92_g 0 n0_12616_14490  0.0480157 
iB22_93_v n1_11771_14660 0  0.0480157 
iB22_93_g 0 n0_12616_14673  0.0480157 
iB22_94_v n1_11771_14687 0  0.0480157 
iB22_94_g 0 n0_12616_14673  0.0480157 
iB22_95_v n1_11771_14720 0  0.0480157 
iB22_95_g 0 n0_12616_14727  0.0480157 
iB22_96_v n1_11771_14903 0  0.0480157 
iB22_96_g 0 n0_12616_14889  0.0480157 
iB22_97_v n1_11771_14936 0  0.0480157 
iB22_97_g 0 n0_12616_14922  0.0480157 
iB22_98_v n1_11771_15119 0  0.0480157 
iB22_98_g 0 n0_12616_15138  0.0480157 
iB22_99_v n1_11771_15152 0  0.0480157 
iB22_99_g 0 n0_12616_15138  0.0480157 
iB22_100_v n1_11771_15335 0  0.0480157 
iB22_100_g 0 n0_12616_15321  0.0480157 
iB22_101_v n1_11771_15368 0  0.0480157 
iB22_101_g 0 n0_12616_15368  0.0480157 
iB22_102_v n1_11771_15551 0  0.0480157 
iB22_102_g 0 n0_12616_15537  0.0480157 
iB22_103_v n1_11771_15584 0  0.0480157 
iB22_103_g 0 n0_12616_15570  0.0480157 
iB22_104_v n1_11771_15740 0  0.0480157 
iB22_104_g 0 n0_12616_15753  0.0480157 
iB22_105_v n1_11771_15767 0  0.0480157 
iB22_105_g 0 n0_12616_15753  0.0480157 
iB22_106_v n1_11771_15800 0  0.0480157 
iB22_106_g 0 n0_12616_15800  0.0480157 
iB22_107_v n1_13833_10799 0  0.0480157 
iB22_107_g 0 n0_13741_10785  0.0480157 
iB22_108_v n1_13833_10832 0  0.0480157 
iB22_108_g 0 n0_13741_10832  0.0480157 
iB22_109_v n1_13833_10988 0  0.0480157 
iB22_109_g 0 n0_13741_11001  0.0480157 
iB22_110_v n1_14021_10799 0  0.0480157 
iB22_110_g 0 n0_13929_10785  0.0480157 
iB22_111_v n1_14021_10832 0  0.0480157 
iB22_111_g 0 n0_13929_10832  0.0480157 
iB22_112_v n1_14021_10988 0  0.0480157 
iB22_112_g 0 n0_13929_11001  0.0480157 
iB22_113_v n1_13833_11015 0  0.0480157 
iB22_113_g 0 n0_13741_11001  0.0480157 
iB22_114_v n1_13833_11048 0  0.0480157 
iB22_114_g 0 n0_13741_11048  0.0480157 
iB22_115_v n1_13833_11204 0  0.0480157 
iB22_115_g 0 n0_13741_11217  0.0480157 
iB22_116_v n1_13833_11231 0  0.0480157 
iB22_116_g 0 n0_13741_11217  0.0480157 
iB22_117_v n1_13833_11264 0  0.0480157 
iB22_117_g 0 n0_13741_11250  0.0480157 
iB22_118_v n1_14021_11015 0  0.0480157 
iB22_118_g 0 n0_13929_11001  0.0480157 
iB22_119_v n1_14021_11048 0  0.0480157 
iB22_119_g 0 n0_13929_11048  0.0480157 
iB22_120_v n1_14021_11204 0  0.0480157 
iB22_120_g 0 n0_13929_11217  0.0480157 
iB22_121_v n1_14021_11231 0  0.0480157 
iB22_121_g 0 n0_13929_11217  0.0480157 
iB22_122_v n1_14021_11264 0  0.0480157 
iB22_122_g 0 n0_13929_11250  0.0480157 
iB22_123_v n1_13833_11447 0  0.0480157 
iB22_123_g 0 n0_13741_11433  0.0480157 
iB22_124_v n1_13833_11480 0  0.0480157 
iB22_124_g 0 n0_13741_11466  0.0480157 
iB22_125_v n1_13833_11663 0  0.0480157 
iB22_125_g 0 n0_13741_11649  0.0480157 
iB22_126_v n1_13833_11696 0  0.0480157 
iB22_126_g 0 n0_13741_11682  0.0480157 
iB22_127_v n1_13880_11663 0  0.0480157 
iB22_127_g 0 n0_13741_11649  0.0480157 
iB22_128_v n1_13880_11696 0  0.0480157 
iB22_128_g 0 n0_13741_11682  0.0480157 
iB22_129_v n1_14021_11447 0  0.0480157 
iB22_129_g 0 n0_13929_11433  0.0480157 
iB22_130_v n1_14021_11480 0  0.0480157 
iB22_130_g 0 n0_13929_11466  0.0480157 
iB22_131_v n1_14021_11663 0  0.0480157 
iB22_131_g 0 n0_13929_11466  0.0480157 
iB22_132_v n1_14021_11696 0  0.0480157 
iB22_132_g 0 n0_13929_11865  0.0480157 
iB22_133_v n1_13833_11879 0  0.0480157 
iB22_133_g 0 n0_13741_11865  0.0480157 
iB22_134_v n1_13833_11912 0  0.0480157 
iB22_134_g 0 n0_13741_11912  0.0480157 
iB22_135_v n1_13833_12068 0  0.0480157 
iB22_135_g 0 n0_13741_12081  0.0480157 
iB22_136_v n1_13833_12095 0  0.0480157 
iB22_136_g 0 n0_13741_12081  0.0480157 
iB22_137_v n1_13833_12128 0  0.0480157 
iB22_137_g 0 n0_13741_12128  0.0480157 
iB22_138_v n1_14021_11879 0  0.0480157 
iB22_138_g 0 n0_13929_11865  0.0480157 
iB22_139_v n1_14021_11912 0  0.0480157 
iB22_139_g 0 n0_13929_11912  0.0480157 
iB22_140_v n1_14021_12068 0  0.0480157 
iB22_140_g 0 n0_13929_12081  0.0480157 
iB22_141_v n1_14021_12095 0  0.0480157 
iB22_141_g 0 n0_13929_12081  0.0480157 
iB22_142_v n1_14021_12128 0  0.0480157 
iB22_142_g 0 n0_13929_12128  0.0480157 
iB22_143_v n1_13833_12284 0  0.0480157 
iB22_143_g 0 n0_13741_12297  0.0480157 
iB22_144_v n1_13833_12311 0  0.0480157 
iB22_144_g 0 n0_13741_12297  0.0480157 
iB22_145_v n1_13833_12344 0  0.0480157 
iB22_145_g 0 n0_13741_12330  0.0480157 
iB22_146_v n1_13833_12527 0  0.0480157 
iB22_146_g 0 n0_13741_12513  0.0480157 
iB22_147_v n1_13833_12560 0  0.0480157 
iB22_147_g 0 n0_13741_12546  0.0480157 
iB22_148_v n1_14021_12284 0  0.0480157 
iB22_148_g 0 n0_13929_12297  0.0480157 
iB22_149_v n1_14021_12311 0  0.0480157 
iB22_149_g 0 n0_13929_12297  0.0480157 
iB22_150_v n1_14021_12344 0  0.0480157 
iB22_150_g 0 n0_13929_12330  0.0480157 
iB22_151_v n1_14021_12527 0  0.0480157 
iB22_151_g 0 n0_13929_12513  0.0480157 
iB22_152_v n1_14021_12560 0  0.0480157 
iB22_152_g 0 n0_13929_12546  0.0480157 
iB22_153_v n1_13833_12743 0  0.0480157 
iB22_153_g 0 n0_13880_12776  0.0480157 
iB22_154_v n1_13833_12959 0  0.0480157 
iB22_154_g 0 n0_13741_12945  0.0480157 
iB22_155_v n1_13833_12992 0  0.0480157 
iB22_155_g 0 n0_13741_12992  0.0480157 
iB22_156_v n1_14021_12743 0  0.0480157 
iB22_156_g 0 n0_13929_12729  0.0480157 
iB22_157_v n1_14021_12776 0  0.0480157 
iB22_157_g 0 n0_13929_12776  0.0480157 
iB22_158_v n1_14021_12959 0  0.0480157 
iB22_158_g 0 n0_13929_12945  0.0480157 
iB22_159_v n1_14021_12992 0  0.0480157 
iB22_159_g 0 n0_13929_12992  0.0480157 
iB22_160_v n1_13833_13175 0  0.0480157 
iB22_160_g 0 n0_13741_13161  0.0480157 
iB22_161_v n1_13833_13208 0  0.0480157 
iB22_161_g 0 n0_13741_13194  0.0480157 
iB22_162_v n1_13833_13391 0  0.0480157 
iB22_162_g 0 n0_13741_13377  0.0480157 
iB22_163_v n1_13833_13424 0  0.0480157 
iB22_163_g 0 n0_13741_13423  0.0480157 
iB22_164_v n1_14021_13175 0  0.0480157 
iB22_164_g 0 n0_13929_13161  0.0480157 
iB22_165_v n1_14021_13208 0  0.0480157 
iB22_165_g 0 n0_13929_13194  0.0480157 
iB22_166_v n1_14021_13391 0  0.0480157 
iB22_166_g 0 n0_13929_13377  0.0480157 
iB22_167_v n1_14021_13424 0  0.0480157 
iB22_167_g 0 n0_13929_13423  0.0480157 
iB22_168_v n1_13833_13607 0  0.0480157 
iB22_168_g 0 n0_13741_13593  0.0480157 
iB22_169_v n1_13833_13640 0  0.0480157 
iB22_169_g 0 n0_13741_13626  0.0480157 
iB22_170_v n1_13833_13823 0  0.0480157 
iB22_170_g 0 n0_13741_13809  0.0480157 
iB22_171_v n1_13833_13856 0  0.0480157 
iB22_171_g 0 n0_13741_13842  0.0480157 
iB22_172_v n1_14021_13607 0  0.0480157 
iB22_172_g 0 n0_13929_13593  0.0480157 
iB22_173_v n1_14021_13640 0  0.0480157 
iB22_173_g 0 n0_13929_13626  0.0480157 
iB22_174_v n1_14021_13823 0  0.0480157 
iB22_174_g 0 n0_13929_13809  0.0480157 
iB22_175_v n1_14021_13856 0  0.0480157 
iB22_175_g 0 n0_13929_13842  0.0480157 
iB22_176_v n1_13833_14039 0  0.0480157 
iB22_176_g 0 n0_13741_13842  0.0480157 
iB22_177_v n1_13833_14072 0  0.0480157 
iB22_177_g 0 n0_13741_13842  0.0480157 
iB22_178_v n1_13833_14220 0  0.0480157 
iB22_178_g 0 n0_13741_13842  0.0480157 
iB22_179_v n1_13833_14255 0  0.0480157 
iB22_179_g 0 n0_13741_13842  0.0480157 
iB22_180_v n1_13880_14039 0  0.0480157 
iB22_180_g 0 n0_13929_13842  0.0480157 
iB22_181_v n1_14021_14039 0  0.0480157 
iB22_181_g 0 n0_13929_13842  0.0480157 
iB22_182_v n1_14021_14072 0  0.0480157 
iB22_182_g 0 n0_13929_13842  0.0480157 
iB22_183_v n1_14021_14220 0  0.0480157 
iB22_183_g 0 n0_13929_13842  0.0480157 
iB22_184_v n1_14021_14255 0  0.0480157 
iB22_184_g 0 n0_13929_13842  0.0480157 
iB22_185_v n1_13833_14288 0  0.0480157 
iB22_185_g 0 n0_13741_13842  0.0480157 
iB22_186_v n1_13833_14471 0  0.0480157 
iB22_186_g 0 n0_13741_13842  0.0480157 
iB22_187_v n1_13833_14504 0  0.0480157 
iB22_187_g 0 n0_13741_13842  0.0480157 
iB22_188_v n1_13833_14652 0  0.0480157 
iB22_188_g 0 n0_13741_13842  0.0480157 
iB22_189_v n1_14021_14288 0  0.0480157 
iB22_189_g 0 n0_13929_13842  0.0480157 
iB22_190_v n1_14021_14471 0  0.0480157 
iB22_190_g 0 n0_13929_13842  0.0480157 
iB22_191_v n1_14021_14504 0  0.0480157 
iB22_191_g 0 n0_13929_13842  0.0480157 
iB22_192_v n1_14021_14652 0  0.0480157 
iB22_192_g 0 n0_13929_13842  0.0480157 
iB22_193_v n1_13833_14687 0  0.0480157 
iB22_193_g 0 n0_13741_13842  0.0480157 
iB22_194_v n1_13833_14720 0  0.0480157 
iB22_194_g 0 n0_13741_13842  0.0480157 
iB22_195_v n1_13833_14868 0  0.0480157 
iB22_195_g 0 n0_12896_14889  0.0480157 
iB22_196_v n1_13833_14903 0  0.0480157 
iB22_196_g 0 n0_12896_14889  0.0480157 
iB22_197_v n1_13833_14936 0  0.0480157 
iB22_197_g 0 n0_12896_14922  0.0480157 
iB22_198_v n1_14021_14687 0  0.0480157 
iB22_198_g 0 n0_13929_13842  0.0480157 
iB22_199_v n1_14021_14720 0  0.0480157 
iB22_199_g 0 n0_13929_13842  0.0480157 
iB22_200_v n1_14021_14868 0  0.0480157 
iB22_200_g 0 n0_14866_14889  0.0480157 
iB22_201_v n1_14021_14903 0  0.0480157 
iB22_201_g 0 n0_14866_14889  0.0480157 
iB22_202_v n1_14021_14936 0  0.0480157 
iB22_202_g 0 n0_14866_14943  0.0480157 
iB22_203_v n1_13833_15335 0  0.0480157 
iB22_203_g 0 n0_12896_15321  0.0480157 
iB22_204_v n1_13833_15368 0  0.0480157 
iB22_204_g 0 n0_12896_15368  0.0480157 
iB22_205_v n1_14021_15119 0  0.0480157 
iB22_205_g 0 n0_14866_15138  0.0480157 
iB22_206_v n1_14021_15152 0  0.0480157 
iB22_206_g 0 n0_14866_15159  0.0480157 
iB22_207_v n1_14021_15335 0  0.0480157 
iB22_207_g 0 n0_14866_15321  0.0480157 
iB22_208_v n1_14021_15368 0  0.0480157 
iB22_208_g 0 n0_14866_15368  0.0480157 
iB22_209_v n1_13833_15524 0  0.0480157 
iB22_209_g 0 n0_12896_15537  0.0480157 
iB22_210_v n1_13833_15551 0  0.0480157 
iB22_210_g 0 n0_12896_15537  0.0480157 
iB22_211_v n1_13833_15584 0  0.0480157 
iB22_211_g 0 n0_12896_15570  0.0480157 
iB22_212_v n1_13833_15767 0  0.0480157 
iB22_212_g 0 n0_12896_15753  0.0480157 
iB22_213_v n1_13833_15800 0  0.0480157 
iB22_213_g 0 n0_12896_15800  0.0480157 
iB22_214_v n1_14021_15524 0  0.0480157 
iB22_214_g 0 n0_14866_15537  0.0480157 
iB22_215_v n1_14021_15551 0  0.0480157 
iB22_215_g 0 n0_14866_15537  0.0480157 
iB22_216_v n1_14021_15584 0  0.0480157 
iB22_216_g 0 n0_14866_15584  0.0480157 
iB22_217_v n1_14021_15767 0  0.0480157 
iB22_217_g 0 n0_14866_15753  0.0480157 
iB22_218_v n1_14021_15800 0  0.0480157 
iB22_218_g 0 n0_14866_15800  0.0480157 
iB23_0_v n1_11583_15948 0  0.0282587 
iB23_0_g 0 n0_10646_15969  0.0282587 
iB23_1_v n1_11583_15956 0  0.0282587 
iB23_1_g 0 n0_10646_15969  0.0282587 
iB23_2_v n1_11583_15983 0  0.0282587 
iB23_2_g 0 n0_10646_15969  0.0282587 
iB23_3_v n1_11583_16016 0  0.0282587 
iB23_3_g 0 n0_10646_16016  0.0282587 
iB23_4_v n1_11583_16172 0  0.0282587 
iB23_4_g 0 n0_10646_16185  0.0282587 
iB23_5_v n1_11583_16199 0  0.0282587 
iB23_5_g 0 n0_10646_16185  0.0282587 
iB23_6_v n1_11583_16232 0  0.0282587 
iB23_6_g 0 n0_10646_16185  0.0282587 
iB23_7_v n1_11630_16172 0  0.0282587 
iB23_7_g 0 n0_10646_16185  0.0282587 
iB23_8_v n1_11630_16199 0  0.0282587 
iB23_8_g 0 n0_10646_16185  0.0282587 
iB23_9_v n1_11630_16232 0  0.0282587 
iB23_9_g 0 n0_10646_16185  0.0282587 
iB23_10_v n1_11583_16415 0  0.0282587 
iB23_10_g 0 n0_10646_16401  0.0282587 
iB23_11_v n1_11583_16448 0  0.0282587 
iB23_11_g 0 n0_10646_16434  0.0282587 
iB23_12_v n1_11583_16604 0  0.0282587 
iB23_12_g 0 n0_10646_16617  0.0282587 
iB23_13_v n1_11583_16631 0  0.0282587 
iB23_13_g 0 n0_10646_16617  0.0282587 
iB23_14_v n1_11583_16664 0  0.0282587 
iB23_14_g 0 n0_10646_16650  0.0282587 
iB23_15_v n1_11583_16847 0  0.0282587 
iB23_15_g 0 n0_10646_16833  0.0282587 
iB23_16_v n1_11583_16880 0  0.0282587 
iB23_16_g 0 n0_10646_16866  0.0282587 
iB23_17_v n1_11583_17063 0  0.0282587 
iB23_17_g 0 n0_10646_17049  0.0282587 
iB23_18_v n1_11583_17096 0  0.0282587 
iB23_18_g 0 n0_10646_17096  0.0282587 
iB23_19_v n1_11583_17244 0  0.0282587 
iB23_19_g 0 n0_10646_17265  0.0282587 
iB23_20_v n1_11583_17468 0  0.0282587 
iB23_20_g 0 n0_10646_17481  0.0282587 
iB23_21_v n1_11583_17495 0  0.0282587 
iB23_21_g 0 n0_10646_17481  0.0282587 
iB23_22_v n1_11583_17528 0  0.0282587 
iB23_22_g 0 n0_10646_17514  0.0282587 
iB23_23_v n1_11583_17684 0  0.0282587 
iB23_23_g 0 n0_10646_17697  0.0282587 
iB23_24_v n1_11583_17711 0  0.0282587 
iB23_24_g 0 n0_10646_17697  0.0282587 
iB23_25_v n1_11583_17744 0  0.0282587 
iB23_25_g 0 n0_10646_17730  0.0282587 
iB23_26_v n1_11583_17927 0  0.0282587 
iB23_26_g 0 n0_10646_17913  0.0282587 
iB23_27_v n1_11583_17960 0  0.0282587 
iB23_27_g 0 n0_10646_17946  0.0282587 
iB23_28_v n1_11583_18143 0  0.0282587 
iB23_28_g 0 n0_10646_18129  0.0282587 
iB23_29_v n1_11583_18176 0  0.0282587 
iB23_29_g 0 n0_10646_18162  0.0282587 
iB23_30_v n1_11583_18332 0  0.0282587 
iB23_30_g 0 n0_10646_18345  0.0282587 
iB23_31_v n1_11400_18527 0  0.0282587 
iB23_31_g 0 n0_10646_18561  0.0282587 
iB23_32_v n1_11400_18548 0  0.0282587 
iB23_32_g 0 n0_10646_18561  0.0282587 
iB23_33_v n1_11400_18575 0  0.0282587 
iB23_33_g 0 n0_10646_18561  0.0282587 
iB23_34_v n1_11400_18608 0  0.0282587 
iB23_34_g 0 n0_10646_18608  0.0282587 
iB23_35_v n1_11583_18359 0  0.0282587 
iB23_35_g 0 n0_10646_18345  0.0282587 
iB23_36_v n1_11583_18392 0  0.0282587 
iB23_36_g 0 n0_10646_18392  0.0282587 
iB23_37_v n1_11583_18527 0  0.0282587 
iB23_37_g 0 n0_10646_18561  0.0282587 
iB23_38_v n1_11583_18548 0  0.0282587 
iB23_38_g 0 n0_10646_18561  0.0282587 
iB23_39_v n1_11583_18575 0  0.0282587 
iB23_39_g 0 n0_10646_18561  0.0282587 
iB23_40_v n1_11583_18608 0  0.0282587 
iB23_40_g 0 n0_10646_18608  0.0282587 
iB23_41_v n1_11630_18392 0  0.0282587 
iB23_41_g 0 n0_10646_18392  0.0282587 
iB23_42_v n1_11630_18527 0  0.0282587 
iB23_42_g 0 n0_10646_18561  0.0282587 
iB23_43_v n1_11630_18548 0  0.0282587 
iB23_43_g 0 n0_10646_18561  0.0282587 
iB23_44_v n1_11400_18764 0  0.0282587 
iB23_44_g 0 n0_10646_18777  0.0282587 
iB23_45_v n1_11400_18791 0  0.0282587 
iB23_45_g 0 n0_10646_18777  0.0282587 
iB23_46_v n1_11400_18824 0  0.0282587 
iB23_46_g 0 n0_10646_18810  0.0282587 
iB23_47_v n1_11400_19007 0  0.0282587 
iB23_47_g 0 n0_10646_18993  0.0282587 
iB23_48_v n1_11400_19040 0  0.0282587 
iB23_48_g 0 n0_10646_19026  0.0282587 
iB23_49_v n1_11583_18764 0  0.0282587 
iB23_49_g 0 n0_10646_18777  0.0282587 
iB23_50_v n1_11583_18791 0  0.0282587 
iB23_50_g 0 n0_10646_18777  0.0282587 
iB23_51_v n1_11583_18824 0  0.0282587 
iB23_51_g 0 n0_10646_18810  0.0282587 
iB23_52_v n1_11583_19007 0  0.0282587 
iB23_52_g 0 n0_10646_18993  0.0282587 
iB23_53_v n1_11583_19040 0  0.0282587 
iB23_53_g 0 n0_10646_19026  0.0282587 
iB23_54_v n1_11400_19223 0  0.0282587 
iB23_54_g 0 n0_10646_19209  0.0282587 
iB23_55_v n1_11400_19256 0  0.0282587 
iB23_55_g 0 n0_10646_19256  0.0282587 
iB23_56_v n1_11400_19412 0  0.0282587 
iB23_56_g 0 n0_10646_19425  0.0282587 
iB23_57_v n1_11400_19439 0  0.0282587 
iB23_57_g 0 n0_10646_19425  0.0282587 
iB23_58_v n1_11400_19472 0  0.0282587 
iB23_58_g 0 n0_10646_19458  0.0282587 
iB23_59_v n1_11583_19223 0  0.0282587 
iB23_59_g 0 n0_10646_19209  0.0282587 
iB23_60_v n1_11583_19256 0  0.0282587 
iB23_60_g 0 n0_10646_19256  0.0282587 
iB23_61_v n1_11583_19404 0  0.0282587 
iB23_61_g 0 n0_10646_19425  0.0282587 
iB23_62_v n1_11583_19412 0  0.0282587 
iB23_62_g 0 n0_10646_19425  0.0282587 
iB23_63_v n1_11583_19439 0  0.0282587 
iB23_63_g 0 n0_10646_19425  0.0282587 
iB23_64_v n1_11583_19472 0  0.0282587 
iB23_64_g 0 n0_10646_19458  0.0282587 
iB23_65_v n1_11400_19655 0  0.0282587 
iB23_65_g 0 n0_10646_19641  0.0282587 
iB23_66_v n1_11400_19688 0  0.0282587 
iB23_66_g 0 n0_10646_19674  0.0282587 
iB23_67_v n1_11400_19871 0  0.0282587 
iB23_67_g 0 n0_10646_19857  0.0282587 
iB23_68_v n1_11400_19904 0  0.0282587 
iB23_68_g 0 n0_10646_19890  0.0282587 
iB23_69_v n1_11583_19871 0  0.0282587 
iB23_69_g 0 n0_10646_19857  0.0282587 
iB23_70_v n1_11583_19904 0  0.0282587 
iB23_70_g 0 n0_10646_19890  0.0282587 
iB23_71_v n1_11400_20087 0  0.0282587 
iB23_71_g 0 n0_10646_20073  0.0282587 
iB23_72_v n1_11400_20120 0  0.0282587 
iB23_72_g 0 n0_10646_20106  0.0282587 
iB23_73_v n1_11400_20303 0  0.0282587 
iB23_73_g 0 n0_10646_20289  0.0282587 
iB23_74_v n1_11400_20336 0  0.0282587 
iB23_74_g 0 n0_10646_20322  0.0282587 
iB23_75_v n1_11583_20087 0  0.0282587 
iB23_75_g 0 n0_10646_20073  0.0282587 
iB23_76_v n1_11583_20120 0  0.0282587 
iB23_76_g 0 n0_10646_20106  0.0282587 
iB23_77_v n1_11583_20303 0  0.0282587 
iB23_77_g 0 n0_10646_20289  0.0282587 
iB23_78_v n1_11583_20336 0  0.0282587 
iB23_78_g 0 n0_10646_20322  0.0282587 
iB23_79_v n1_11400_20519 0  0.0282587 
iB23_79_g 0 n0_10646_20505  0.0282587 
iB23_80_v n1_11400_20552 0  0.0282587 
iB23_80_g 0 n0_10646_20538  0.0282587 
iB23_81_v n1_11400_20687 0  0.0282587 
iB23_81_g 0 n0_10646_20754  0.0282587 
iB23_82_v n1_11400_20735 0  0.0282587 
iB23_82_g 0 n0_10646_20754  0.0282587 
iB23_83_v n1_11400_20768 0  0.0282587 
iB23_83_g 0 n0_10646_20754  0.0282587 
iB23_84_v n1_11583_20519 0  0.0282587 
iB23_84_g 0 n0_10646_20505  0.0282587 
iB23_85_v n1_11583_20552 0  0.0282587 
iB23_85_g 0 n0_10646_20538  0.0282587 
iB23_86_v n1_11583_20687 0  0.0282587 
iB23_86_g 0 n0_10646_20754  0.0282587 
iB23_87_v n1_11583_20735 0  0.0282587 
iB23_87_g 0 n0_10646_20754  0.0282587 
iB23_88_v n1_11583_20768 0  0.0282587 
iB23_88_g 0 n0_10646_20754  0.0282587 
iB23_89_v n1_11630_20687 0  0.0282587 
iB23_89_g 0 n0_10646_20754  0.0282587 
iB23_90_v n1_11630_20735 0  0.0282587 
iB23_90_g 0 n0_10646_20754  0.0282587 
iB23_91_v n1_11630_20768 0  0.0282587 
iB23_91_g 0 n0_10646_20754  0.0282587 
iB23_92_v n1_11400_20951 0  0.0282587 
iB23_92_g 0 n0_10646_20937  0.0282587 
iB23_93_v n1_11400_20984 0  0.0282587 
iB23_93_g 0 n0_10646_20970  0.0282587 
iB23_94_v n1_11583_20951 0  0.0282587 
iB23_94_g 0 n0_10646_20937  0.0282587 
iB23_95_v n1_11583_20984 0  0.0282587 
iB23_95_g 0 n0_10646_20970  0.0282587 
iB23_96_v n1_11771_15948 0  0.0282587 
iB23_96_g 0 n0_12616_15969  0.0282587 
iB23_97_v n1_11771_15956 0  0.0282587 
iB23_97_g 0 n0_12616_15969  0.0282587 
iB23_98_v n1_11771_15983 0  0.0282587 
iB23_98_g 0 n0_12616_15969  0.0282587 
iB23_99_v n1_11771_16016 0  0.0282587 
iB23_99_g 0 n0_12616_16002  0.0282587 
iB23_100_v n1_11771_16172 0  0.0282587 
iB23_100_g 0 n0_12616_16185  0.0282587 
iB23_101_v n1_11771_16199 0  0.0282587 
iB23_101_g 0 n0_12616_16185  0.0282587 
iB23_102_v n1_11771_16415 0  0.0282587 
iB23_102_g 0 n0_12616_16401  0.0282587 
iB23_103_v n1_11771_16448 0  0.0282587 
iB23_103_g 0 n0_12616_16448  0.0282587 
iB23_104_v n1_11771_16604 0  0.0282587 
iB23_104_g 0 n0_12616_16617  0.0282587 
iB23_105_v n1_11771_16631 0  0.0282587 
iB23_105_g 0 n0_12616_16617  0.0282587 
iB23_106_v n1_11771_16664 0  0.0282587 
iB23_106_g 0 n0_12616_16650  0.0282587 
iB23_107_v n1_11771_16847 0  0.0282587 
iB23_107_g 0 n0_12616_16833  0.0282587 
iB23_108_v n1_11771_16880 0  0.0282587 
iB23_108_g 0 n0_12616_16866  0.0282587 
iB23_109_v n1_11771_17063 0  0.0282587 
iB23_109_g 0 n0_12616_17049  0.0282587 
iB23_110_v n1_11771_17096 0  0.0282587 
iB23_110_g 0 n0_12616_17096  0.0282587 
iB23_111_v n1_11771_17244 0  0.0282587 
iB23_111_g 0 n0_12616_17265  0.0282587 
iB23_112_v n1_11771_17279 0  0.0282587 
iB23_112_g 0 n0_12616_17265  0.0282587 
iB23_113_v n1_11771_17312 0  0.0282587 
iB23_113_g 0 n0_12616_17298  0.0282587 
iB23_114_v n1_11771_17468 0  0.0282587 
iB23_114_g 0 n0_12616_17481  0.0282587 
iB23_115_v n1_11771_17495 0  0.0282587 
iB23_115_g 0 n0_12616_17481  0.0282587 
iB23_116_v n1_11771_17528 0  0.0282587 
iB23_116_g 0 n0_12616_17528  0.0282587 
iB23_117_v n1_11771_17684 0  0.0282587 
iB23_117_g 0 n0_12616_17697  0.0282587 
iB23_118_v n1_11771_17711 0  0.0282587 
iB23_118_g 0 n0_12616_17697  0.0282587 
iB23_119_v n1_11771_17744 0  0.0282587 
iB23_119_g 0 n0_12616_17730  0.0282587 
iB23_120_v n1_11771_17927 0  0.0282587 
iB23_120_g 0 n0_12616_17913  0.0282587 
iB23_121_v n1_11771_17960 0  0.0282587 
iB23_121_g 0 n0_12616_17946  0.0282587 
iB23_122_v n1_11771_18143 0  0.0282587 
iB23_122_g 0 n0_12616_18129  0.0282587 
iB23_123_v n1_11771_18176 0  0.0282587 
iB23_123_g 0 n0_12616_18176  0.0282587 
iB23_124_v n1_11771_18332 0  0.0282587 
iB23_124_g 0 n0_12616_18345  0.0282587 
iB23_125_v n1_11771_18359 0  0.0282587 
iB23_125_g 0 n0_12616_18345  0.0282587 
iB23_126_v n1_11771_18392 0  0.0282587 
iB23_126_g 0 n0_12616_18378  0.0282587 
iB23_127_v n1_11771_18527 0  0.0282587 
iB23_127_g 0 n0_12616_18561  0.0282587 
iB23_128_v n1_11771_18548 0  0.0282587 
iB23_128_g 0 n0_12616_18561  0.0282587 
iB23_129_v n1_11771_18575 0  0.0282587 
iB23_129_g 0 n0_12616_18561  0.0282587 
iB23_130_v n1_11771_18608 0  0.0282587 
iB23_130_g 0 n0_12616_18608  0.0282587 
iB23_131_v n1_11864_18527 0  0.0282587 
iB23_131_g 0 n0_12616_18561  0.0282587 
iB23_132_v n1_11864_18575 0  0.0282587 
iB23_132_g 0 n0_12616_18561  0.0282587 
iB23_133_v n1_11864_18608 0  0.0282587 
iB23_133_g 0 n0_12616_18608  0.0282587 
iB23_134_v n1_11771_18764 0  0.0282587 
iB23_134_g 0 n0_12616_18777  0.0282587 
iB23_135_v n1_11771_18791 0  0.0282587 
iB23_135_g 0 n0_12616_18777  0.0282587 
iB23_136_v n1_11771_18824 0  0.0282587 
iB23_136_g 0 n0_12616_18810  0.0282587 
iB23_137_v n1_11771_19007 0  0.0282587 
iB23_137_g 0 n0_12616_18993  0.0282587 
iB23_138_v n1_11771_19040 0  0.0282587 
iB23_138_g 0 n0_12616_19026  0.0282587 
iB23_139_v n1_11864_18764 0  0.0282587 
iB23_139_g 0 n0_12616_18777  0.0282587 
iB23_140_v n1_11864_18791 0  0.0282587 
iB23_140_g 0 n0_12616_18777  0.0282587 
iB23_141_v n1_11864_18824 0  0.0282587 
iB23_141_g 0 n0_12616_18810  0.0282587 
iB23_142_v n1_11864_19007 0  0.0282587 
iB23_142_g 0 n0_12616_18993  0.0282587 
iB23_143_v n1_11864_19040 0  0.0282587 
iB23_143_g 0 n0_12616_19026  0.0282587 
iB23_144_v n1_11771_19223 0  0.0282587 
iB23_144_g 0 n0_12616_19209  0.0282587 
iB23_145_v n1_11771_19256 0  0.0282587 
iB23_145_g 0 n0_12616_19256  0.0282587 
iB23_146_v n1_11771_19404 0  0.0282587 
iB23_146_g 0 n0_12616_19425  0.0282587 
iB23_147_v n1_11771_19412 0  0.0282587 
iB23_147_g 0 n0_12616_19425  0.0282587 
iB23_148_v n1_11771_19439 0  0.0282587 
iB23_148_g 0 n0_12616_19425  0.0282587 
iB23_149_v n1_11771_19472 0  0.0282587 
iB23_149_g 0 n0_12616_19458  0.0282587 
iB23_150_v n1_11864_19223 0  0.0282587 
iB23_150_g 0 n0_12616_19209  0.0282587 
iB23_151_v n1_11864_19256 0  0.0282587 
iB23_151_g 0 n0_12616_19256  0.0282587 
iB23_152_v n1_11864_19404 0  0.0282587 
iB23_152_g 0 n0_12616_19425  0.0282587 
iB23_153_v n1_11864_19439 0  0.0282587 
iB23_153_g 0 n0_12616_19425  0.0282587 
iB23_154_v n1_11864_19472 0  0.0282587 
iB23_154_g 0 n0_12616_19458  0.0282587 
iB23_155_v n1_11771_19655 0  0.0282587 
iB23_155_g 0 n0_12616_19641  0.0282587 
iB23_156_v n1_11771_19688 0  0.0282587 
iB23_156_g 0 n0_12616_19674  0.0282587 
iB23_157_v n1_11771_19871 0  0.0282587 
iB23_157_g 0 n0_12616_19857  0.0282587 
iB23_158_v n1_11771_19904 0  0.0282587 
iB23_158_g 0 n0_12616_19890  0.0282587 
iB23_159_v n1_11864_19655 0  0.0282587 
iB23_159_g 0 n0_12616_19641  0.0282587 
iB23_160_v n1_11864_19688 0  0.0282587 
iB23_160_g 0 n0_12616_19674  0.0282587 
iB23_161_v n1_11864_19871 0  0.0282587 
iB23_161_g 0 n0_12616_19857  0.0282587 
iB23_162_v n1_11864_19904 0  0.0282587 
iB23_162_g 0 n0_12616_19890  0.0282587 
iB23_163_v n1_11771_20087 0  0.0282587 
iB23_163_g 0 n0_12616_20073  0.0282587 
iB23_164_v n1_11771_20120 0  0.0282587 
iB23_164_g 0 n0_12616_20106  0.0282587 
iB23_165_v n1_11771_20303 0  0.0282587 
iB23_165_g 0 n0_12616_20289  0.0282587 
iB23_166_v n1_11771_20336 0  0.0282587 
iB23_166_g 0 n0_12616_20322  0.0282587 
iB23_167_v n1_11864_20087 0  0.0282587 
iB23_167_g 0 n0_12616_20073  0.0282587 
iB23_168_v n1_11864_20120 0  0.0282587 
iB23_168_g 0 n0_12616_20106  0.0282587 
iB23_169_v n1_11864_20303 0  0.0282587 
iB23_169_g 0 n0_12616_20289  0.0282587 
iB23_170_v n1_11864_20336 0  0.0282587 
iB23_170_g 0 n0_12616_20322  0.0282587 
iB23_171_v n1_11771_20519 0  0.0282587 
iB23_171_g 0 n0_12616_20505  0.0282587 
iB23_172_v n1_11771_20552 0  0.0282587 
iB23_172_g 0 n0_12616_20538  0.0282587 
iB23_173_v n1_11771_20687 0  0.0282587 
iB23_173_g 0 n0_12616_20754  0.0282587 
iB23_174_v n1_11771_20768 0  0.0282587 
iB23_174_g 0 n0_12616_20754  0.0282587 
iB23_175_v n1_11864_20519 0  0.0282587 
iB23_175_g 0 n0_12616_20505  0.0282587 
iB23_176_v n1_11864_20552 0  0.0282587 
iB23_176_g 0 n0_12616_20538  0.0282587 
iB23_177_v n1_11864_20687 0  0.0282587 
iB23_177_g 0 n0_12616_20754  0.0282587 
iB23_178_v n1_11864_20735 0  0.0282587 
iB23_178_g 0 n0_12616_20754  0.0282587 
iB23_179_v n1_11864_20768 0  0.0282587 
iB23_179_g 0 n0_12616_20754  0.0282587 
iB23_180_v n1_11771_20951 0  0.0282587 
iB23_180_g 0 n0_12616_20937  0.0282587 
iB23_181_v n1_11771_20984 0  0.0282587 
iB23_181_g 0 n0_12616_20970  0.0282587 
iB23_182_v n1_11864_20951 0  0.0282587 
iB23_182_g 0 n0_12616_20937  0.0282587 
iB23_183_v n1_11864_20984 0  0.0282587 
iB23_183_g 0 n0_12616_20970  0.0282587 
iB23_184_v n1_13650_18527 0  0.0282587 
iB23_184_g 0 n0_12896_18561  0.0282587 
iB23_185_v n1_13650_18575 0  0.0282587 
iB23_185_g 0 n0_12896_18561  0.0282587 
iB23_186_v n1_13650_18608 0  0.0282587 
iB23_186_g 0 n0_12896_18608  0.0282587 
iB23_187_v n1_13650_18764 0  0.0282587 
iB23_187_g 0 n0_12896_18777  0.0282587 
iB23_188_v n1_13650_18791 0  0.0282587 
iB23_188_g 0 n0_12896_18777  0.0282587 
iB23_189_v n1_13650_18824 0  0.0282587 
iB23_189_g 0 n0_12896_18810  0.0282587 
iB23_190_v n1_13650_19007 0  0.0282587 
iB23_190_g 0 n0_12896_18993  0.0282587 
iB23_191_v n1_13650_19040 0  0.0282587 
iB23_191_g 0 n0_12896_19026  0.0282587 
iB23_192_v n1_13650_19223 0  0.0282587 
iB23_192_g 0 n0_12896_19209  0.0282587 
iB23_193_v n1_13650_19256 0  0.0282587 
iB23_193_g 0 n0_12896_19256  0.0282587 
iB23_194_v n1_13650_19412 0  0.0282587 
iB23_194_g 0 n0_12896_19425  0.0282587 
iB23_195_v n1_13650_19439 0  0.0282587 
iB23_195_g 0 n0_12896_19425  0.0282587 
iB23_196_v n1_13650_19472 0  0.0282587 
iB23_196_g 0 n0_12896_19458  0.0282587 
iB23_197_v n1_13650_19655 0  0.0282587 
iB23_197_g 0 n0_12896_19641  0.0282587 
iB23_198_v n1_13650_19688 0  0.0282587 
iB23_198_g 0 n0_12896_19674  0.0282587 
iB23_199_v n1_13650_19871 0  0.0282587 
iB23_199_g 0 n0_12896_19857  0.0282587 
iB23_200_v n1_13650_19904 0  0.0282587 
iB23_200_g 0 n0_12896_19890  0.0282587 
iB23_201_v n1_13650_20087 0  0.0282587 
iB23_201_g 0 n0_12896_20073  0.0282587 
iB23_202_v n1_13650_20120 0  0.0282587 
iB23_202_g 0 n0_12896_20106  0.0282587 
iB23_203_v n1_13650_20303 0  0.0282587 
iB23_203_g 0 n0_12896_20289  0.0282587 
iB23_204_v n1_13650_20336 0  0.0282587 
iB23_204_g 0 n0_12896_20322  0.0282587 
iB23_205_v n1_13650_20519 0  0.0282587 
iB23_205_g 0 n0_12896_20505  0.0282587 
iB23_206_v n1_13650_20552 0  0.0282587 
iB23_206_g 0 n0_12896_20538  0.0282587 
iB23_207_v n1_13650_20687 0  0.0282587 
iB23_207_g 0 n0_12896_20754  0.0282587 
iB23_208_v n1_13650_20735 0  0.0282587 
iB23_208_g 0 n0_12896_20754  0.0282587 
iB23_209_v n1_13650_20768 0  0.0282587 
iB23_209_g 0 n0_12896_20754  0.0282587 
iB23_210_v n1_13650_20951 0  0.0282587 
iB23_210_g 0 n0_12896_20937  0.0282587 
iB23_211_v n1_13650_20984 0  0.0282587 
iB23_211_g 0 n0_12896_20970  0.0282587 
iB23_212_v n1_13833_15956 0  0.0282587 
iB23_212_g 0 n0_12896_15969  0.0282587 
iB23_213_v n1_13833_15983 0  0.0282587 
iB23_213_g 0 n0_12896_15969  0.0282587 
iB23_214_v n1_13833_16016 0  0.0282587 
iB23_214_g 0 n0_12896_16002  0.0282587 
iB23_215_v n1_13833_16199 0  0.0282587 
iB23_215_g 0 n0_12896_16185  0.0282587 
iB23_216_v n1_13833_16232 0  0.0282587 
iB23_216_g 0 n0_12896_16185  0.0282587 
iB23_217_v n1_13880_16199 0  0.0282587 
iB23_217_g 0 n0_12896_16185  0.0282587 
iB23_218_v n1_13880_16232 0  0.0282587 
iB23_218_g 0 n0_12896_16185  0.0282587 
iB23_219_v n1_14021_15956 0  0.0282587 
iB23_219_g 0 n0_14866_15969  0.0282587 
iB23_220_v n1_14021_15983 0  0.0282587 
iB23_220_g 0 n0_14866_15969  0.0282587 
iB23_221_v n1_14021_16016 0  0.0282587 
iB23_221_g 0 n0_14866_16002  0.0282587 
iB23_222_v n1_14021_16199 0  0.0282587 
iB23_222_g 0 n0_14866_16185  0.0282587 
iB23_223_v n1_13833_16415 0  0.0282587 
iB23_223_g 0 n0_12896_16401  0.0282587 
iB23_224_v n1_13833_16448 0  0.0282587 
iB23_224_g 0 n0_12896_16448  0.0282587 
iB23_225_v n1_13833_16604 0  0.0282587 
iB23_225_g 0 n0_12896_16617  0.0282587 
iB23_226_v n1_13833_16631 0  0.0282587 
iB23_226_g 0 n0_12896_16617  0.0282587 
iB23_227_v n1_13833_16664 0  0.0282587 
iB23_227_g 0 n0_12896_16650  0.0282587 
iB23_228_v n1_14021_16415 0  0.0282587 
iB23_228_g 0 n0_14866_16401  0.0282587 
iB23_229_v n1_14021_16448 0  0.0282587 
iB23_229_g 0 n0_14866_16448  0.0282587 
iB23_230_v n1_14021_16604 0  0.0282587 
iB23_230_g 0 n0_14866_16617  0.0282587 
iB23_231_v n1_14021_16631 0  0.0282587 
iB23_231_g 0 n0_14866_16617  0.0282587 
iB23_232_v n1_14021_16664 0  0.0282587 
iB23_232_g 0 n0_14866_16650  0.0282587 
iB23_233_v n1_13833_16847 0  0.0282587 
iB23_233_g 0 n0_12896_16833  0.0282587 
iB23_234_v n1_13833_16880 0  0.0282587 
iB23_234_g 0 n0_12896_16866  0.0282587 
iB23_235_v n1_13833_17063 0  0.0282587 
iB23_235_g 0 n0_12896_17049  0.0282587 
iB23_236_v n1_13833_17096 0  0.0282587 
iB23_236_g 0 n0_12896_17096  0.0282587 
iB23_237_v n1_14021_16847 0  0.0282587 
iB23_237_g 0 n0_14866_16833  0.0282587 
iB23_238_v n1_14021_16880 0  0.0282587 
iB23_238_g 0 n0_14866_16866  0.0282587 
iB23_239_v n1_14021_17063 0  0.0282587 
iB23_239_g 0 n0_14866_17049  0.0282587 
iB23_240_v n1_14021_17096 0  0.0282587 
iB23_240_g 0 n0_14866_17096  0.0282587 
iB23_241_v n1_13833_17495 0  0.0282587 
iB23_241_g 0 n0_12896_17481  0.0282587 
iB23_242_v n1_14021_17252 0  0.0282587 
iB23_242_g 0 n0_14866_17265  0.0282587 
iB23_243_v n1_14021_17279 0  0.0282587 
iB23_243_g 0 n0_14866_17265  0.0282587 
iB23_244_v n1_14021_17312 0  0.0282587 
iB23_244_g 0 n0_14866_17298  0.0282587 
iB23_245_v n1_14021_17495 0  0.0282587 
iB23_245_g 0 n0_14866_17481  0.0282587 
iB23_246_v n1_13833_17528 0  0.0282587 
iB23_246_g 0 n0_12896_17528  0.0282587 
iB23_247_v n1_13833_17684 0  0.0282587 
iB23_247_g 0 n0_12896_17697  0.0282587 
iB23_248_v n1_13833_17711 0  0.0282587 
iB23_248_g 0 n0_12896_17697  0.0282587 
iB23_249_v n1_13833_17744 0  0.0282587 
iB23_249_g 0 n0_12896_17730  0.0282587 
iB23_250_v n1_13833_17927 0  0.0282587 
iB23_250_g 0 n0_12896_17913  0.0282587 
iB23_251_v n1_14021_17528 0  0.0282587 
iB23_251_g 0 n0_14866_17528  0.0282587 
iB23_252_v n1_14021_17684 0  0.0282587 
iB23_252_g 0 n0_14866_17697  0.0282587 
iB23_253_v n1_14021_17711 0  0.0282587 
iB23_253_g 0 n0_14866_17697  0.0282587 
iB23_254_v n1_14021_17744 0  0.0282587 
iB23_254_g 0 n0_14866_17730  0.0282587 
iB23_255_v n1_14021_17927 0  0.0282587 
iB23_255_g 0 n0_14866_17913  0.0282587 
iB23_256_v n1_13833_17960 0  0.0282587 
iB23_256_g 0 n0_12896_17946  0.0282587 
iB23_257_v n1_13833_18094 0  0.0282587 
iB23_257_g 0 n0_12896_18129  0.0282587 
iB23_258_v n1_13833_18143 0  0.0282587 
iB23_258_g 0 n0_12896_18129  0.0282587 
iB23_259_v n1_13833_18176 0  0.0282587 
iB23_259_g 0 n0_12896_18176  0.0282587 
iB23_260_v n1_13833_18324 0  0.0282587 
iB23_260_g 0 n0_12896_18345  0.0282587 
iB23_261_v n1_13833_18332 0  0.0282587 
iB23_261_g 0 n0_12896_18345  0.0282587 
iB23_262_v n1_14021_17960 0  0.0282587 
iB23_262_g 0 n0_14866_17946  0.0282587 
iB23_263_v n1_14021_18094 0  0.0282587 
iB23_263_g 0 n0_14866_18129  0.0282587 
iB23_264_v n1_14021_18143 0  0.0282587 
iB23_264_g 0 n0_14866_18129  0.0282587 
iB23_265_v n1_14021_18176 0  0.0282587 
iB23_265_g 0 n0_14866_18176  0.0282587 
iB23_266_v n1_14021_18324 0  0.0282587 
iB23_266_g 0 n0_14866_18345  0.0282587 
iB23_267_v n1_14021_18332 0  0.0282587 
iB23_267_g 0 n0_14866_18345  0.0282587 
iB23_268_v n1_13833_18359 0  0.0282587 
iB23_268_g 0 n0_12896_18345  0.0282587 
iB23_269_v n1_13833_18392 0  0.0282587 
iB23_269_g 0 n0_12896_18378  0.0282587 
iB23_270_v n1_13833_18527 0  0.0282587 
iB23_270_g 0 n0_12896_18561  0.0282587 
iB23_271_v n1_13833_18575 0  0.0282587 
iB23_271_g 0 n0_12896_18561  0.0282587 
iB23_272_v n1_13833_18608 0  0.0282587 
iB23_272_g 0 n0_12896_18608  0.0282587 
iB23_273_v n1_13880_18392 0  0.0282587 
iB23_273_g 0 n0_12896_18378  0.0282587 
iB23_274_v n1_13880_18527 0  0.0282587 
iB23_274_g 0 n0_12896_18561  0.0282587 
iB23_275_v n1_14021_18359 0  0.0282587 
iB23_275_g 0 n0_14866_18345  0.0282587 
iB23_276_v n1_14021_18392 0  0.0282587 
iB23_276_g 0 n0_14866_18378  0.0282587 
iB23_277_v n1_14021_18527 0  0.0282587 
iB23_277_g 0 n0_14866_18561  0.0282587 
iB23_278_v n1_14021_18575 0  0.0282587 
iB23_278_g 0 n0_14866_18561  0.0282587 
iB23_279_v n1_14021_18608 0  0.0282587 
iB23_279_g 0 n0_14866_18608  0.0282587 
iB23_280_v n1_14114_18527 0  0.0282587 
iB23_280_g 0 n0_14866_18561  0.0282587 
iB23_281_v n1_14114_18575 0  0.0282587 
iB23_281_g 0 n0_14866_18561  0.0282587 
iB23_282_v n1_14114_18608 0  0.0282587 
iB23_282_g 0 n0_14866_18608  0.0282587 
iB23_283_v n1_13833_18764 0  0.0282587 
iB23_283_g 0 n0_12896_18777  0.0282587 
iB23_284_v n1_13833_18791 0  0.0282587 
iB23_284_g 0 n0_12896_18777  0.0282587 
iB23_285_v n1_13833_18824 0  0.0282587 
iB23_285_g 0 n0_12896_18810  0.0282587 
iB23_286_v n1_13833_19007 0  0.0282587 
iB23_286_g 0 n0_12896_18993  0.0282587 
iB23_287_v n1_13833_19040 0  0.0282587 
iB23_287_g 0 n0_12896_19026  0.0282587 
iB23_288_v n1_14021_18764 0  0.0282587 
iB23_288_g 0 n0_14866_18777  0.0282587 
iB23_289_v n1_14021_18791 0  0.0282587 
iB23_289_g 0 n0_14866_18777  0.0282587 
iB23_290_v n1_14021_18824 0  0.0282587 
iB23_290_g 0 n0_14866_18810  0.0282587 
iB23_291_v n1_14021_19007 0  0.0282587 
iB23_291_g 0 n0_14866_18993  0.0282587 
iB23_292_v n1_14021_19040 0  0.0282587 
iB23_292_g 0 n0_14866_19026  0.0282587 
iB23_293_v n1_14114_18764 0  0.0282587 
iB23_293_g 0 n0_14866_18777  0.0282587 
iB23_294_v n1_14114_18791 0  0.0282587 
iB23_294_g 0 n0_14866_18777  0.0282587 
iB23_295_v n1_14114_18824 0  0.0282587 
iB23_295_g 0 n0_14866_18810  0.0282587 
iB23_296_v n1_14114_19007 0  0.0282587 
iB23_296_g 0 n0_14866_18993  0.0282587 
iB23_297_v n1_14114_19040 0  0.0282587 
iB23_297_g 0 n0_14866_19026  0.0282587 
iB23_298_v n1_13833_19223 0  0.0282587 
iB23_298_g 0 n0_12896_19209  0.0282587 
iB23_299_v n1_13833_19256 0  0.0282587 
iB23_299_g 0 n0_12896_19256  0.0282587 
iB23_300_v n1_13833_19404 0  0.0282587 
iB23_300_g 0 n0_12896_19425  0.0282587 
iB23_301_v n1_13833_19412 0  0.0282587 
iB23_301_g 0 n0_12896_19425  0.0282587 
iB23_302_v n1_13833_19439 0  0.0282587 
iB23_302_g 0 n0_12896_19425  0.0282587 
iB23_303_v n1_13833_19472 0  0.0282587 
iB23_303_g 0 n0_12896_19458  0.0282587 
iB23_304_v n1_14021_19223 0  0.0282587 
iB23_304_g 0 n0_14866_19209  0.0282587 
iB23_305_v n1_14021_19256 0  0.0282587 
iB23_305_g 0 n0_14866_19256  0.0282587 
iB23_306_v n1_14021_19404 0  0.0282587 
iB23_306_g 0 n0_14866_19425  0.0282587 
iB23_307_v n1_14021_19412 0  0.0282587 
iB23_307_g 0 n0_14866_19425  0.0282587 
iB23_308_v n1_14021_19439 0  0.0282587 
iB23_308_g 0 n0_14866_19425  0.0282587 
iB23_309_v n1_14021_19472 0  0.0282587 
iB23_309_g 0 n0_14866_19458  0.0282587 
iB23_310_v n1_14114_19223 0  0.0282587 
iB23_310_g 0 n0_14866_19209  0.0282587 
iB23_311_v n1_14114_19256 0  0.0282587 
iB23_311_g 0 n0_14866_19256  0.0282587 
iB23_312_v n1_14114_19404 0  0.0282587 
iB23_312_g 0 n0_14866_19425  0.0282587 
iB23_313_v n1_14114_19439 0  0.0282587 
iB23_313_g 0 n0_14866_19425  0.0282587 
iB23_314_v n1_14114_19472 0  0.0282587 
iB23_314_g 0 n0_14866_19458  0.0282587 
iB23_315_v n1_13833_19871 0  0.0282587 
iB23_315_g 0 n0_12896_19857  0.0282587 
iB23_316_v n1_13833_19904 0  0.0282587 
iB23_316_g 0 n0_12896_19890  0.0282587 
iB23_317_v n1_14021_19655 0  0.0282587 
iB23_317_g 0 n0_14866_19641  0.0282587 
iB23_318_v n1_14021_19688 0  0.0282587 
iB23_318_g 0 n0_14866_19674  0.0282587 
iB23_319_v n1_14021_19871 0  0.0282587 
iB23_319_g 0 n0_14866_19857  0.0282587 
iB23_320_v n1_14021_19904 0  0.0282587 
iB23_320_g 0 n0_14866_19890  0.0282587 
iB23_321_v n1_14114_19655 0  0.0282587 
iB23_321_g 0 n0_14866_19641  0.0282587 
iB23_322_v n1_14114_19688 0  0.0282587 
iB23_322_g 0 n0_14866_19674  0.0282587 
iB23_323_v n1_14114_19871 0  0.0282587 
iB23_323_g 0 n0_14866_19857  0.0282587 
iB23_324_v n1_14114_19904 0  0.0282587 
iB23_324_g 0 n0_14866_19890  0.0282587 
iB23_325_v n1_13833_20087 0  0.0282587 
iB23_325_g 0 n0_12896_20073  0.0282587 
iB23_326_v n1_13833_20120 0  0.0282587 
iB23_326_g 0 n0_12896_20106  0.0282587 
iB23_327_v n1_13833_20303 0  0.0282587 
iB23_327_g 0 n0_12896_20289  0.0282587 
iB23_328_v n1_13833_20336 0  0.0282587 
iB23_328_g 0 n0_12896_20322  0.0282587 
iB23_329_v n1_14021_20087 0  0.0282587 
iB23_329_g 0 n0_14866_20073  0.0282587 
iB23_330_v n1_14021_20120 0  0.0282587 
iB23_330_g 0 n0_14866_20106  0.0282587 
iB23_331_v n1_14021_20303 0  0.0282587 
iB23_331_g 0 n0_14866_20289  0.0282587 
iB23_332_v n1_14021_20336 0  0.0282587 
iB23_332_g 0 n0_14866_20322  0.0282587 
iB23_333_v n1_14114_20087 0  0.0282587 
iB23_333_g 0 n0_14866_20073  0.0282587 
iB23_334_v n1_14114_20120 0  0.0282587 
iB23_334_g 0 n0_14866_20106  0.0282587 
iB23_335_v n1_14114_20303 0  0.0282587 
iB23_335_g 0 n0_14866_20289  0.0282587 
iB23_336_v n1_14114_20336 0  0.0282587 
iB23_336_g 0 n0_14866_20322  0.0282587 
iB23_337_v n1_13833_20519 0  0.0282587 
iB23_337_g 0 n0_12896_20505  0.0282587 
iB23_338_v n1_13833_20552 0  0.0282587 
iB23_338_g 0 n0_12896_20538  0.0282587 
iB23_339_v n1_13833_20687 0  0.0282587 
iB23_339_g 0 n0_12896_20754  0.0282587 
iB23_340_v n1_13833_20735 0  0.0282587 
iB23_340_g 0 n0_12896_20754  0.0282587 
iB23_341_v n1_13833_20768 0  0.0282587 
iB23_341_g 0 n0_12896_20754  0.0282587 
iB23_342_v n1_13880_20687 0  0.0282587 
iB23_342_g 0 n0_12896_20754  0.0282587 
iB23_343_v n1_13880_20735 0  0.0282587 
iB23_343_g 0 n0_12896_20754  0.0282587 
iB23_344_v n1_13880_20768 0  0.0282587 
iB23_344_g 0 n0_12896_20754  0.0282587 
iB23_345_v n1_14021_20519 0  0.0282587 
iB23_345_g 0 n0_14866_20505  0.0282587 
iB23_346_v n1_14021_20552 0  0.0282587 
iB23_346_g 0 n0_14866_20538  0.0282587 
iB23_347_v n1_14021_20687 0  0.0282587 
iB23_347_g 0 n0_14866_20754  0.0282587 
iB23_348_v n1_14021_20768 0  0.0282587 
iB23_348_g 0 n0_14866_20754  0.0282587 
iB23_349_v n1_14114_20519 0  0.0282587 
iB23_349_g 0 n0_14866_20505  0.0282587 
iB23_350_v n1_14114_20552 0  0.0282587 
iB23_350_g 0 n0_14866_20538  0.0282587 
iB23_351_v n1_14114_20687 0  0.0282587 
iB23_351_g 0 n0_14866_20754  0.0282587 
iB23_352_v n1_14114_20735 0  0.0282587 
iB23_352_g 0 n0_14866_20754  0.0282587 
iB23_353_v n1_14114_20768 0  0.0282587 
iB23_353_g 0 n0_14866_20754  0.0282587 
iB23_354_v n1_13833_20951 0  0.0282587 
iB23_354_g 0 n0_12896_20937  0.0282587 
iB23_355_v n1_13833_20984 0  0.0282587 
iB23_355_g 0 n0_12896_20970  0.0282587 
iB23_356_v n1_14021_20951 0  0.0282587 
iB23_356_g 0 n0_14866_20937  0.0282587 
iB23_357_v n1_14021_20984 0  0.0282587 
iB23_357_g 0 n0_14866_20970  0.0282587 
iB23_358_v n1_14114_20951 0  0.0282587 
iB23_358_g 0 n0_14866_20937  0.0282587 
iB23_359_v n1_14114_20984 0  0.0282587 
iB23_359_g 0 n0_14866_20970  0.0282587 
iB23_360_v n1_15900_18527 0  0.0282587 
iB23_360_g 0 n0_15146_18561  0.0282587 
iB23_361_v n1_15900_18575 0  0.0282587 
iB23_361_g 0 n0_15146_18561  0.0282587 
iB23_362_v n1_15900_18608 0  0.0282587 
iB23_362_g 0 n0_15146_18608  0.0282587 
iB23_363_v n1_15900_18764 0  0.0282587 
iB23_363_g 0 n0_15146_18777  0.0282587 
iB23_364_v n1_15900_18791 0  0.0282587 
iB23_364_g 0 n0_15146_18777  0.0282587 
iB23_365_v n1_15900_18824 0  0.0282587 
iB23_365_g 0 n0_15146_18810  0.0282587 
iB23_366_v n1_15900_19007 0  0.0282587 
iB23_366_g 0 n0_15146_18993  0.0282587 
iB23_367_v n1_15900_19040 0  0.0282587 
iB23_367_g 0 n0_15146_19026  0.0282587 
iB23_368_v n1_15900_19223 0  0.0282587 
iB23_368_g 0 n0_15146_19209  0.0282587 
iB23_369_v n1_15900_19256 0  0.0282587 
iB23_369_g 0 n0_15146_19256  0.0282587 
iB23_370_v n1_15900_19412 0  0.0282587 
iB23_370_g 0 n0_15146_19425  0.0282587 
iB23_371_v n1_15900_19439 0  0.0282587 
iB23_371_g 0 n0_15146_19425  0.0282587 
iB23_372_v n1_15900_19472 0  0.0282587 
iB23_372_g 0 n0_15146_19458  0.0282587 
iB23_373_v n1_15900_19655 0  0.0282587 
iB23_373_g 0 n0_15146_19641  0.0282587 
iB23_374_v n1_15900_19688 0  0.0282587 
iB23_374_g 0 n0_15146_19674  0.0282587 
iB23_375_v n1_15900_19871 0  0.0282587 
iB23_375_g 0 n0_15146_19857  0.0282587 
iB23_376_v n1_15900_19904 0  0.0282587 
iB23_376_g 0 n0_15146_19890  0.0282587 
iB23_377_v n1_15900_20087 0  0.0282587 
iB23_377_g 0 n0_15146_20073  0.0282587 
iB23_378_v n1_15900_20120 0  0.0282587 
iB23_378_g 0 n0_15146_20106  0.0282587 
iB23_379_v n1_15900_20303 0  0.0282587 
iB23_379_g 0 n0_15146_20289  0.0282587 
iB23_380_v n1_15900_20336 0  0.0282587 
iB23_380_g 0 n0_15146_20322  0.0282587 
iB23_381_v n1_15900_20519 0  0.0282587 
iB23_381_g 0 n0_15146_20505  0.0282587 
iB23_382_v n1_15900_20552 0  0.0282587 
iB23_382_g 0 n0_15146_20538  0.0282587 
iB23_383_v n1_15900_20687 0  0.0282587 
iB23_383_g 0 n0_15146_20754  0.0282587 
iB23_384_v n1_15900_20735 0  0.0282587 
iB23_384_g 0 n0_15146_20754  0.0282587 
iB23_385_v n1_15900_20768 0  0.0282587 
iB23_385_g 0 n0_15146_20754  0.0282587 
iB23_386_v n1_15900_20951 0  0.0282587 
iB23_386_g 0 n0_15146_20937  0.0282587 
iB23_387_v n1_15900_20984 0  0.0282587 
iB23_387_g 0 n0_15146_20970  0.0282587 
iB10_0_v n1_6900_215 0  0.0186858 
iB10_0_g 0 n0_6146_201  0.0186858 
iB10_1_v n1_6900_248 0  0.0186858 
iB10_1_g 0 n0_6146_234  0.0186858 
iB10_2_v n1_6900_383 0  0.0186858 
iB10_2_g 0 n0_6146_356  0.0186858 
iB10_3_v n1_6900_431 0  0.0186858 
iB10_3_g 0 n0_6146_417  0.0186858 
iB10_4_v n1_6900_464 0  0.0186858 
iB10_4_g 0 n0_6146_450  0.0186858 
iB10_5_v n1_6900_647 0  0.0186858 
iB10_5_g 0 n0_6146_633  0.0186858 
iB10_6_v n1_6900_680 0  0.0186858 
iB10_6_g 0 n0_6146_666  0.0186858 
iB10_7_v n1_6900_863 0  0.0186858 
iB10_7_g 0 n0_6146_849  0.0186858 
iB10_8_v n1_6900_896 0  0.0186858 
iB10_8_g 0 n0_6146_882  0.0186858 
iB10_9_v n1_6900_1079 0  0.0186858 
iB10_9_g 0 n0_6146_1065  0.0186858 
iB10_10_v n1_6900_1112 0  0.0186858 
iB10_10_g 0 n0_6146_1098  0.0186858 
iB10_11_v n1_6900_1295 0  0.0186858 
iB10_11_g 0 n0_6146_1281  0.0186858 
iB10_12_v n1_6900_1328 0  0.0186858 
iB10_12_g 0 n0_6146_1314  0.0186858 
iB10_13_v n1_6900_1511 0  0.0186858 
iB10_13_g 0 n0_6146_1497  0.0186858 
iB10_14_v n1_6900_1544 0  0.0186858 
iB10_14_g 0 n0_6146_1530  0.0186858 
iB10_15_v n1_6900_1727 0  0.0186858 
iB10_15_g 0 n0_6146_1713  0.0186858 
iB10_16_v n1_6900_1760 0  0.0186858 
iB10_16_g 0 n0_6146_1760  0.0186858 
iB10_17_v n1_6900_1916 0  0.0186858 
iB10_17_g 0 n0_6146_1929  0.0186858 
iB10_18_v n1_6900_1943 0  0.0186858 
iB10_18_g 0 n0_6146_1929  0.0186858 
iB10_19_v n1_6900_1976 0  0.0186858 
iB10_19_g 0 n0_6146_1962  0.0186858 
iB10_20_v n1_6900_2159 0  0.0186858 
iB10_20_g 0 n0_6146_2145  0.0186858 
iB10_21_v n1_6900_2192 0  0.0186858 
iB10_21_g 0 n0_6146_2178  0.0186858 
iB10_22_v n1_6900_2375 0  0.0186858 
iB10_22_g 0 n0_6146_2361  0.0186858 
iB10_23_v n1_6900_2408 0  0.0186858 
iB10_23_g 0 n0_6146_2408  0.0186858 
iB10_24_v n1_6900_2543 0  0.0186858 
iB10_24_g 0 n0_6146_2577  0.0186858 
iB10_25_v n1_6900_2564 0  0.0186858 
iB10_25_g 0 n0_6146_2577  0.0186858 
iB10_26_v n1_6900_2591 0  0.0186858 
iB10_26_g 0 n0_6146_2577  0.0186858 
iB10_27_v n1_6900_2624 0  0.0186858 
iB10_27_g 0 n0_6146_2610  0.0186858 
iB10_28_v n1_7083_215 0  0.0186858 
iB10_28_g 0 n0_6146_201  0.0186858 
iB10_29_v n1_7083_248 0  0.0186858 
iB10_29_g 0 n0_6146_234  0.0186858 
iB10_30_v n1_7083_383 0  0.0186858 
iB10_30_g 0 n0_6146_356  0.0186858 
iB10_31_v n1_7271_215 0  0.0186858 
iB10_31_g 0 n0_8116_201  0.0186858 
iB10_32_v n1_7271_248 0  0.0186858 
iB10_32_g 0 n0_8116_234  0.0186858 
iB10_33_v n1_7271_383 0  0.0186858 
iB10_33_g 0 n0_8116_417  0.0186858 
iB10_34_v n1_7083_431 0  0.0186858 
iB10_34_g 0 n0_6146_417  0.0186858 
iB10_35_v n1_7083_464 0  0.0186858 
iB10_35_g 0 n0_6146_450  0.0186858 
iB10_36_v n1_7083_647 0  0.0186858 
iB10_36_g 0 n0_6146_633  0.0186858 
iB10_37_v n1_7083_680 0  0.0186858 
iB10_37_g 0 n0_6146_666  0.0186858 
iB10_38_v n1_7130_431 0  0.0186858 
iB10_38_g 0 n0_6146_417  0.0186858 
iB10_39_v n1_7130_464 0  0.0186858 
iB10_39_g 0 n0_6146_450  0.0186858 
iB10_40_v n1_7271_431 0  0.0186858 
iB10_40_g 0 n0_8116_417  0.0186858 
iB10_41_v n1_7271_647 0  0.0186858 
iB10_41_g 0 n0_8116_633  0.0186858 
iB10_42_v n1_7271_680 0  0.0186858 
iB10_42_g 0 n0_8116_666  0.0186858 
iB10_43_v n1_7083_863 0  0.0186858 
iB10_43_g 0 n0_6146_849  0.0186858 
iB10_44_v n1_7083_896 0  0.0186858 
iB10_44_g 0 n0_6146_882  0.0186858 
iB10_45_v n1_7083_1079 0  0.0186858 
iB10_45_g 0 n0_6146_1065  0.0186858 
iB10_46_v n1_7083_1112 0  0.0186858 
iB10_46_g 0 n0_6146_1098  0.0186858 
iB10_47_v n1_7271_863 0  0.0186858 
iB10_47_g 0 n0_8116_849  0.0186858 
iB10_48_v n1_7271_896 0  0.0186858 
iB10_48_g 0 n0_8116_882  0.0186858 
iB10_49_v n1_7271_1079 0  0.0186858 
iB10_49_g 0 n0_8116_1065  0.0186858 
iB10_50_v n1_7271_1112 0  0.0186858 
iB10_50_g 0 n0_8116_1098  0.0186858 
iB10_51_v n1_7083_1295 0  0.0186858 
iB10_51_g 0 n0_6146_1281  0.0186858 
iB10_52_v n1_7083_1328 0  0.0186858 
iB10_52_g 0 n0_6146_1314  0.0186858 
iB10_53_v n1_7271_1295 0  0.0186858 
iB10_53_g 0 n0_8116_1281  0.0186858 
iB10_54_v n1_7271_1328 0  0.0186858 
iB10_54_g 0 n0_8116_1314  0.0186858 
iB10_55_v n1_7271_1511 0  0.0186858 
iB10_55_g 0 n0_8116_1497  0.0186858 
iB10_56_v n1_7271_1544 0  0.0186858 
iB10_56_g 0 n0_8116_1530  0.0186858 
iB10_57_v n1_7083_1727 0  0.0186858 
iB10_57_g 0 n0_6146_1713  0.0186858 
iB10_58_v n1_7083_1760 0  0.0186858 
iB10_58_g 0 n0_6146_1760  0.0186858 
iB10_59_v n1_7083_1916 0  0.0186858 
iB10_59_g 0 n0_6146_1929  0.0186858 
iB10_60_v n1_7083_1943 0  0.0186858 
iB10_60_g 0 n0_6146_1929  0.0186858 
iB10_61_v n1_7083_1976 0  0.0186858 
iB10_61_g 0 n0_6146_1962  0.0186858 
iB10_62_v n1_7271_1727 0  0.0186858 
iB10_62_g 0 n0_8116_1713  0.0186858 
iB10_63_v n1_7271_1760 0  0.0186858 
iB10_63_g 0 n0_8116_1760  0.0186858 
iB10_64_v n1_7271_1916 0  0.0186858 
iB10_64_g 0 n0_8116_1929  0.0186858 
iB10_65_v n1_7271_1943 0  0.0186858 
iB10_65_g 0 n0_8116_1929  0.0186858 
iB10_66_v n1_7271_1976 0  0.0186858 
iB10_66_g 0 n0_8116_1962  0.0186858 
iB10_67_v n1_7083_2159 0  0.0186858 
iB10_67_g 0 n0_6146_2145  0.0186858 
iB10_68_v n1_7083_2192 0  0.0186858 
iB10_68_g 0 n0_6146_2178  0.0186858 
iB10_69_v n1_7083_2375 0  0.0186858 
iB10_69_g 0 n0_6146_2361  0.0186858 
iB10_70_v n1_7083_2408 0  0.0186858 
iB10_70_g 0 n0_6146_2408  0.0186858 
iB10_71_v n1_7271_2159 0  0.0186858 
iB10_71_g 0 n0_8116_2145  0.0186858 
iB10_72_v n1_7271_2192 0  0.0186858 
iB10_72_g 0 n0_8116_2178  0.0186858 
iB10_73_v n1_7271_2375 0  0.0186858 
iB10_73_g 0 n0_8116_2361  0.0186858 
iB10_74_v n1_7271_2408 0  0.0186858 
iB10_74_g 0 n0_8116_2408  0.0186858 
iB10_75_v n1_7083_2543 0  0.0186858 
iB10_75_g 0 n0_6146_2577  0.0186858 
iB10_76_v n1_7083_2564 0  0.0186858 
iB10_76_g 0 n0_6146_2577  0.0186858 
iB10_77_v n1_7083_2591 0  0.0186858 
iB10_77_g 0 n0_6146_2577  0.0186858 
iB10_78_v n1_7083_2624 0  0.0186858 
iB10_78_g 0 n0_6146_2610  0.0186858 
iB10_79_v n1_7083_2807 0  0.0186858 
iB10_79_g 0 n0_6146_2793  0.0186858 
iB10_80_v n1_7083_2840 0  0.0186858 
iB10_80_g 0 n0_6146_2840  0.0186858 
iB10_81_v n1_7271_2543 0  0.0186858 
iB10_81_g 0 n0_8116_2577  0.0186858 
iB10_82_v n1_7271_2564 0  0.0186858 
iB10_82_g 0 n0_8116_2577  0.0186858 
iB10_83_v n1_7271_2591 0  0.0186858 
iB10_83_g 0 n0_8116_2577  0.0186858 
iB10_84_v n1_7271_2624 0  0.0186858 
iB10_84_g 0 n0_8116_2610  0.0186858 
iB10_85_v n1_7271_2807 0  0.0186858 
iB10_85_g 0 n0_8116_2793  0.0186858 
iB10_86_v n1_7271_2840 0  0.0186858 
iB10_86_g 0 n0_8116_2840  0.0186858 
iB10_87_v n1_7083_2974 0  0.0186858 
iB10_87_g 0 n0_6146_3009  0.0186858 
iB10_88_v n1_7083_2996 0  0.0186858 
iB10_88_g 0 n0_6146_3009  0.0186858 
iB10_89_v n1_7083_3023 0  0.0186858 
iB10_89_g 0 n0_6146_3009  0.0186858 
iB10_90_v n1_7083_3056 0  0.0186858 
iB10_90_g 0 n0_6146_3056  0.0186858 
iB10_91_v n1_7083_3239 0  0.0186858 
iB10_91_g 0 n0_6146_3225  0.0186858 
iB10_92_v n1_7271_2974 0  0.0186858 
iB10_92_g 0 n0_8116_3009  0.0186858 
iB10_93_v n1_7271_2996 0  0.0186858 
iB10_93_g 0 n0_8116_3009  0.0186858 
iB10_94_v n1_7271_3023 0  0.0186858 
iB10_94_g 0 n0_8116_3009  0.0186858 
iB10_95_v n1_7271_3056 0  0.0186858 
iB10_95_g 0 n0_8116_3042  0.0186858 
iB10_96_v n1_7271_3239 0  0.0186858 
iB10_96_g 0 n0_8116_3225  0.0186858 
iB10_97_v n1_7083_3272 0  0.0186858 
iB10_97_g 0 n0_6146_3258  0.0186858 
iB10_98_v n1_7083_3455 0  0.0186858 
iB10_98_g 0 n0_6146_3441  0.0186858 
iB10_99_v n1_7083_3488 0  0.0186858 
iB10_99_g 0 n0_6146_3488  0.0186858 
iB10_100_v n1_7083_3644 0  0.0186858 
iB10_100_g 0 n0_6146_3657  0.0186858 
iB10_101_v n1_7083_3671 0  0.0186858 
iB10_101_g 0 n0_6146_3657  0.0186858 
iB10_102_v n1_7271_3272 0  0.0186858 
iB10_102_g 0 n0_8116_3258  0.0186858 
iB10_103_v n1_7271_3455 0  0.0186858 
iB10_103_g 0 n0_8116_3441  0.0186858 
iB10_104_v n1_7271_3488 0  0.0186858 
iB10_104_g 0 n0_8116_3488  0.0186858 
iB10_105_v n1_7271_3644 0  0.0186858 
iB10_105_g 0 n0_8116_3657  0.0186858 
iB10_106_v n1_7271_3671 0  0.0186858 
iB10_106_g 0 n0_8116_3657  0.0186858 
iB10_107_v n1_7083_3704 0  0.0186858 
iB10_107_g 0 n0_6146_3690  0.0186858 
iB10_108_v n1_7271_3704 0  0.0186858 
iB10_108_g 0 n0_8116_3690  0.0186858 
iB10_109_v n1_7271_3887 0  0.0186858 
iB10_109_g 0 n0_8116_3873  0.0186858 
iB10_110_v n1_7271_3920 0  0.0186858 
iB10_110_g 0 n0_8116_3906  0.0186858 
iB10_111_v n1_7083_4103 0  0.0186858 
iB10_111_g 0 n0_6146_4089  0.0186858 
iB10_112_v n1_7083_4136 0  0.0186858 
iB10_112_g 0 n0_6146_4136  0.0186858 
iB10_113_v n1_7083_4292 0  0.0186858 
iB10_113_g 0 n0_6146_4305  0.0186858 
iB10_114_v n1_7083_4319 0  0.0186858 
iB10_114_g 0 n0_6146_4305  0.0186858 
iB10_115_v n1_7083_4352 0  0.0186858 
iB10_115_g 0 n0_6146_4352  0.0186858 
iB10_116_v n1_7271_4103 0  0.0186858 
iB10_116_g 0 n0_8116_4089  0.0186858 
iB10_117_v n1_7271_4136 0  0.0186858 
iB10_117_g 0 n0_8116_4136  0.0186858 
iB10_118_v n1_7271_4292 0  0.0186858 
iB10_118_g 0 n0_8116_4305  0.0186858 
iB10_119_v n1_7271_4319 0  0.0186858 
iB10_119_g 0 n0_8116_4305  0.0186858 
iB10_120_v n1_7271_4352 0  0.0186858 
iB10_120_g 0 n0_8116_4338  0.0186858 
iB10_121_v n1_7083_4535 0  0.0186858 
iB10_121_g 0 n0_6146_4521  0.0186858 
iB10_122_v n1_7083_4568 0  0.0186858 
iB10_122_g 0 n0_6146_4568  0.0186858 
iB10_123_v n1_7083_4724 0  0.0186858 
iB10_123_g 0 n0_6146_4737  0.0186858 
iB10_124_v n1_7083_4751 0  0.0186858 
iB10_124_g 0 n0_6146_4737  0.0186858 
iB10_125_v n1_7083_4784 0  0.0186858 
iB10_125_g 0 n0_6146_4770  0.0186858 
iB10_126_v n1_7271_4535 0  0.0186858 
iB10_126_g 0 n0_8116_4521  0.0186858 
iB10_127_v n1_7271_4568 0  0.0186858 
iB10_127_g 0 n0_8116_4568  0.0186858 
iB10_128_v n1_7271_4724 0  0.0186858 
iB10_128_g 0 n0_8116_4737  0.0186858 
iB10_129_v n1_7271_4751 0  0.0186858 
iB10_129_g 0 n0_8116_4737  0.0186858 
iB10_130_v n1_7271_4784 0  0.0186858 
iB10_130_g 0 n0_8116_4770  0.0186858 
iB10_131_v n1_7083_4967 0  0.0186858 
iB10_131_g 0 n0_6146_4953  0.0186858 
iB10_132_v n1_7083_5000 0  0.0186858 
iB10_132_g 0 n0_6146_4953  0.0186858 
iB10_133_v n1_7083_5183 0  0.0186858 
iB10_133_g 0 n0_6146_5169  0.0186858 
iB10_134_v n1_7083_5216 0  0.0186858 
iB10_134_g 0 n0_6146_5216  0.0186858 
iB10_135_v n1_7130_4967 0  0.0186858 
iB10_135_g 0 n0_6146_4953  0.0186858 
iB10_136_v n1_7130_5000 0  0.0186858 
iB10_136_g 0 n0_6146_4953  0.0186858 
iB10_137_v n1_7271_5000 0  0.0186858 
iB10_137_g 0 n0_8116_4953  0.0186858 
iB10_138_v n1_7271_5183 0  0.0186858 
iB10_138_g 0 n0_8116_5169  0.0186858 
iB10_139_v n1_7271_5216 0  0.0186858 
iB10_139_g 0 n0_8116_5216  0.0186858 
iB10_140_v n1_7364_215 0  0.0186858 
iB10_140_g 0 n0_8116_201  0.0186858 
iB10_141_v n1_7364_248 0  0.0186858 
iB10_141_g 0 n0_8116_234  0.0186858 
iB10_142_v n1_7364_383 0  0.0186858 
iB10_142_g 0 n0_8116_417  0.0186858 
iB10_143_v n1_7364_431 0  0.0186858 
iB10_143_g 0 n0_8116_417  0.0186858 
iB10_144_v n1_7364_464 0  0.0186858 
iB10_144_g 0 n0_8116_450  0.0186858 
iB10_145_v n1_7364_647 0  0.0186858 
iB10_145_g 0 n0_8116_633  0.0186858 
iB10_146_v n1_7364_680 0  0.0186858 
iB10_146_g 0 n0_8116_666  0.0186858 
iB10_147_v n1_7364_863 0  0.0186858 
iB10_147_g 0 n0_8116_849  0.0186858 
iB10_148_v n1_7364_896 0  0.0186858 
iB10_148_g 0 n0_8116_882  0.0186858 
iB10_149_v n1_7364_1079 0  0.0186858 
iB10_149_g 0 n0_8116_1065  0.0186858 
iB10_150_v n1_7364_1112 0  0.0186858 
iB10_150_g 0 n0_8116_1098  0.0186858 
iB10_151_v n1_7364_1295 0  0.0186858 
iB10_151_g 0 n0_8116_1281  0.0186858 
iB10_152_v n1_7364_1328 0  0.0186858 
iB10_152_g 0 n0_8116_1314  0.0186858 
iB10_153_v n1_7364_1511 0  0.0186858 
iB10_153_g 0 n0_8116_1497  0.0186858 
iB10_154_v n1_7364_1544 0  0.0186858 
iB10_154_g 0 n0_8116_1530  0.0186858 
iB10_155_v n1_7364_1727 0  0.0186858 
iB10_155_g 0 n0_8116_1713  0.0186858 
iB10_156_v n1_7364_1760 0  0.0186858 
iB10_156_g 0 n0_8116_1760  0.0186858 
iB10_157_v n1_7364_1916 0  0.0186858 
iB10_157_g 0 n0_8116_1929  0.0186858 
iB10_158_v n1_7364_1943 0  0.0186858 
iB10_158_g 0 n0_8116_1929  0.0186858 
iB10_159_v n1_7364_1976 0  0.0186858 
iB10_159_g 0 n0_8116_1962  0.0186858 
iB10_160_v n1_7364_2159 0  0.0186858 
iB10_160_g 0 n0_8116_2145  0.0186858 
iB10_161_v n1_7364_2192 0  0.0186858 
iB10_161_g 0 n0_8116_2178  0.0186858 
iB10_162_v n1_7364_2375 0  0.0186858 
iB10_162_g 0 n0_8116_2361  0.0186858 
iB10_163_v n1_7364_2408 0  0.0186858 
iB10_163_g 0 n0_8116_2408  0.0186858 
iB10_164_v n1_7364_2543 0  0.0186858 
iB10_164_g 0 n0_8116_2577  0.0186858 
iB10_165_v n1_7364_2564 0  0.0186858 
iB10_165_g 0 n0_8116_2577  0.0186858 
iB10_166_v n1_7364_2591 0  0.0186858 
iB10_166_g 0 n0_8116_2577  0.0186858 
iB10_167_v n1_7364_2624 0  0.0186858 
iB10_167_g 0 n0_8116_2610  0.0186858 
iB10_168_v n1_9150_215 0  0.0186858 
iB10_168_g 0 n0_8396_201  0.0186858 
iB10_169_v n1_9150_248 0  0.0186858 
iB10_169_g 0 n0_8396_234  0.0186858 
iB10_170_v n1_9150_383 0  0.0186858 
iB10_170_g 0 n0_8396_417  0.0186858 
iB10_171_v n1_9333_215 0  0.0186858 
iB10_171_g 0 n0_8396_201  0.0186858 
iB10_172_v n1_9333_248 0  0.0186858 
iB10_172_g 0 n0_8396_234  0.0186858 
iB10_173_v n1_9333_383 0  0.0186858 
iB10_173_g 0 n0_8396_417  0.0186858 
iB10_174_v n1_9150_431 0  0.0186858 
iB10_174_g 0 n0_8396_417  0.0186858 
iB10_175_v n1_9150_464 0  0.0186858 
iB10_175_g 0 n0_8396_450  0.0186858 
iB10_176_v n1_9150_647 0  0.0186858 
iB10_176_g 0 n0_8396_633  0.0186858 
iB10_177_v n1_9150_680 0  0.0186858 
iB10_177_g 0 n0_8396_666  0.0186858 
iB10_178_v n1_9333_431 0  0.0186858 
iB10_178_g 0 n0_8396_417  0.0186858 
iB10_179_v n1_9333_464 0  0.0186858 
iB10_179_g 0 n0_8396_450  0.0186858 
iB10_180_v n1_9333_647 0  0.0186858 
iB10_180_g 0 n0_8396_633  0.0186858 
iB10_181_v n1_9333_680 0  0.0186858 
iB10_181_g 0 n0_8396_666  0.0186858 
iB10_182_v n1_9150_863 0  0.0186858 
iB10_182_g 0 n0_8396_849  0.0186858 
iB10_183_v n1_9150_896 0  0.0186858 
iB10_183_g 0 n0_8396_882  0.0186858 
iB10_184_v n1_9150_1079 0  0.0186858 
iB10_184_g 0 n0_8396_1065  0.0186858 
iB10_185_v n1_9150_1112 0  0.0186858 
iB10_185_g 0 n0_8396_1098  0.0186858 
iB10_186_v n1_9333_863 0  0.0186858 
iB10_186_g 0 n0_8396_849  0.0186858 
iB10_187_v n1_9333_896 0  0.0186858 
iB10_187_g 0 n0_8396_882  0.0186858 
iB10_188_v n1_9333_1079 0  0.0186858 
iB10_188_g 0 n0_8396_1065  0.0186858 
iB10_189_v n1_9333_1112 0  0.0186858 
iB10_189_g 0 n0_8396_1098  0.0186858 
iB10_190_v n1_9150_1295 0  0.0186858 
iB10_190_g 0 n0_8396_1281  0.0186858 
iB10_191_v n1_9150_1328 0  0.0186858 
iB10_191_g 0 n0_8396_1314  0.0186858 
iB10_192_v n1_9150_1511 0  0.0186858 
iB10_192_g 0 n0_8396_1497  0.0186858 
iB10_193_v n1_9150_1544 0  0.0186858 
iB10_193_g 0 n0_8396_1530  0.0186858 
iB10_194_v n1_9333_1295 0  0.0186858 
iB10_194_g 0 n0_8396_1281  0.0186858 
iB10_195_v n1_9333_1328 0  0.0186858 
iB10_195_g 0 n0_8396_1314  0.0186858 
iB10_196_v n1_9150_1727 0  0.0186858 
iB10_196_g 0 n0_8396_1713  0.0186858 
iB10_197_v n1_9150_1760 0  0.0186858 
iB10_197_g 0 n0_8396_1760  0.0186858 
iB10_198_v n1_9150_1894 0  0.0186858 
iB10_198_g 0 n0_8396_1929  0.0186858 
iB10_199_v n1_9150_1943 0  0.0186858 
iB10_199_g 0 n0_8396_1929  0.0186858 
iB10_200_v n1_9150_1976 0  0.0186858 
iB10_200_g 0 n0_8396_1962  0.0186858 
iB10_201_v n1_9333_1727 0  0.0186858 
iB10_201_g 0 n0_8396_1713  0.0186858 
iB10_202_v n1_9333_1760 0  0.0186858 
iB10_202_g 0 n0_8396_1760  0.0186858 
iB10_203_v n1_9333_1894 0  0.0186858 
iB10_203_g 0 n0_8396_1929  0.0186858 
iB10_204_v n1_9333_1916 0  0.0186858 
iB10_204_g 0 n0_8396_1929  0.0186858 
iB10_205_v n1_9333_1943 0  0.0186858 
iB10_205_g 0 n0_8396_1929  0.0186858 
iB10_206_v n1_9333_1976 0  0.0186858 
iB10_206_g 0 n0_8396_1962  0.0186858 
iB10_207_v n1_9150_2159 0  0.0186858 
iB10_207_g 0 n0_8396_2145  0.0186858 
iB10_208_v n1_9150_2192 0  0.0186858 
iB10_208_g 0 n0_8396_2178  0.0186858 
iB10_209_v n1_9150_2375 0  0.0186858 
iB10_209_g 0 n0_8396_2361  0.0186858 
iB10_210_v n1_9150_2408 0  0.0186858 
iB10_210_g 0 n0_8396_2408  0.0186858 
iB10_211_v n1_9333_2159 0  0.0186858 
iB10_211_g 0 n0_8396_2145  0.0186858 
iB10_212_v n1_9333_2192 0  0.0186858 
iB10_212_g 0 n0_8396_2178  0.0186858 
iB10_213_v n1_9333_2375 0  0.0186858 
iB10_213_g 0 n0_8396_2361  0.0186858 
iB10_214_v n1_9333_2408 0  0.0186858 
iB10_214_g 0 n0_8396_2408  0.0186858 
iB10_215_v n1_9150_2543 0  0.0186858 
iB10_215_g 0 n0_8396_2577  0.0186858 
iB10_216_v n1_9150_2564 0  0.0186858 
iB10_216_g 0 n0_8396_2577  0.0186858 
iB10_217_v n1_9150_2591 0  0.0186858 
iB10_217_g 0 n0_8396_2577  0.0186858 
iB10_218_v n1_9150_2624 0  0.0186858 
iB10_218_g 0 n0_8396_2610  0.0186858 
iB10_219_v n1_9333_2543 0  0.0186858 
iB10_219_g 0 n0_8396_2577  0.0186858 
iB10_220_v n1_9333_2564 0  0.0186858 
iB10_220_g 0 n0_8396_2577  0.0186858 
iB10_221_v n1_9333_2591 0  0.0186858 
iB10_221_g 0 n0_8396_2577  0.0186858 
iB10_222_v n1_9333_2624 0  0.0186858 
iB10_222_g 0 n0_8396_2610  0.0186858 
iB10_223_v n1_9333_2807 0  0.0186858 
iB10_223_g 0 n0_8396_2793  0.0186858 
iB10_224_v n1_9333_2840 0  0.0186858 
iB10_224_g 0 n0_8396_2840  0.0186858 
iB10_225_v n1_9333_2996 0  0.0186858 
iB10_225_g 0 n0_8396_3009  0.0186858 
iB10_226_v n1_9333_3023 0  0.0186858 
iB10_226_g 0 n0_8396_3009  0.0186858 
iB10_227_v n1_9333_3056 0  0.0186858 
iB10_227_g 0 n0_8396_3042  0.0186858 
iB10_228_v n1_9333_3239 0  0.0186858 
iB10_228_g 0 n0_8396_3225  0.0186858 
iB10_229_v n1_9333_3272 0  0.0186858 
iB10_229_g 0 n0_8396_3258  0.0186858 
iB10_230_v n1_9333_3455 0  0.0186858 
iB10_230_g 0 n0_8396_3441  0.0186858 
iB10_231_v n1_9333_3488 0  0.0186858 
iB10_231_g 0 n0_8396_3488  0.0186858 
iB10_232_v n1_9333_3644 0  0.0186858 
iB10_232_g 0 n0_8396_3657  0.0186858 
iB10_233_v n1_9333_3671 0  0.0186858 
iB10_233_g 0 n0_8396_3657  0.0186858 
iB10_234_v n1_9333_3704 0  0.0186858 
iB10_234_g 0 n0_8396_3690  0.0186858 
iB10_235_v n1_9333_4103 0  0.0186858 
iB10_235_g 0 n0_8396_4089  0.0186858 
iB10_236_v n1_9333_4136 0  0.0186858 
iB10_236_g 0 n0_8396_4136  0.0186858 
iB10_237_v n1_9333_4292 0  0.0186858 
iB10_237_g 0 n0_8396_4305  0.0186858 
iB10_238_v n1_9333_4319 0  0.0186858 
iB10_238_g 0 n0_8396_4305  0.0186858 
iB10_239_v n1_9333_4352 0  0.0186858 
iB10_239_g 0 n0_8396_4338  0.0186858 
iB10_240_v n1_9333_4535 0  0.0186858 
iB10_240_g 0 n0_8396_4521  0.0186858 
iB10_241_v n1_9333_4568 0  0.0186858 
iB10_241_g 0 n0_8396_4568  0.0186858 
iB10_242_v n1_9333_4724 0  0.0186858 
iB10_242_g 0 n0_8396_4737  0.0186858 
iB10_243_v n1_9333_4751 0  0.0186858 
iB10_243_g 0 n0_8396_4737  0.0186858 
iB10_244_v n1_9333_4784 0  0.0186858 
iB10_244_g 0 n0_8396_4770  0.0186858 
iB10_245_v n1_9333_4967 0  0.0186858 
iB10_245_g 0 n0_8396_4953  0.0186858 
iB10_246_v n1_9333_5000 0  0.0186858 
iB10_246_g 0 n0_8396_4953  0.0186858 
iB10_247_v n1_9333_5183 0  0.0186858 
iB10_247_g 0 n0_8396_5169  0.0186858 
iB10_248_v n1_9333_5216 0  0.0186858 
iB10_248_g 0 n0_8396_5216  0.0186858 
iB10_249_v n1_9521_215 0  0.0186858 
iB10_249_g 0 n0_10366_201  0.0186858 
iB10_250_v n1_9521_248 0  0.0186858 
iB10_250_g 0 n0_10366_234  0.0186858 
iB10_251_v n1_9521_383 0  0.0186858 
iB10_251_g 0 n0_10366_417  0.0186858 
iB10_252_v n1_9614_215 0  0.0186858 
iB10_252_g 0 n0_10366_201  0.0186858 
iB10_253_v n1_9614_248 0  0.0186858 
iB10_253_g 0 n0_10366_234  0.0186858 
iB10_254_v n1_9614_383 0  0.0186858 
iB10_254_g 0 n0_10366_417  0.0186858 
iB10_255_v n1_9380_431 0  0.0186858 
iB10_255_g 0 n0_8396_417  0.0186858 
iB10_256_v n1_9380_464 0  0.0186858 
iB10_256_g 0 n0_8396_450  0.0186858 
iB10_257_v n1_9521_431 0  0.0186858 
iB10_257_g 0 n0_10366_417  0.0186858 
iB10_258_v n1_9521_647 0  0.0186858 
iB10_258_g 0 n0_10366_633  0.0186858 
iB10_259_v n1_9521_680 0  0.0186858 
iB10_259_g 0 n0_10366_666  0.0186858 
iB10_260_v n1_9614_431 0  0.0186858 
iB10_260_g 0 n0_10366_417  0.0186858 
iB10_261_v n1_9614_464 0  0.0186858 
iB10_261_g 0 n0_10366_450  0.0186858 
iB10_262_v n1_9614_647 0  0.0186858 
iB10_262_g 0 n0_10366_633  0.0186858 
iB10_263_v n1_9614_680 0  0.0186858 
iB10_263_g 0 n0_10366_666  0.0186858 
iB10_264_v n1_9521_863 0  0.0186858 
iB10_264_g 0 n0_10366_849  0.0186858 
iB10_265_v n1_9521_896 0  0.0186858 
iB10_265_g 0 n0_10366_882  0.0186858 
iB10_266_v n1_9521_1079 0  0.0186858 
iB10_266_g 0 n0_10366_1065  0.0186858 
iB10_267_v n1_9521_1112 0  0.0186858 
iB10_267_g 0 n0_10366_1098  0.0186858 
iB10_268_v n1_9614_863 0  0.0186858 
iB10_268_g 0 n0_10366_849  0.0186858 
iB10_269_v n1_9614_896 0  0.0186858 
iB10_269_g 0 n0_10366_882  0.0186858 
iB10_270_v n1_9614_1079 0  0.0186858 
iB10_270_g 0 n0_10366_1065  0.0186858 
iB10_271_v n1_9614_1112 0  0.0186858 
iB10_271_g 0 n0_10366_1098  0.0186858 
iB10_272_v n1_9521_1295 0  0.0186858 
iB10_272_g 0 n0_10366_1281  0.0186858 
iB10_273_v n1_9521_1328 0  0.0186858 
iB10_273_g 0 n0_10366_1314  0.0186858 
iB10_274_v n1_9521_1511 0  0.0186858 
iB10_274_g 0 n0_10366_1497  0.0186858 
iB10_275_v n1_9521_1544 0  0.0186858 
iB10_275_g 0 n0_10366_1530  0.0186858 
iB10_276_v n1_9614_1295 0  0.0186858 
iB10_276_g 0 n0_10366_1281  0.0186858 
iB10_277_v n1_9614_1328 0  0.0186858 
iB10_277_g 0 n0_10366_1314  0.0186858 
iB10_278_v n1_9614_1511 0  0.0186858 
iB10_278_g 0 n0_10366_1497  0.0186858 
iB10_279_v n1_9614_1544 0  0.0186858 
iB10_279_g 0 n0_10366_1530  0.0186858 
iB10_280_v n1_9521_1727 0  0.0186858 
iB10_280_g 0 n0_10366_1713  0.0186858 
iB10_281_v n1_9521_1760 0  0.0186858 
iB10_281_g 0 n0_10366_1760  0.0186858 
iB10_282_v n1_9521_1894 0  0.0186858 
iB10_282_g 0 n0_10366_1929  0.0186858 
iB10_283_v n1_9521_1916 0  0.0186858 
iB10_283_g 0 n0_10366_1929  0.0186858 
iB10_284_v n1_9521_1943 0  0.0186858 
iB10_284_g 0 n0_10366_1929  0.0186858 
iB10_285_v n1_9521_1976 0  0.0186858 
iB10_285_g 0 n0_10366_1962  0.0186858 
iB10_286_v n1_9614_1727 0  0.0186858 
iB10_286_g 0 n0_10366_1713  0.0186858 
iB10_287_v n1_9614_1760 0  0.0186858 
iB10_287_g 0 n0_10366_1760  0.0186858 
iB10_288_v n1_9614_1916 0  0.0186858 
iB10_288_g 0 n0_10366_1929  0.0186858 
iB10_289_v n1_9614_1943 0  0.0186858 
iB10_289_g 0 n0_10366_1929  0.0186858 
iB10_290_v n1_9614_1976 0  0.0186858 
iB10_290_g 0 n0_10366_1962  0.0186858 
iB10_291_v n1_9521_2159 0  0.0186858 
iB10_291_g 0 n0_10366_2145  0.0186858 
iB10_292_v n1_9521_2192 0  0.0186858 
iB10_292_g 0 n0_10366_2178  0.0186858 
iB10_293_v n1_9521_2375 0  0.0186858 
iB10_293_g 0 n0_10366_2361  0.0186858 
iB10_294_v n1_9521_2408 0  0.0186858 
iB10_294_g 0 n0_10366_2408  0.0186858 
iB10_295_v n1_9614_2159 0  0.0186858 
iB10_295_g 0 n0_10366_2145  0.0186858 
iB10_296_v n1_9614_2192 0  0.0186858 
iB10_296_g 0 n0_10366_2178  0.0186858 
iB10_297_v n1_9614_2375 0  0.0186858 
iB10_297_g 0 n0_10366_2361  0.0186858 
iB10_298_v n1_9614_2408 0  0.0186858 
iB10_298_g 0 n0_10366_2408  0.0186858 
iB10_299_v n1_9521_2543 0  0.0186858 
iB10_299_g 0 n0_10366_2577  0.0186858 
iB10_300_v n1_9521_2564 0  0.0186858 
iB10_300_g 0 n0_10366_2577  0.0186858 
iB10_301_v n1_9521_2591 0  0.0186858 
iB10_301_g 0 n0_10366_2577  0.0186858 
iB10_302_v n1_9521_2624 0  0.0186858 
iB10_302_g 0 n0_10366_2610  0.0186858 
iB10_303_v n1_9521_2807 0  0.0186858 
iB10_303_g 0 n0_10366_2793  0.0186858 
iB10_304_v n1_9521_2840 0  0.0186858 
iB10_304_g 0 n0_10366_2840  0.0186858 
iB10_305_v n1_9614_2543 0  0.0186858 
iB10_305_g 0 n0_10366_2577  0.0186858 
iB10_306_v n1_9614_2564 0  0.0186858 
iB10_306_g 0 n0_10366_2577  0.0186858 
iB10_307_v n1_9614_2591 0  0.0186858 
iB10_307_g 0 n0_10366_2577  0.0186858 
iB10_308_v n1_9614_2624 0  0.0186858 
iB10_308_g 0 n0_10366_2610  0.0186858 
iB10_309_v n1_9521_2996 0  0.0186858 
iB10_309_g 0 n0_10366_3009  0.0186858 
iB10_310_v n1_9521_3023 0  0.0186858 
iB10_310_g 0 n0_10366_3009  0.0186858 
iB10_311_v n1_9521_3056 0  0.0186858 
iB10_311_g 0 n0_10366_3042  0.0186858 
iB10_312_v n1_9521_3239 0  0.0186858 
iB10_312_g 0 n0_10366_3225  0.0186858 
iB10_313_v n1_9521_3272 0  0.0186858 
iB10_313_g 0 n0_10366_3258  0.0186858 
iB10_314_v n1_9521_3455 0  0.0186858 
iB10_314_g 0 n0_10366_3441  0.0186858 
iB10_315_v n1_9521_3488 0  0.0186858 
iB10_315_g 0 n0_10366_3488  0.0186858 
iB10_316_v n1_9521_3644 0  0.0186858 
iB10_316_g 0 n0_10366_3657  0.0186858 
iB10_317_v n1_9521_3671 0  0.0186858 
iB10_317_g 0 n0_10366_3657  0.0186858 
iB10_318_v n1_9521_3704 0  0.0186858 
iB10_318_g 0 n0_10366_3690  0.0186858 
iB10_319_v n1_9521_3887 0  0.0186858 
iB10_319_g 0 n0_10366_3873  0.0186858 
iB10_320_v n1_9521_3920 0  0.0186858 
iB10_320_g 0 n0_10366_3906  0.0186858 
iB10_321_v n1_9521_4103 0  0.0186858 
iB10_321_g 0 n0_10366_4089  0.0186858 
iB10_322_v n1_9521_4136 0  0.0186858 
iB10_322_g 0 n0_10366_4136  0.0186858 
iB10_323_v n1_9521_4292 0  0.0186858 
iB10_323_g 0 n0_10366_4305  0.0186858 
iB10_324_v n1_9521_4319 0  0.0186858 
iB10_324_g 0 n0_10366_4305  0.0186858 
iB10_325_v n1_9521_4352 0  0.0186858 
iB10_325_g 0 n0_10366_4338  0.0186858 
iB10_326_v n1_9521_4535 0  0.0186858 
iB10_326_g 0 n0_10366_4521  0.0186858 
iB10_327_v n1_9521_4568 0  0.0186858 
iB10_327_g 0 n0_10366_4568  0.0186858 
iB10_328_v n1_9521_4724 0  0.0186858 
iB10_328_g 0 n0_10366_4737  0.0186858 
iB10_329_v n1_9521_4751 0  0.0186858 
iB10_329_g 0 n0_10366_4737  0.0186858 
iB10_330_v n1_9521_4784 0  0.0186858 
iB10_330_g 0 n0_10366_4770  0.0186858 
iB10_331_v n1_9380_4967 0  0.0186858 
iB10_331_g 0 n0_8396_4953  0.0186858 
iB10_332_v n1_9380_5000 0  0.0186858 
iB10_332_g 0 n0_8396_4953  0.0186858 
iB10_333_v n1_9521_5000 0  0.0186858 
iB10_333_g 0 n0_10366_4953  0.0186858 
iB10_334_v n1_9521_5183 0  0.0186858 
iB10_334_g 0 n0_10366_5169  0.0186858 
iB10_335_v n1_9521_5216 0  0.0186858 
iB10_335_g 0 n0_10366_5202  0.0186858 
iB11_0_v n1_7083_5372 0  0.0483404 
iB11_0_g 0 n0_6146_5385  0.0483404 
iB11_1_v n1_7083_5399 0  0.0483404 
iB11_1_g 0 n0_6146_5385  0.0483404 
iB11_2_v n1_7083_5432 0  0.0483404 
iB11_2_g 0 n0_6146_5432  0.0483404 
iB11_3_v n1_7083_5566 0  0.0483404 
iB11_3_g 0 n0_6146_5601  0.0483404 
iB11_4_v n1_7083_5588 0  0.0483404 
iB11_4_g 0 n0_6146_5601  0.0483404 
iB11_5_v n1_7083_5615 0  0.0483404 
iB11_5_g 0 n0_6146_5601  0.0483404 
iB11_6_v n1_7083_5648 0  0.0483404 
iB11_6_g 0 n0_6146_5634  0.0483404 
iB11_7_v n1_7271_5372 0  0.0483404 
iB11_7_g 0 n0_8116_5385  0.0483404 
iB11_8_v n1_7271_5399 0  0.0483404 
iB11_8_g 0 n0_8116_5385  0.0483404 
iB11_9_v n1_7271_5432 0  0.0483404 
iB11_9_g 0 n0_8116_5432  0.0483404 
iB11_10_v n1_7271_5566 0  0.0483404 
iB11_10_g 0 n0_8116_5601  0.0483404 
iB11_11_v n1_7271_5588 0  0.0483404 
iB11_11_g 0 n0_8116_5601  0.0483404 
iB11_12_v n1_7271_5615 0  0.0483404 
iB11_12_g 0 n0_8116_5601  0.0483404 
iB11_13_v n1_7271_5648 0  0.0483404 
iB11_13_g 0 n0_8116_5634  0.0483404 
iB11_14_v n1_7083_5831 0  0.0483404 
iB11_14_g 0 n0_6146_5817  0.0483404 
iB11_15_v n1_7083_5864 0  0.0483404 
iB11_15_g 0 n0_6146_5850  0.0483404 
iB11_16_v n1_7271_5831 0  0.0483404 
iB11_16_g 0 n0_8116_5817  0.0483404 
iB11_17_v n1_7271_5864 0  0.0483404 
iB11_17_g 0 n0_8116_5850  0.0483404 
iB11_18_v n1_7271_6047 0  0.0483404 
iB11_18_g 0 n0_8116_6033  0.0483404 
iB11_19_v n1_7271_6080 0  0.0483404 
iB11_19_g 0 n0_8116_6066  0.0483404 
iB11_20_v n1_7083_6263 0  0.0483404 
iB11_20_g 0 n0_8116_6249  0.0483404 
iB11_21_v n1_7083_6296 0  0.0483404 
iB11_21_g 0 n0_8116_6282  0.0483404 
iB11_22_v n1_7083_6479 0  0.0483404 
iB11_22_g 0 n0_6991_7329  0.0483404 
iB11_23_v n1_7083_6512 0  0.0483404 
iB11_23_g 0 n0_6991_7329  0.0483404 
iB11_24_v n1_7271_6263 0  0.0483404 
iB11_24_g 0 n0_8116_6249  0.0483404 
iB11_25_v n1_7271_6296 0  0.0483404 
iB11_25_g 0 n0_8116_6282  0.0483404 
iB11_26_v n1_7271_6479 0  0.0483404 
iB11_26_g 0 n0_7179_7329  0.0483404 
iB11_27_v n1_7271_6512 0  0.0483404 
iB11_27_g 0 n0_7179_7329  0.0483404 
iB11_28_v n1_7083_6646 0  0.0483404 
iB11_28_g 0 n0_6991_7329  0.0483404 
iB11_29_v n1_7083_6695 0  0.0483404 
iB11_29_g 0 n0_6991_7329  0.0483404 
iB11_30_v n1_7083_6728 0  0.0483404 
iB11_30_g 0 n0_6991_7329  0.0483404 
iB11_31_v n1_7083_6911 0  0.0483404 
iB11_31_g 0 n0_6991_7329  0.0483404 
iB11_32_v n1_7271_6646 0  0.0483404 
iB11_32_g 0 n0_7179_7329  0.0483404 
iB11_33_v n1_7271_6695 0  0.0483404 
iB11_33_g 0 n0_7179_7329  0.0483404 
iB11_34_v n1_7271_6728 0  0.0483404 
iB11_34_g 0 n0_7179_7329  0.0483404 
iB11_35_v n1_7271_6911 0  0.0483404 
iB11_35_g 0 n0_7179_7329  0.0483404 
iB11_36_v n1_7083_6944 0  0.0483404 
iB11_36_g 0 n0_6991_7329  0.0483404 
iB11_37_v n1_7083_7127 0  0.0483404 
iB11_37_g 0 n0_6991_7329  0.0483404 
iB11_38_v n1_7083_7160 0  0.0483404 
iB11_38_g 0 n0_6991_7329  0.0483404 
iB11_39_v n1_7130_7160 0  0.0483404 
iB11_39_g 0 n0_7179_7329  0.0483404 
iB11_40_v n1_7271_6944 0  0.0483404 
iB11_40_g 0 n0_7179_7329  0.0483404 
iB11_41_v n1_7271_7127 0  0.0483404 
iB11_41_g 0 n0_7179_7329  0.0483404 
iB11_42_v n1_7271_7160 0  0.0483404 
iB11_42_g 0 n0_7179_7329  0.0483404 
iB11_43_v n1_7083_7343 0  0.0483404 
iB11_43_g 0 n0_6991_7329  0.0483404 
iB11_44_v n1_7083_7376 0  0.0483404 
iB11_44_g 0 n0_6991_7362  0.0483404 
iB11_45_v n1_7083_7559 0  0.0483404 
iB11_45_g 0 n0_6991_7545  0.0483404 
iB11_46_v n1_7083_7592 0  0.0483404 
iB11_46_g 0 n0_6991_7578  0.0483404 
iB11_47_v n1_7271_7343 0  0.0483404 
iB11_47_g 0 n0_7179_7329  0.0483404 
iB11_48_v n1_7271_7376 0  0.0483404 
iB11_48_g 0 n0_7179_7362  0.0483404 
iB11_49_v n1_7271_7559 0  0.0483404 
iB11_49_g 0 n0_7179_7545  0.0483404 
iB11_50_v n1_7271_7592 0  0.0483404 
iB11_50_g 0 n0_7179_7578  0.0483404 
iB11_51_v n1_7083_7775 0  0.0483404 
iB11_51_g 0 n0_6991_7761  0.0483404 
iB11_52_v n1_7083_7808 0  0.0483404 
iB11_52_g 0 n0_6991_7808  0.0483404 
iB11_53_v n1_7083_7822 0  0.0483404 
iB11_53_g 0 n0_6991_7808  0.0483404 
iB11_54_v n1_7083_7964 0  0.0483404 
iB11_54_g 0 n0_6991_7977  0.0483404 
iB11_55_v n1_7083_7991 0  0.0483404 
iB11_55_g 0 n0_6991_7977  0.0483404 
iB11_56_v n1_7083_8024 0  0.0483404 
iB11_56_g 0 n0_6991_8010  0.0483404 
iB11_57_v n1_7271_7775 0  0.0483404 
iB11_57_g 0 n0_7179_7761  0.0483404 
iB11_58_v n1_7271_7808 0  0.0483404 
iB11_58_g 0 n0_7179_7808  0.0483404 
iB11_59_v n1_7271_7822 0  0.0483404 
iB11_59_g 0 n0_7179_7808  0.0483404 
iB11_60_v n1_7271_7964 0  0.0483404 
iB11_60_g 0 n0_7179_7977  0.0483404 
iB11_61_v n1_7271_7991 0  0.0483404 
iB11_61_g 0 n0_7179_7977  0.0483404 
iB11_62_v n1_7271_8024 0  0.0483404 
iB11_62_g 0 n0_7179_8010  0.0483404 
iB11_63_v n1_7083_8207 0  0.0483404 
iB11_63_g 0 n0_6991_8193  0.0483404 
iB11_64_v n1_7083_8240 0  0.0483404 
iB11_64_g 0 n0_6991_8226  0.0483404 
iB11_65_v n1_7083_8456 0  0.0483404 
iB11_65_g 0 n0_7130_8409  0.0483404 
iB11_66_v n1_7271_8207 0  0.0483404 
iB11_66_g 0 n0_7179_8193  0.0483404 
iB11_67_v n1_7271_8240 0  0.0483404 
iB11_67_g 0 n0_7179_8226  0.0483404 
iB11_68_v n1_7271_8423 0  0.0483404 
iB11_68_g 0 n0_7179_8409  0.0483404 
iB11_69_v n1_7271_8456 0  0.0483404 
iB11_69_g 0 n0_7179_8442  0.0483404 
iB11_70_v n1_7083_8639 0  0.0483404 
iB11_70_g 0 n0_6991_8625  0.0483404 
iB11_71_v n1_7083_8672 0  0.0483404 
iB11_71_g 0 n0_6991_8658  0.0483404 
iB11_72_v n1_7083_8855 0  0.0483404 
iB11_72_g 0 n0_6991_8841  0.0483404 
iB11_73_v n1_7083_8888 0  0.0483404 
iB11_73_g 0 n0_6991_8888  0.0483404 
iB11_74_v n1_7083_8902 0  0.0483404 
iB11_74_g 0 n0_6991_8888  0.0483404 
iB11_75_v n1_7271_8639 0  0.0483404 
iB11_75_g 0 n0_7179_8625  0.0483404 
iB11_76_v n1_7271_8672 0  0.0483404 
iB11_76_g 0 n0_7179_8658  0.0483404 
iB11_77_v n1_7271_8855 0  0.0483404 
iB11_77_g 0 n0_7179_8841  0.0483404 
iB11_78_v n1_7271_8888 0  0.0483404 
iB11_78_g 0 n0_7179_8888  0.0483404 
iB11_79_v n1_7271_8902 0  0.0483404 
iB11_79_g 0 n0_7179_8888  0.0483404 
iB11_80_v n1_7083_9044 0  0.0483404 
iB11_80_g 0 n0_6991_9057  0.0483404 
iB11_81_v n1_7083_9071 0  0.0483404 
iB11_81_g 0 n0_6991_9057  0.0483404 
iB11_82_v n1_7083_9104 0  0.0483404 
iB11_82_g 0 n0_6991_9090  0.0483404 
iB11_83_v n1_7083_9287 0  0.0483404 
iB11_83_g 0 n0_6991_9273  0.0483404 
iB11_84_v n1_7083_9320 0  0.0483404 
iB11_84_g 0 n0_6991_9306  0.0483404 
iB11_85_v n1_7271_9044 0  0.0483404 
iB11_85_g 0 n0_7179_9057  0.0483404 
iB11_86_v n1_7271_9071 0  0.0483404 
iB11_86_g 0 n0_7179_9057  0.0483404 
iB11_87_v n1_7271_9104 0  0.0483404 
iB11_87_g 0 n0_7179_9090  0.0483404 
iB11_88_v n1_7271_9287 0  0.0483404 
iB11_88_g 0 n0_7179_9273  0.0483404 
iB11_89_v n1_7271_9320 0  0.0483404 
iB11_89_g 0 n0_7179_9306  0.0483404 
iB11_90_v n1_7083_9503 0  0.0483404 
iB11_90_g 0 n0_6991_9489  0.0483404 
iB11_91_v n1_7083_9536 0  0.0483404 
iB11_91_g 0 n0_6991_9522  0.0483404 
iB11_92_v n1_7083_9719 0  0.0483404 
iB11_92_g 0 n0_6991_9705  0.0483404 
iB11_93_v n1_7083_9752 0  0.0483404 
iB11_93_g 0 n0_6991_9738  0.0483404 
iB11_94_v n1_7130_9503 0  0.0483404 
iB11_94_g 0 n0_6991_9489  0.0483404 
iB11_95_v n1_7130_9536 0  0.0483404 
iB11_95_g 0 n0_6991_9522  0.0483404 
iB11_96_v n1_7271_9503 0  0.0483404 
iB11_96_g 0 n0_7179_9306  0.0483404 
iB11_97_v n1_7271_9536 0  0.0483404 
iB11_97_g 0 n0_7179_9705  0.0483404 
iB11_98_v n1_7271_9719 0  0.0483404 
iB11_98_g 0 n0_7179_9705  0.0483404 
iB11_99_v n1_7271_9752 0  0.0483404 
iB11_99_g 0 n0_7179_9738  0.0483404 
iB11_100_v n1_7083_9935 0  0.0483404 
iB11_100_g 0 n0_6991_9921  0.0483404 
iB11_101_v n1_7083_9968 0  0.0483404 
iB11_101_g 0 n0_6991_9968  0.0483404 
iB11_102_v n1_7083_9982 0  0.0483404 
iB11_102_g 0 n0_6991_9968  0.0483404 
iB11_103_v n1_7083_10124 0  0.0483404 
iB11_103_g 0 n0_6991_10137  0.0483404 
iB11_104_v n1_7083_10151 0  0.0483404 
iB11_104_g 0 n0_6991_10137  0.0483404 
iB11_105_v n1_7083_10184 0  0.0483404 
iB11_105_g 0 n0_6991_10170  0.0483404 
iB11_106_v n1_7271_9935 0  0.0483404 
iB11_106_g 0 n0_7179_9921  0.0483404 
iB11_107_v n1_7271_9968 0  0.0483404 
iB11_107_g 0 n0_7179_9968  0.0483404 
iB11_108_v n1_7271_9982 0  0.0483404 
iB11_108_g 0 n0_7179_9968  0.0483404 
iB11_109_v n1_7271_10124 0  0.0483404 
iB11_109_g 0 n0_7179_10137  0.0483404 
iB11_110_v n1_7271_10151 0  0.0483404 
iB11_110_g 0 n0_7179_10137  0.0483404 
iB11_111_v n1_7271_10184 0  0.0483404 
iB11_111_g 0 n0_7179_10170  0.0483404 
iB11_112_v n1_7083_10367 0  0.0483404 
iB11_112_g 0 n0_6991_10353  0.0483404 
iB11_113_v n1_7083_10400 0  0.0483404 
iB11_113_g 0 n0_6991_10386  0.0483404 
iB11_114_v n1_7271_10367 0  0.0483404 
iB11_114_g 0 n0_7179_10353  0.0483404 
iB11_115_v n1_7271_10400 0  0.0483404 
iB11_115_g 0 n0_7179_10386  0.0483404 
iB11_116_v n1_7271_10616 0  0.0483404 
iB11_116_g 0 n0_7179_10602  0.0483404 
iB11_117_v n1_9333_5350 0  0.0483404 
iB11_117_g 0 n0_8396_5385  0.0483404 
iB11_118_v n1_9333_5372 0  0.0483404 
iB11_118_g 0 n0_8396_5385  0.0483404 
iB11_119_v n1_9333_5399 0  0.0483404 
iB11_119_g 0 n0_8396_5385  0.0483404 
iB11_120_v n1_9333_5432 0  0.0483404 
iB11_120_g 0 n0_8396_5432  0.0483404 
iB11_121_v n1_9333_5588 0  0.0483404 
iB11_121_g 0 n0_8396_5601  0.0483404 
iB11_122_v n1_9333_5615 0  0.0483404 
iB11_122_g 0 n0_8396_5601  0.0483404 
iB11_123_v n1_9333_5648 0  0.0483404 
iB11_123_g 0 n0_8396_5634  0.0483404 
iB11_124_v n1_9333_5831 0  0.0483404 
iB11_124_g 0 n0_8396_5817  0.0483404 
iB11_125_v n1_9333_5864 0  0.0483404 
iB11_125_g 0 n0_8396_5850  0.0483404 
iB11_126_v n1_9333_6263 0  0.0483404 
iB11_126_g 0 n0_8396_6249  0.0483404 
iB11_127_v n1_9333_6296 0  0.0483404 
iB11_127_g 0 n0_8396_6282  0.0483404 
iB11_128_v n1_9333_6479 0  0.0483404 
iB11_128_g 0 n0_8396_6465  0.0483404 
iB11_129_v n1_9333_6512 0  0.0483404 
iB11_129_g 0 n0_8396_6512  0.0483404 
iB11_130_v n1_9333_6668 0  0.0483404 
iB11_130_g 0 n0_8396_6681  0.0483404 
iB11_131_v n1_9333_6695 0  0.0483404 
iB11_131_g 0 n0_8396_6681  0.0483404 
iB11_132_v n1_9333_6728 0  0.0483404 
iB11_132_g 0 n0_8396_6714  0.0483404 
iB11_133_v n1_9333_6911 0  0.0483404 
iB11_133_g 0 n0_8396_6897  0.0483404 
iB11_134_v n1_9333_6944 0  0.0483404 
iB11_134_g 0 n0_8396_6944  0.0483404 
iB11_135_v n1_9333_7100 0  0.0483404 
iB11_135_g 0 n0_8396_7113  0.0483404 
iB11_136_v n1_9333_7127 0  0.0483404 
iB11_136_g 0 n0_8396_7113  0.0483404 
iB11_137_v n1_9333_7160 0  0.0483404 
iB11_137_g 0 n0_8396_7160  0.0483404 
iB11_138_v n1_9333_7316 0  0.0483404 
iB11_138_g 0 n0_8396_7329  0.0483404 
iB11_139_v n1_9333_7343 0  0.0483404 
iB11_139_g 0 n0_8396_7329  0.0483404 
iB11_140_v n1_9333_7376 0  0.0483404 
iB11_140_g 0 n0_8396_7376  0.0483404 
iB11_141_v n1_9333_7532 0  0.0483404 
iB11_141_g 0 n0_8396_7545  0.0483404 
iB11_142_v n1_9333_7559 0  0.0483404 
iB11_142_g 0 n0_8396_7545  0.0483404 
iB11_143_v n1_9333_7592 0  0.0483404 
iB11_143_g 0 n0_8396_7578  0.0483404 
iB11_144_v n1_9333_7775 0  0.0483404 
iB11_144_g 0 n0_8396_7761  0.0483404 
iB11_145_v n1_9333_7808 0  0.0483404 
iB11_145_g 0 n0_8396_7808  0.0483404 
iB11_146_v n1_9333_7991 0  0.0483404 
iB11_146_g 0 n0_8396_7977  0.0483404 
iB11_147_v n1_9333_8024 0  0.0483404 
iB11_147_g 0 n0_8396_8010  0.0483404 
iB11_148_v n1_9333_8207 0  0.0483404 
iB11_148_g 0 n0_8396_8193  0.0483404 
iB11_149_v n1_9333_8240 0  0.0483404 
iB11_149_g 0 n0_8396_8226  0.0483404 
iB11_150_v n1_9333_8456 0  0.0483404 
iB11_150_g 0 n0_8304_8442  0.0483404 
iB11_151_v n1_9333_8639 0  0.0483404 
iB11_151_g 0 n0_9241_9489  0.0483404 
iB11_152_v n1_9333_8672 0  0.0483404 
iB11_152_g 0 n0_9241_9489  0.0483404 
iB11_153_v n1_9333_8855 0  0.0483404 
iB11_153_g 0 n0_9241_9489  0.0483404 
iB11_154_v n1_9333_8888 0  0.0483404 
iB11_154_g 0 n0_9241_9489  0.0483404 
iB11_155_v n1_9333_9071 0  0.0483404 
iB11_155_g 0 n0_9241_9489  0.0483404 
iB11_156_v n1_9333_9104 0  0.0483404 
iB11_156_g 0 n0_9241_9489  0.0483404 
iB11_157_v n1_9333_9287 0  0.0483404 
iB11_157_g 0 n0_9241_9489  0.0483404 
iB11_158_v n1_9333_9320 0  0.0483404 
iB11_158_g 0 n0_9241_9489  0.0483404 
iB11_159_v n1_9333_9503 0  0.0483404 
iB11_159_g 0 n0_9241_9489  0.0483404 
iB11_160_v n1_9333_9536 0  0.0483404 
iB11_160_g 0 n0_9241_9522  0.0483404 
iB11_161_v n1_9333_9719 0  0.0483404 
iB11_161_g 0 n0_9241_9705  0.0483404 
iB11_162_v n1_9333_9752 0  0.0483404 
iB11_162_g 0 n0_9241_9738  0.0483404 
iB11_163_v n1_9333_9935 0  0.0483404 
iB11_163_g 0 n0_9241_9921  0.0483404 
iB11_164_v n1_9333_9968 0  0.0483404 
iB11_164_g 0 n0_9241_9954  0.0483404 
iB11_165_v n1_9333_10151 0  0.0483404 
iB11_165_g 0 n0_9241_10137  0.0483404 
iB11_166_v n1_9333_10184 0  0.0483404 
iB11_166_g 0 n0_9241_10170  0.0483404 
iB11_167_v n1_9333_10367 0  0.0483404 
iB11_167_g 0 n0_9241_10353  0.0483404 
iB11_168_v n1_9333_10400 0  0.0483404 
iB11_168_g 0 n0_9241_10386  0.0483404 
iB11_169_v n1_9521_5350 0  0.0483404 
iB11_169_g 0 n0_10366_5385  0.0483404 
iB11_170_v n1_9521_5372 0  0.0483404 
iB11_170_g 0 n0_10366_5385  0.0483404 
iB11_171_v n1_9521_5399 0  0.0483404 
iB11_171_g 0 n0_10366_5385  0.0483404 
iB11_172_v n1_9521_5432 0  0.0483404 
iB11_172_g 0 n0_10366_5432  0.0483404 
iB11_173_v n1_9521_5588 0  0.0483404 
iB11_173_g 0 n0_10366_5601  0.0483404 
iB11_174_v n1_9521_5615 0  0.0483404 
iB11_174_g 0 n0_10366_5601  0.0483404 
iB11_175_v n1_9521_5648 0  0.0483404 
iB11_175_g 0 n0_10366_5634  0.0483404 
iB11_176_v n1_9521_5831 0  0.0483404 
iB11_176_g 0 n0_10366_5817  0.0483404 
iB11_177_v n1_9521_5864 0  0.0483404 
iB11_177_g 0 n0_10366_5850  0.0483404 
iB11_178_v n1_9521_6047 0  0.0483404 
iB11_178_g 0 n0_10366_6033  0.0483404 
iB11_179_v n1_9521_6080 0  0.0483404 
iB11_179_g 0 n0_10366_6066  0.0483404 
iB11_180_v n1_9521_6263 0  0.0483404 
iB11_180_g 0 n0_10366_6249  0.0483404 
iB11_181_v n1_9521_6296 0  0.0483404 
iB11_181_g 0 n0_10366_6282  0.0483404 
iB11_182_v n1_9521_6479 0  0.0483404 
iB11_182_g 0 n0_10366_6465  0.0483404 
iB11_183_v n1_9521_6512 0  0.0483404 
iB11_183_g 0 n0_10366_6512  0.0483404 
iB11_184_v n1_9521_6668 0  0.0483404 
iB11_184_g 0 n0_10366_6681  0.0483404 
iB11_185_v n1_9521_6695 0  0.0483404 
iB11_185_g 0 n0_10366_6681  0.0483404 
iB11_186_v n1_9521_6728 0  0.0483404 
iB11_186_g 0 n0_10366_6714  0.0483404 
iB11_187_v n1_9521_6911 0  0.0483404 
iB11_187_g 0 n0_10366_6897  0.0483404 
iB11_188_v n1_9380_7160 0  0.0483404 
iB11_188_g 0 n0_8396_7160  0.0483404 
iB11_189_v n1_9521_6944 0  0.0483404 
iB11_189_g 0 n0_10366_6944  0.0483404 
iB11_190_v n1_9521_7100 0  0.0483404 
iB11_190_g 0 n0_10366_7113  0.0483404 
iB11_191_v n1_9521_7127 0  0.0483404 
iB11_191_g 0 n0_10366_7113  0.0483404 
iB11_192_v n1_9521_7160 0  0.0483404 
iB11_192_g 0 n0_10366_7160  0.0483404 
iB11_193_v n1_9521_7316 0  0.0483404 
iB11_193_g 0 n0_10366_7329  0.0483404 
iB11_194_v n1_9521_7343 0  0.0483404 
iB11_194_g 0 n0_10366_7329  0.0483404 
iB11_195_v n1_9521_7376 0  0.0483404 
iB11_195_g 0 n0_10366_7376  0.0483404 
iB11_196_v n1_9521_7532 0  0.0483404 
iB11_196_g 0 n0_10366_7545  0.0483404 
iB11_197_v n1_9521_7559 0  0.0483404 
iB11_197_g 0 n0_10366_7545  0.0483404 
iB11_198_v n1_9521_7592 0  0.0483404 
iB11_198_g 0 n0_10366_7578  0.0483404 
iB11_199_v n1_9521_7775 0  0.0483404 
iB11_199_g 0 n0_10366_7761  0.0483404 
iB11_200_v n1_9521_7808 0  0.0483404 
iB11_200_g 0 n0_10366_7794  0.0483404 
iB11_201_v n1_9521_7991 0  0.0483404 
iB11_201_g 0 n0_10366_7977  0.0483404 
iB11_202_v n1_9521_8024 0  0.0483404 
iB11_202_g 0 n0_10366_8010  0.0483404 
iB11_203_v n1_9521_8207 0  0.0483404 
iB11_203_g 0 n0_10366_8193  0.0483404 
iB11_204_v n1_9521_8240 0  0.0483404 
iB11_204_g 0 n0_10366_8226  0.0483404 
iB11_205_v n1_9521_8423 0  0.0483404 
iB11_205_g 0 n0_10366_8409  0.0483404 
iB11_206_v n1_9521_8456 0  0.0483404 
iB11_206_g 0 n0_10366_8442  0.0483404 
iB11_207_v n1_9521_8639 0  0.0483404 
iB11_207_g 0 n0_10366_8625  0.0483404 
iB11_208_v n1_9521_8672 0  0.0483404 
iB11_208_g 0 n0_10366_8658  0.0483404 
iB11_209_v n1_9521_8855 0  0.0483404 
iB11_209_g 0 n0_10366_8841  0.0483404 
iB11_210_v n1_9521_8888 0  0.0483404 
iB11_210_g 0 n0_10366_8874  0.0483404 
iB11_211_v n1_9521_9071 0  0.0483404 
iB11_211_g 0 n0_9241_9489  0.0483404 
iB11_212_v n1_9521_9104 0  0.0483404 
iB11_212_g 0 n0_9241_9489  0.0483404 
iB11_213_v n1_9521_9287 0  0.0483404 
iB11_213_g 0 n0_9241_9489  0.0483404 
iB11_214_v n1_9521_9320 0  0.0483404 
iB11_214_g 0 n0_9241_9489  0.0483404 
iB11_215_v n1_9380_9503 0  0.0483404 
iB11_215_g 0 n0_9241_9489  0.0483404 
iB11_216_v n1_9380_9536 0  0.0483404 
iB11_216_g 0 n0_9241_9522  0.0483404 
iB11_217_v n1_9521_9503 0  0.0483404 
iB11_217_g 0 n0_9241_9489  0.0483404 
iB11_218_v n1_9521_9536 0  0.0483404 
iB11_218_g 0 n0_9429_9705  0.0483404 
iB11_219_v n1_9521_9719 0  0.0483404 
iB11_219_g 0 n0_9429_9705  0.0483404 
iB11_220_v n1_9521_9752 0  0.0483404 
iB11_220_g 0 n0_9429_9738  0.0483404 
iB11_221_v n1_9521_9935 0  0.0483404 
iB11_221_g 0 n0_9429_9921  0.0483404 
iB11_222_v n1_9521_9968 0  0.0483404 
iB11_222_g 0 n0_9429_9954  0.0483404 
iB11_223_v n1_9521_10151 0  0.0483404 
iB11_223_g 0 n0_9429_10137  0.0483404 
iB11_224_v n1_9521_10184 0  0.0483404 
iB11_224_g 0 n0_9429_10170  0.0483404 
iB11_225_v n1_9521_10367 0  0.0483404 
iB11_225_g 0 n0_9429_10353  0.0483404 
iB11_226_v n1_9521_10400 0  0.0483404 
iB11_226_g 0 n0_9429_10386  0.0483404 
iB11_227_v n1_9521_10616 0  0.0483404 
iB11_227_g 0 n0_9429_10602  0.0483404 
iB30_0_v n1_16083_215 0  0.0142751 
iB30_0_g 0 n0_15146_201  0.0142751 
iB30_1_v n1_16083_248 0  0.0142751 
iB30_1_g 0 n0_15146_234  0.0142751 
iB30_2_v n1_16083_383 0  0.0142751 
iB30_2_g 0 n0_15146_417  0.0142751 
iB30_3_v n1_16083_431 0  0.0142751 
iB30_3_g 0 n0_15146_417  0.0142751 
iB30_4_v n1_16083_464 0  0.0142751 
iB30_4_g 0 n0_15146_450  0.0142751 
iB30_5_v n1_16083_647 0  0.0142751 
iB30_5_g 0 n0_15146_633  0.0142751 
iB30_6_v n1_16083_680 0  0.0142751 
iB30_6_g 0 n0_15146_666  0.0142751 
iB30_7_v n1_16130_431 0  0.0142751 
iB30_7_g 0 n0_17116_417  0.0142751 
iB30_8_v n1_16130_464 0  0.0142751 
iB30_8_g 0 n0_17116_450  0.0142751 
iB30_9_v n1_16083_863 0  0.0142751 
iB30_9_g 0 n0_15146_849  0.0142751 
iB30_10_v n1_16083_896 0  0.0142751 
iB30_10_g 0 n0_15146_882  0.0142751 
iB30_11_v n1_16083_1079 0  0.0142751 
iB30_11_g 0 n0_15146_1065  0.0142751 
iB30_12_v n1_16083_1112 0  0.0142751 
iB30_12_g 0 n0_15146_1098  0.0142751 
iB30_13_v n1_16083_1295 0  0.0142751 
iB30_13_g 0 n0_15146_1281  0.0142751 
iB30_14_v n1_16083_1328 0  0.0142751 
iB30_14_g 0 n0_15146_1314  0.0142751 
iB30_15_v n1_16083_1727 0  0.0142751 
iB30_15_g 0 n0_15146_1713  0.0142751 
iB30_16_v n1_16083_1760 0  0.0142751 
iB30_16_g 0 n0_15146_1746  0.0142751 
iB30_17_v n1_16083_1894 0  0.0142751 
iB30_17_g 0 n0_15146_1929  0.0142751 
iB30_18_v n1_16083_1943 0  0.0142751 
iB30_18_g 0 n0_15146_1929  0.0142751 
iB30_19_v n1_16083_1976 0  0.0142751 
iB30_19_g 0 n0_15146_1962  0.0142751 
iB30_20_v n1_16083_2159 0  0.0142751 
iB30_20_g 0 n0_15146_2145  0.0142751 
iB30_21_v n1_16083_2192 0  0.0142751 
iB30_21_g 0 n0_15146_2178  0.0142751 
iB30_22_v n1_16083_2375 0  0.0142751 
iB30_22_g 0 n0_15146_2361  0.0142751 
iB30_23_v n1_16083_2408 0  0.0142751 
iB30_23_g 0 n0_15146_2394  0.0142751 
iB30_24_v n1_16083_2445 0  0.0142751 
iB30_24_g 0 n0_15146_2431  0.0142751 
iB30_25_v n1_16083_2542 0  0.0142751 
iB30_25_g 0 n0_15146_2577  0.0142751 
iB30_26_v n1_16083_2543 0  0.0142751 
iB30_26_g 0 n0_15146_2577  0.0142751 
iB30_27_v n1_16083_2591 0  0.0142751 
iB30_27_g 0 n0_15146_2577  0.0142751 
iB30_28_v n1_16083_2624 0  0.0142751 
iB30_28_g 0 n0_15146_2610  0.0142751 
iB30_29_v n1_16083_2807 0  0.0142751 
iB30_29_g 0 n0_15146_2793  0.0142751 
iB30_30_v n1_16083_2840 0  0.0142751 
iB30_30_g 0 n0_15146_2826  0.0142751 
iB30_31_v n1_16083_2877 0  0.0142751 
iB30_31_g 0 n0_15146_2863  0.0142751 
iB30_32_v n1_16083_2974 0  0.0142751 
iB30_32_g 0 n0_15146_3009  0.0142751 
iB30_33_v n1_16083_3023 0  0.0142751 
iB30_33_g 0 n0_15146_3009  0.0142751 
iB30_34_v n1_16083_3056 0  0.0142751 
iB30_34_g 0 n0_15146_3042  0.0142751 
iB30_35_v n1_16083_3239 0  0.0142751 
iB30_35_g 0 n0_15146_3225  0.0142751 
iB30_36_v n1_16083_3272 0  0.0142751 
iB30_36_g 0 n0_15146_3258  0.0142751 
iB30_37_v n1_16083_3406 0  0.0142751 
iB30_37_g 0 n0_15146_3441  0.0142751 
iB30_38_v n1_16083_3455 0  0.0142751 
iB30_38_g 0 n0_15146_3441  0.0142751 
iB30_39_v n1_16083_3488 0  0.0142751 
iB30_39_g 0 n0_15146_3474  0.0142751 
iB30_40_v n1_16083_3671 0  0.0142751 
iB30_40_g 0 n0_15146_3657  0.0142751 
iB30_41_v n1_16083_3704 0  0.0142751 
iB30_41_g 0 n0_15146_3690  0.0142751 
iB30_42_v n1_16083_4103 0  0.0142751 
iB30_42_g 0 n0_15146_4089  0.0142751 
iB30_43_v n1_16083_4136 0  0.0142751 
iB30_43_g 0 n0_15146_4122  0.0142751 
iB30_44_v n1_16083_4319 0  0.0142751 
iB30_44_g 0 n0_15991_5023  0.0142751 
iB30_45_v n1_16083_4352 0  0.0142751 
iB30_45_g 0 n0_15991_5023  0.0142751 
iB30_46_v n1_16083_4486 0  0.0142751 
iB30_46_g 0 n0_15991_5023  0.0142751 
iB30_47_v n1_16083_4535 0  0.0142751 
iB30_47_g 0 n0_15991_5023  0.0142751 
iB30_48_v n1_16083_4568 0  0.0142751 
iB30_48_g 0 n0_15991_5023  0.0142751 
iB30_49_v n1_16083_4702 0  0.0142751 
iB30_49_g 0 n0_15991_5023  0.0142751 
iB30_50_v n1_16083_4751 0  0.0142751 
iB30_50_g 0 n0_15991_5023  0.0142751 
iB30_51_v n1_16083_4784 0  0.0142751 
iB30_51_g 0 n0_15991_5023  0.0142751 
iB30_52_v n1_16083_4919 0  0.0142751 
iB30_52_g 0 n0_15991_5023  0.0142751 
iB30_53_v n1_16083_4967 0  0.0142751 
iB30_53_g 0 n0_15991_5023  0.0142751 
iB30_54_v n1_16083_5000 0  0.0142751 
iB30_54_g 0 n0_15991_5023  0.0142751 
iB30_55_v n1_16083_5134 0  0.0142751 
iB30_55_g 0 n0_15991_5169  0.0142751 
iB30_56_v n1_16083_5183 0  0.0142751 
iB30_56_g 0 n0_15991_5169  0.0142751 
iB30_57_v n1_16083_5216 0  0.0142751 
iB30_57_g 0 n0_15991_5202  0.0142751 
iB30_58_v n1_16083_5253 0  0.0142751 
iB30_58_g 0 n0_15991_5239  0.0142751 
iB30_59_v n1_16130_4919 0  0.0142751 
iB30_59_g 0 n0_15991_5023  0.0142751 
iB30_60_v n1_16130_4967 0  0.0142751 
iB30_60_g 0 n0_15991_5023  0.0142751 
iB30_61_v n1_16130_5000 0  0.0142751 
iB30_61_g 0 n0_15991_5023  0.0142751 
iB30_62_v n1_16271_215 0  0.0142751 
iB30_62_g 0 n0_17116_201  0.0142751 
iB30_63_v n1_16271_248 0  0.0142751 
iB30_63_g 0 n0_17116_234  0.0142751 
iB30_64_v n1_16271_383 0  0.0142751 
iB30_64_g 0 n0_17116_417  0.0142751 
iB30_65_v n1_16364_215 0  0.0142751 
iB30_65_g 0 n0_17116_201  0.0142751 
iB30_66_v n1_16364_248 0  0.0142751 
iB30_66_g 0 n0_17116_234  0.0142751 
iB30_67_v n1_16364_383 0  0.0142751 
iB30_67_g 0 n0_17116_417  0.0142751 
iB30_68_v n1_16271_431 0  0.0142751 
iB30_68_g 0 n0_17116_417  0.0142751 
iB30_69_v n1_16271_647 0  0.0142751 
iB30_69_g 0 n0_17116_633  0.0142751 
iB30_70_v n1_16271_680 0  0.0142751 
iB30_70_g 0 n0_17116_666  0.0142751 
iB30_71_v n1_16364_431 0  0.0142751 
iB30_71_g 0 n0_17116_417  0.0142751 
iB30_72_v n1_16364_464 0  0.0142751 
iB30_72_g 0 n0_17116_450  0.0142751 
iB30_73_v n1_16364_647 0  0.0142751 
iB30_73_g 0 n0_17116_633  0.0142751 
iB30_74_v n1_16364_680 0  0.0142751 
iB30_74_g 0 n0_17116_666  0.0142751 
iB30_75_v n1_16271_863 0  0.0142751 
iB30_75_g 0 n0_17116_849  0.0142751 
iB30_76_v n1_16271_896 0  0.0142751 
iB30_76_g 0 n0_17116_882  0.0142751 
iB30_77_v n1_16271_1079 0  0.0142751 
iB30_77_g 0 n0_17116_1065  0.0142751 
iB30_78_v n1_16271_1112 0  0.0142751 
iB30_78_g 0 n0_17116_1098  0.0142751 
iB30_79_v n1_16364_863 0  0.0142751 
iB30_79_g 0 n0_17116_849  0.0142751 
iB30_80_v n1_16364_896 0  0.0142751 
iB30_80_g 0 n0_17116_882  0.0142751 
iB30_81_v n1_16364_1079 0  0.0142751 
iB30_81_g 0 n0_17116_1065  0.0142751 
iB30_82_v n1_16364_1112 0  0.0142751 
iB30_82_g 0 n0_17116_1098  0.0142751 
iB30_83_v n1_16271_1295 0  0.0142751 
iB30_83_g 0 n0_17116_1281  0.0142751 
iB30_84_v n1_16271_1328 0  0.0142751 
iB30_84_g 0 n0_17116_1314  0.0142751 
iB30_85_v n1_16271_1511 0  0.0142751 
iB30_85_g 0 n0_17116_1497  0.0142751 
iB30_86_v n1_16271_1544 0  0.0142751 
iB30_86_g 0 n0_17116_1530  0.0142751 
iB30_87_v n1_16364_1295 0  0.0142751 
iB30_87_g 0 n0_17116_1281  0.0142751 
iB30_88_v n1_16364_1328 0  0.0142751 
iB30_88_g 0 n0_17116_1314  0.0142751 
iB30_89_v n1_16364_1511 0  0.0142751 
iB30_89_g 0 n0_17116_1497  0.0142751 
iB30_90_v n1_16364_1544 0  0.0142751 
iB30_90_g 0 n0_17116_1530  0.0142751 
iB30_91_v n1_16271_1727 0  0.0142751 
iB30_91_g 0 n0_17116_1713  0.0142751 
iB30_92_v n1_16271_1760 0  0.0142751 
iB30_92_g 0 n0_17116_1746  0.0142751 
iB30_93_v n1_16271_1894 0  0.0142751 
iB30_93_g 0 n0_17116_1929  0.0142751 
iB30_94_v n1_16271_1943 0  0.0142751 
iB30_94_g 0 n0_17116_1929  0.0142751 
iB30_95_v n1_16271_1976 0  0.0142751 
iB30_95_g 0 n0_17116_1962  0.0142751 
iB30_96_v n1_16364_1727 0  0.0142751 
iB30_96_g 0 n0_17116_1713  0.0142751 
iB30_97_v n1_16364_1760 0  0.0142751 
iB30_97_g 0 n0_17116_1746  0.0142751 
iB30_98_v n1_16364_1894 0  0.0142751 
iB30_98_g 0 n0_17116_1929  0.0142751 
iB30_99_v n1_16364_1943 0  0.0142751 
iB30_99_g 0 n0_17116_1929  0.0142751 
iB30_100_v n1_16364_1976 0  0.0142751 
iB30_100_g 0 n0_17116_1962  0.0142751 
iB30_101_v n1_16271_2159 0  0.0142751 
iB30_101_g 0 n0_17116_2145  0.0142751 
iB30_102_v n1_16271_2192 0  0.0142751 
iB30_102_g 0 n0_17116_2178  0.0142751 
iB30_103_v n1_16271_2375 0  0.0142751 
iB30_103_g 0 n0_17116_2361  0.0142751 
iB30_104_v n1_16271_2408 0  0.0142751 
iB30_104_g 0 n0_17116_2394  0.0142751 
iB30_105_v n1_16271_2445 0  0.0142751 
iB30_105_g 0 n0_17116_2431  0.0142751 
iB30_106_v n1_16364_2159 0  0.0142751 
iB30_106_g 0 n0_17116_2145  0.0142751 
iB30_107_v n1_16364_2192 0  0.0142751 
iB30_107_g 0 n0_17116_2178  0.0142751 
iB30_108_v n1_16364_2375 0  0.0142751 
iB30_108_g 0 n0_17116_2361  0.0142751 
iB30_109_v n1_16364_2408 0  0.0142751 
iB30_109_g 0 n0_17116_2394  0.0142751 
iB30_110_v n1_16364_2445 0  0.0142751 
iB30_110_g 0 n0_17116_2431  0.0142751 
iB30_111_v n1_16271_2542 0  0.0142751 
iB30_111_g 0 n0_17116_2577  0.0142751 
iB30_112_v n1_16271_2543 0  0.0142751 
iB30_112_g 0 n0_17116_2577  0.0142751 
iB30_113_v n1_16271_2591 0  0.0142751 
iB30_113_g 0 n0_17116_2577  0.0142751 
iB30_114_v n1_16271_2624 0  0.0142751 
iB30_114_g 0 n0_17116_2610  0.0142751 
iB30_115_v n1_16271_2807 0  0.0142751 
iB30_115_g 0 n0_17116_2793  0.0142751 
iB30_116_v n1_16271_2840 0  0.0142751 
iB30_116_g 0 n0_17116_2826  0.0142751 
iB30_117_v n1_16364_2542 0  0.0142751 
iB30_117_g 0 n0_17116_2577  0.0142751 
iB30_118_v n1_16364_2543 0  0.0142751 
iB30_118_g 0 n0_17116_2577  0.0142751 
iB30_119_v n1_16364_2591 0  0.0142751 
iB30_119_g 0 n0_17116_2577  0.0142751 
iB30_120_v n1_16364_2624 0  0.0142751 
iB30_120_g 0 n0_17116_2610  0.0142751 
iB30_121_v n1_16271_2877 0  0.0142751 
iB30_121_g 0 n0_17116_2863  0.0142751 
iB30_122_v n1_16271_2974 0  0.0142751 
iB30_122_g 0 n0_17116_3009  0.0142751 
iB30_123_v n1_16271_3023 0  0.0142751 
iB30_123_g 0 n0_17116_3009  0.0142751 
iB30_124_v n1_16271_3056 0  0.0142751 
iB30_124_g 0 n0_17116_3042  0.0142751 
iB30_125_v n1_16271_3239 0  0.0142751 
iB30_125_g 0 n0_17116_3225  0.0142751 
iB30_126_v n1_16271_3272 0  0.0142751 
iB30_126_g 0 n0_17116_3258  0.0142751 
iB30_127_v n1_16271_3406 0  0.0142751 
iB30_127_g 0 n0_17116_3441  0.0142751 
iB30_128_v n1_16271_3455 0  0.0142751 
iB30_128_g 0 n0_17116_3441  0.0142751 
iB30_129_v n1_16271_3488 0  0.0142751 
iB30_129_g 0 n0_17116_3474  0.0142751 
iB30_130_v n1_16271_3671 0  0.0142751 
iB30_130_g 0 n0_17116_3657  0.0142751 
iB30_131_v n1_16271_3704 0  0.0142751 
iB30_131_g 0 n0_17116_3690  0.0142751 
iB30_132_v n1_16271_3887 0  0.0142751 
iB30_132_g 0 n0_17116_3873  0.0142751 
iB30_133_v n1_16271_3920 0  0.0142751 
iB30_133_g 0 n0_17116_3906  0.0142751 
iB30_134_v n1_16271_4103 0  0.0142751 
iB30_134_g 0 n0_17116_4089  0.0142751 
iB30_135_v n1_16271_4136 0  0.0142751 
iB30_135_g 0 n0_17116_4122  0.0142751 
iB30_136_v n1_16271_4319 0  0.0142751 
iB30_136_g 0 n0_15991_5023  0.0142751 
iB30_137_v n1_16271_4352 0  0.0142751 
iB30_137_g 0 n0_15991_5023  0.0142751 
iB30_138_v n1_16271_4486 0  0.0142751 
iB30_138_g 0 n0_15991_5023  0.0142751 
iB30_139_v n1_16271_4535 0  0.0142751 
iB30_139_g 0 n0_15991_5023  0.0142751 
iB30_140_v n1_16271_4568 0  0.0142751 
iB30_140_g 0 n0_15991_5023  0.0142751 
iB30_141_v n1_16271_4702 0  0.0142751 
iB30_141_g 0 n0_15991_5023  0.0142751 
iB30_142_v n1_16271_4751 0  0.0142751 
iB30_142_g 0 n0_15991_5023  0.0142751 
iB30_143_v n1_16271_4784 0  0.0142751 
iB30_143_g 0 n0_15991_5023  0.0142751 
iB30_144_v n1_16271_4919 0  0.0142751 
iB30_144_g 0 n0_16179_5169  0.0142751 
iB30_145_v n1_16271_5000 0  0.0142751 
iB30_145_g 0 n0_16179_5169  0.0142751 
iB30_146_v n1_16271_5134 0  0.0142751 
iB30_146_g 0 n0_16179_5169  0.0142751 
iB30_147_v n1_16271_5183 0  0.0142751 
iB30_147_g 0 n0_16179_5169  0.0142751 
iB30_148_v n1_16271_5216 0  0.0142751 
iB30_148_g 0 n0_16179_5202  0.0142751 
iB30_149_v n1_16271_5253 0  0.0142751 
iB30_149_g 0 n0_16179_5239  0.0142751 
iB30_150_v n1_18150_215 0  0.0142751 
iB30_150_g 0 n0_17396_201  0.0142751 
iB30_151_v n1_18150_248 0  0.0142751 
iB30_151_g 0 n0_17396_234  0.0142751 
iB30_152_v n1_18150_383 0  0.0142751 
iB30_152_g 0 n0_17396_417  0.0142751 
iB30_153_v n1_18150_431 0  0.0142751 
iB30_153_g 0 n0_17396_417  0.0142751 
iB30_154_v n1_18150_464 0  0.0142751 
iB30_154_g 0 n0_17396_450  0.0142751 
iB30_155_v n1_18150_647 0  0.0142751 
iB30_155_g 0 n0_17396_633  0.0142751 
iB30_156_v n1_18150_680 0  0.0142751 
iB30_156_g 0 n0_17396_666  0.0142751 
iB30_157_v n1_18150_863 0  0.0142751 
iB30_157_g 0 n0_17396_849  0.0142751 
iB30_158_v n1_18150_896 0  0.0142751 
iB30_158_g 0 n0_17396_882  0.0142751 
iB30_159_v n1_18150_1079 0  0.0142751 
iB30_159_g 0 n0_17396_1065  0.0142751 
iB30_160_v n1_18150_1112 0  0.0142751 
iB30_160_g 0 n0_17396_1098  0.0142751 
iB30_161_v n1_18150_1295 0  0.0142751 
iB30_161_g 0 n0_17396_1281  0.0142751 
iB30_162_v n1_18150_1328 0  0.0142751 
iB30_162_g 0 n0_17396_1314  0.0142751 
iB30_163_v n1_18150_1511 0  0.0142751 
iB30_163_g 0 n0_17396_1497  0.0142751 
iB30_164_v n1_18150_1544 0  0.0142751 
iB30_164_g 0 n0_17396_1530  0.0142751 
iB30_165_v n1_18150_1727 0  0.0142751 
iB30_165_g 0 n0_17396_1713  0.0142751 
iB30_166_v n1_18150_1760 0  0.0142751 
iB30_166_g 0 n0_17396_1746  0.0142751 
iB30_167_v n1_18150_1894 0  0.0142751 
iB30_167_g 0 n0_17396_1929  0.0142751 
iB30_168_v n1_18150_1943 0  0.0142751 
iB30_168_g 0 n0_17396_1929  0.0142751 
iB30_169_v n1_18150_1976 0  0.0142751 
iB30_169_g 0 n0_17396_1962  0.0142751 
iB30_170_v n1_18150_2159 0  0.0142751 
iB30_170_g 0 n0_18241_2793  0.0142751 
iB30_171_v n1_18150_2192 0  0.0142751 
iB30_171_g 0 n0_18241_2793  0.0142751 
iB30_172_v n1_18150_2375 0  0.0142751 
iB30_172_g 0 n0_18241_2793  0.0142751 
iB30_173_v n1_18150_2408 0  0.0142751 
iB30_173_g 0 n0_18241_2793  0.0142751 
iB30_174_v n1_18150_2542 0  0.0142751 
iB30_174_g 0 n0_18241_2793  0.0142751 
iB30_175_v n1_18150_2543 0  0.0142751 
iB30_175_g 0 n0_18241_2793  0.0142751 
iB30_176_v n1_18150_2591 0  0.0142751 
iB30_176_g 0 n0_18241_2793  0.0142751 
iB30_177_v n1_18150_2624 0  0.0142751 
iB30_177_g 0 n0_18241_2793  0.0142751 
iB30_178_v n1_18333_215 0  0.0142751 
iB30_178_g 0 n0_17396_201  0.0142751 
iB30_179_v n1_18333_248 0  0.0142751 
iB30_179_g 0 n0_17396_234  0.0142751 
iB30_180_v n1_18333_383 0  0.0142751 
iB30_180_g 0 n0_17396_417  0.0142751 
iB30_181_v n1_18521_215 0  0.0142751 
iB30_181_g 0 n0_19366_201  0.0142751 
iB30_182_v n1_18521_248 0  0.0142751 
iB30_182_g 0 n0_19366_234  0.0142751 
iB30_183_v n1_18521_383 0  0.0142751 
iB30_183_g 0 n0_19366_417  0.0142751 
iB30_184_v n1_18333_431 0  0.0142751 
iB30_184_g 0 n0_17396_417  0.0142751 
iB30_185_v n1_18333_464 0  0.0142751 
iB30_185_g 0 n0_17396_450  0.0142751 
iB30_186_v n1_18333_647 0  0.0142751 
iB30_186_g 0 n0_17396_633  0.0142751 
iB30_187_v n1_18333_680 0  0.0142751 
iB30_187_g 0 n0_17396_666  0.0142751 
iB30_188_v n1_18380_431 0  0.0142751 
iB30_188_g 0 n0_17396_417  0.0142751 
iB30_189_v n1_18380_464 0  0.0142751 
iB30_189_g 0 n0_17396_450  0.0142751 
iB30_190_v n1_18521_431 0  0.0142751 
iB30_190_g 0 n0_19366_417  0.0142751 
iB30_191_v n1_18521_647 0  0.0142751 
iB30_191_g 0 n0_19366_633  0.0142751 
iB30_192_v n1_18521_680 0  0.0142751 
iB30_192_g 0 n0_19366_666  0.0142751 
iB30_193_v n1_18333_863 0  0.0142751 
iB30_193_g 0 n0_17396_849  0.0142751 
iB30_194_v n1_18333_896 0  0.0142751 
iB30_194_g 0 n0_17396_882  0.0142751 
iB30_195_v n1_18333_1079 0  0.0142751 
iB30_195_g 0 n0_17396_1065  0.0142751 
iB30_196_v n1_18333_1112 0  0.0142751 
iB30_196_g 0 n0_17396_1098  0.0142751 
iB30_197_v n1_18521_863 0  0.0142751 
iB30_197_g 0 n0_19366_849  0.0142751 
iB30_198_v n1_18521_896 0  0.0142751 
iB30_198_g 0 n0_19366_882  0.0142751 
iB30_199_v n1_18521_1079 0  0.0142751 
iB30_199_g 0 n0_19366_1065  0.0142751 
iB30_200_v n1_18521_1112 0  0.0142751 
iB30_200_g 0 n0_19366_1098  0.0142751 
iB30_201_v n1_18333_1295 0  0.0142751 
iB30_201_g 0 n0_17396_1281  0.0142751 
iB30_202_v n1_18333_1328 0  0.0142751 
iB30_202_g 0 n0_17396_1314  0.0142751 
iB30_203_v n1_18521_1295 0  0.0142751 
iB30_203_g 0 n0_19366_1281  0.0142751 
iB30_204_v n1_18521_1328 0  0.0142751 
iB30_204_g 0 n0_19366_1314  0.0142751 
iB30_205_v n1_18521_1511 0  0.0142751 
iB30_205_g 0 n0_19366_1497  0.0142751 
iB30_206_v n1_18521_1544 0  0.0142751 
iB30_206_g 0 n0_19366_1530  0.0142751 
iB30_207_v n1_18333_1727 0  0.0142751 
iB30_207_g 0 n0_17396_1713  0.0142751 
iB30_208_v n1_18333_1760 0  0.0142751 
iB30_208_g 0 n0_17396_1746  0.0142751 
iB30_209_v n1_18333_1894 0  0.0142751 
iB30_209_g 0 n0_17396_1929  0.0142751 
iB30_210_v n1_18333_1943 0  0.0142751 
iB30_210_g 0 n0_18241_2793  0.0142751 
iB30_211_v n1_18333_1976 0  0.0142751 
iB30_211_g 0 n0_18241_2793  0.0142751 
iB30_212_v n1_18521_1727 0  0.0142751 
iB30_212_g 0 n0_19366_1713  0.0142751 
iB30_213_v n1_18521_1760 0  0.0142751 
iB30_213_g 0 n0_19366_1746  0.0142751 
iB30_214_v n1_18521_1894 0  0.0142751 
iB30_214_g 0 n0_19366_1929  0.0142751 
iB30_215_v n1_18521_1943 0  0.0142751 
iB30_215_g 0 n0_19366_1929  0.0142751 
iB30_216_v n1_18521_1976 0  0.0142751 
iB30_216_g 0 n0_18429_2826  0.0142751 
iB30_217_v n1_18333_2110 0  0.0142751 
iB30_217_g 0 n0_18241_2793  0.0142751 
iB30_218_v n1_18333_2159 0  0.0142751 
iB30_218_g 0 n0_18241_2793  0.0142751 
iB30_219_v n1_18333_2192 0  0.0142751 
iB30_219_g 0 n0_18241_2793  0.0142751 
iB30_220_v n1_18333_2375 0  0.0142751 
iB30_220_g 0 n0_18241_2793  0.0142751 
iB30_221_v n1_18333_2408 0  0.0142751 
iB30_221_g 0 n0_18241_2793  0.0142751 
iB30_222_v n1_18521_2110 0  0.0142751 
iB30_222_g 0 n0_18429_2826  0.0142751 
iB30_223_v n1_18521_2159 0  0.0142751 
iB30_223_g 0 n0_18429_2826  0.0142751 
iB30_224_v n1_18521_2192 0  0.0142751 
iB30_224_g 0 n0_18429_2826  0.0142751 
iB30_225_v n1_18521_2375 0  0.0142751 
iB30_225_g 0 n0_18429_2826  0.0142751 
iB30_226_v n1_18521_2408 0  0.0142751 
iB30_226_g 0 n0_18429_2826  0.0142751 
iB30_227_v n1_18333_2542 0  0.0142751 
iB30_227_g 0 n0_18241_2793  0.0142751 
iB30_228_v n1_18333_2543 0  0.0142751 
iB30_228_g 0 n0_18241_2793  0.0142751 
iB30_229_v n1_18333_2591 0  0.0142751 
iB30_229_g 0 n0_18241_2793  0.0142751 
iB30_230_v n1_18333_2624 0  0.0142751 
iB30_230_g 0 n0_18241_2793  0.0142751 
iB30_231_v n1_18333_2807 0  0.0142751 
iB30_231_g 0 n0_18241_2793  0.0142751 
iB30_232_v n1_18333_2840 0  0.0142751 
iB30_232_g 0 n0_18241_2826  0.0142751 
iB30_233_v n1_18521_2542 0  0.0142751 
iB30_233_g 0 n0_18429_2826  0.0142751 
iB30_234_v n1_18521_2543 0  0.0142751 
iB30_234_g 0 n0_18429_2826  0.0142751 
iB30_235_v n1_18521_2591 0  0.0142751 
iB30_235_g 0 n0_18429_2826  0.0142751 
iB30_236_v n1_18521_2624 0  0.0142751 
iB30_236_g 0 n0_18429_2826  0.0142751 
iB30_237_v n1_18521_2807 0  0.0142751 
iB30_237_g 0 n0_18429_2826  0.0142751 
iB30_238_v n1_18521_2840 0  0.0142751 
iB30_238_g 0 n0_18429_2826  0.0142751 
iB30_239_v n1_18333_3023 0  0.0142751 
iB30_239_g 0 n0_18241_3009  0.0142751 
iB30_240_v n1_18333_3056 0  0.0142751 
iB30_240_g 0 n0_18241_3042  0.0142751 
iB30_241_v n1_18333_3239 0  0.0142751 
iB30_241_g 0 n0_18241_3225  0.0142751 
iB30_242_v n1_18521_3023 0  0.0142751 
iB30_242_g 0 n0_18429_3009  0.0142751 
iB30_243_v n1_18521_3056 0  0.0142751 
iB30_243_g 0 n0_18429_3042  0.0142751 
iB30_244_v n1_18521_3239 0  0.0142751 
iB30_244_g 0 n0_18429_3225  0.0142751 
iB30_245_v n1_18333_3272 0  0.0142751 
iB30_245_g 0 n0_18241_3258  0.0142751 
iB30_246_v n1_18333_3406 0  0.0142751 
iB30_246_g 0 n0_18241_3441  0.0142751 
iB30_247_v n1_18333_3455 0  0.0142751 
iB30_247_g 0 n0_18241_3441  0.0142751 
iB30_248_v n1_18333_3488 0  0.0142751 
iB30_248_g 0 n0_18241_3474  0.0142751 
iB30_249_v n1_18333_3671 0  0.0142751 
iB30_249_g 0 n0_18241_3657  0.0142751 
iB30_250_v n1_18521_3272 0  0.0142751 
iB30_250_g 0 n0_18429_3258  0.0142751 
iB30_251_v n1_18521_3406 0  0.0142751 
iB30_251_g 0 n0_18429_3441  0.0142751 
iB30_252_v n1_18521_3455 0  0.0142751 
iB30_252_g 0 n0_18429_3441  0.0142751 
iB30_253_v n1_18521_3488 0  0.0142751 
iB30_253_g 0 n0_18429_3474  0.0142751 
iB30_254_v n1_18521_3671 0  0.0142751 
iB30_254_g 0 n0_18429_3657  0.0142751 
iB30_255_v n1_18333_3704 0  0.0142751 
iB30_255_g 0 n0_18241_3690  0.0142751 
iB30_256_v n1_18521_3704 0  0.0142751 
iB30_256_g 0 n0_18429_3690  0.0142751 
iB30_257_v n1_18521_3887 0  0.0142751 
iB30_257_g 0 n0_18429_3873  0.0142751 
iB30_258_v n1_18521_3920 0  0.0142751 
iB30_258_g 0 n0_18429_3906  0.0142751 
iB30_259_v n1_18333_4103 0  0.0142751 
iB30_259_g 0 n0_18241_4089  0.0142751 
iB30_260_v n1_18333_4136 0  0.0142751 
iB30_260_g 0 n0_18241_4122  0.0142751 
iB30_261_v n1_18333_4319 0  0.0142751 
iB30_261_g 0 n0_18241_4305  0.0142751 
iB30_262_v n1_18333_4352 0  0.0142751 
iB30_262_g 0 n0_18241_4338  0.0142751 
iB30_263_v n1_18333_4486 0  0.0142751 
iB30_263_g 0 n0_18241_4521  0.0142751 
iB30_264_v n1_18521_4103 0  0.0142751 
iB30_264_g 0 n0_18429_4089  0.0142751 
iB30_265_v n1_18521_4136 0  0.0142751 
iB30_265_g 0 n0_18429_4122  0.0142751 
iB30_266_v n1_18521_4319 0  0.0142751 
iB30_266_g 0 n0_18429_4305  0.0142751 
iB30_267_v n1_18521_4352 0  0.0142751 
iB30_267_g 0 n0_18429_4338  0.0142751 
iB30_268_v n1_18521_4486 0  0.0142751 
iB30_268_g 0 n0_18429_4521  0.0142751 
iB30_269_v n1_18333_4535 0  0.0142751 
iB30_269_g 0 n0_18241_4521  0.0142751 
iB30_270_v n1_18333_4568 0  0.0142751 
iB30_270_g 0 n0_18241_4554  0.0142751 
iB30_271_v n1_18333_4702 0  0.0142751 
iB30_271_g 0 n0_18241_4737  0.0142751 
iB30_272_v n1_18333_4751 0  0.0142751 
iB30_272_g 0 n0_18241_4737  0.0142751 
iB30_273_v n1_18333_4784 0  0.0142751 
iB30_273_g 0 n0_18241_4770  0.0142751 
iB30_274_v n1_18521_4535 0  0.0142751 
iB30_274_g 0 n0_18429_4521  0.0142751 
iB30_275_v n1_18521_4568 0  0.0142751 
iB30_275_g 0 n0_18429_4554  0.0142751 
iB30_276_v n1_18521_4702 0  0.0142751 
iB30_276_g 0 n0_18429_4737  0.0142751 
iB30_277_v n1_18521_4751 0  0.0142751 
iB30_277_g 0 n0_18429_4737  0.0142751 
iB30_278_v n1_18521_4784 0  0.0142751 
iB30_278_g 0 n0_18429_4770  0.0142751 
iB30_279_v n1_18333_4920 0  0.0142751 
iB30_279_g 0 n0_18241_4953  0.0142751 
iB30_280_v n1_18333_4967 0  0.0142751 
iB30_280_g 0 n0_18241_4953  0.0142751 
iB30_281_v n1_18333_5000 0  0.0142751 
iB30_281_g 0 n0_18241_4986  0.0142751 
iB30_282_v n1_18333_5134 0  0.0142751 
iB30_282_g 0 n0_18241_5169  0.0142751 
iB30_283_v n1_18333_5183 0  0.0142751 
iB30_283_g 0 n0_18241_5169  0.0142751 
iB30_284_v n1_18333_5216 0  0.0142751 
iB30_284_g 0 n0_18241_5202  0.0142751 
iB30_285_v n1_18333_5253 0  0.0142751 
iB30_285_g 0 n0_18241_5239  0.0142751 
iB30_286_v n1_18380_4920 0  0.0142751 
iB30_286_g 0 n0_18429_4807  0.0142751 
iB30_287_v n1_18380_4967 0  0.0142751 
iB30_287_g 0 n0_18241_4953  0.0142751 
iB30_288_v n1_18380_5000 0  0.0142751 
iB30_288_g 0 n0_18241_4986  0.0142751 
iB30_289_v n1_18521_4920 0  0.0142751 
iB30_289_g 0 n0_18429_4807  0.0142751 
iB30_290_v n1_18521_5000 0  0.0142751 
iB30_290_g 0 n0_18429_5169  0.0142751 
iB30_291_v n1_18521_5134 0  0.0142751 
iB30_291_g 0 n0_18429_5169  0.0142751 
iB30_292_v n1_18521_5183 0  0.0142751 
iB30_292_g 0 n0_18429_5169  0.0142751 
iB30_293_v n1_18521_5216 0  0.0142751 
iB30_293_g 0 n0_18429_5202  0.0142751 
iB30_294_v n1_18521_5253 0  0.0142751 
iB30_294_g 0 n0_18429_5239  0.0142751 
iB30_295_v n1_18614_215 0  0.0142751 
iB30_295_g 0 n0_19366_201  0.0142751 
iB30_296_v n1_18614_248 0  0.0142751 
iB30_296_g 0 n0_19366_234  0.0142751 
iB30_297_v n1_18614_383 0  0.0142751 
iB30_297_g 0 n0_19366_417  0.0142751 
iB30_298_v n1_18614_431 0  0.0142751 
iB30_298_g 0 n0_19366_417  0.0142751 
iB30_299_v n1_18614_464 0  0.0142751 
iB30_299_g 0 n0_19366_450  0.0142751 
iB30_300_v n1_18614_647 0  0.0142751 
iB30_300_g 0 n0_19366_633  0.0142751 
iB30_301_v n1_18614_680 0  0.0142751 
iB30_301_g 0 n0_19366_666  0.0142751 
iB30_302_v n1_18614_863 0  0.0142751 
iB30_302_g 0 n0_19366_849  0.0142751 
iB30_303_v n1_18614_896 0  0.0142751 
iB30_303_g 0 n0_19366_882  0.0142751 
iB30_304_v n1_18614_1079 0  0.0142751 
iB30_304_g 0 n0_19366_1065  0.0142751 
iB30_305_v n1_18614_1112 0  0.0142751 
iB30_305_g 0 n0_19366_1098  0.0142751 
iB30_306_v n1_18614_1295 0  0.0142751 
iB30_306_g 0 n0_19366_1281  0.0142751 
iB30_307_v n1_18614_1328 0  0.0142751 
iB30_307_g 0 n0_19366_1314  0.0142751 
iB30_308_v n1_18614_1511 0  0.0142751 
iB30_308_g 0 n0_19366_1497  0.0142751 
iB30_309_v n1_18614_1544 0  0.0142751 
iB30_309_g 0 n0_19366_1530  0.0142751 
iB30_310_v n1_18614_1727 0  0.0142751 
iB30_310_g 0 n0_19366_1713  0.0142751 
iB30_311_v n1_18614_1760 0  0.0142751 
iB30_311_g 0 n0_19366_1746  0.0142751 
iB30_312_v n1_18614_1943 0  0.0142751 
iB30_312_g 0 n0_19366_1929  0.0142751 
iB30_313_v n1_18614_1976 0  0.0142751 
iB30_313_g 0 n0_18429_2826  0.0142751 
iB30_314_v n1_18614_2110 0  0.0142751 
iB30_314_g 0 n0_18429_2826  0.0142751 
iB30_315_v n1_18614_2159 0  0.0142751 
iB30_315_g 0 n0_18429_2826  0.0142751 
iB30_316_v n1_18614_2192 0  0.0142751 
iB30_316_g 0 n0_18429_2826  0.0142751 
iB30_317_v n1_18614_2375 0  0.0142751 
iB30_317_g 0 n0_18429_2826  0.0142751 
iB30_318_v n1_18614_2408 0  0.0142751 
iB30_318_g 0 n0_18429_2826  0.0142751 
iB30_319_v n1_18614_2543 0  0.0142751 
iB30_319_g 0 n0_18429_2826  0.0142751 
iB30_320_v n1_18614_2591 0  0.0142751 
iB30_320_g 0 n0_18429_2826  0.0142751 
iB30_321_v n1_18614_2624 0  0.0142751 
iB30_321_g 0 n0_18429_2826  0.0142751 
iB30_322_v n1_20583_215 0  0.0142751 
iB30_322_g 0 n0_20491_633  0.0142751 
iB30_323_v n1_20583_248 0  0.0142751 
iB30_323_g 0 n0_20491_633  0.0142751 
iB30_324_v n1_20583_383 0  0.0142751 
iB30_324_g 0 n0_20491_633  0.0142751 
iB30_325_v n1_20583_431 0  0.0142751 
iB30_325_g 0 n0_20491_633  0.0142751 
iB30_326_v n1_20583_464 0  0.0142751 
iB30_326_g 0 n0_20491_633  0.0142751 
iB30_327_v n1_20583_647 0  0.0142751 
iB30_327_g 0 n0_20491_633  0.0142751 
iB30_328_v n1_20583_680 0  0.0142751 
iB30_328_g 0 n0_20491_666  0.0142751 
iB30_329_v n1_20630_431 0  0.0142751 
iB30_329_g 0 n0_20679_633  0.0142751 
iB30_330_v n1_20630_464 0  0.0142751 
iB30_330_g 0 n0_20679_633  0.0142751 
iB30_331_v n1_20771_647 0  0.0142751 
iB30_331_g 0 n0_20679_633  0.0142751 
iB30_332_v n1_20771_680 0  0.0142751 
iB30_332_g 0 n0_20679_666  0.0142751 
iB30_333_v n1_20583_863 0  0.0142751 
iB30_333_g 0 n0_20491_849  0.0142751 
iB30_334_v n1_20583_896 0  0.0142751 
iB30_334_g 0 n0_20491_882  0.0142751 
iB30_335_v n1_20583_1079 0  0.0142751 
iB30_335_g 0 n0_20491_1065  0.0142751 
iB30_336_v n1_20583_1112 0  0.0142751 
iB30_336_g 0 n0_20491_1098  0.0142751 
iB30_337_v n1_20771_863 0  0.0142751 
iB30_337_g 0 n0_20679_849  0.0142751 
iB30_338_v n1_20771_896 0  0.0142751 
iB30_338_g 0 n0_20679_882  0.0142751 
iB30_339_v n1_20771_1079 0  0.0142751 
iB30_339_g 0 n0_20679_1065  0.0142751 
iB30_340_v n1_20771_1112 0  0.0142751 
iB30_340_g 0 n0_20679_1098  0.0142751 
iB30_341_v n1_20583_1295 0  0.0142751 
iB30_341_g 0 n0_20491_1281  0.0142751 
iB30_342_v n1_20583_1328 0  0.0142751 
iB30_342_g 0 n0_20491_1314  0.0142751 
iB30_343_v n1_20771_1295 0  0.0142751 
iB30_343_g 0 n0_20679_1281  0.0142751 
iB30_344_v n1_20771_1328 0  0.0142751 
iB30_344_g 0 n0_20679_1314  0.0142751 
iB30_345_v n1_20771_1511 0  0.0142751 
iB30_345_g 0 n0_20679_1497  0.0142751 
iB30_346_v n1_20771_1544 0  0.0142751 
iB30_346_g 0 n0_20679_1530  0.0142751 
iB30_347_v n1_20583_1727 0  0.0142751 
iB30_347_g 0 n0_20491_1713  0.0142751 
iB30_348_v n1_20583_1760 0  0.0142751 
iB30_348_g 0 n0_20491_1746  0.0142751 
iB30_349_v n1_20583_1943 0  0.0142751 
iB30_349_g 0 n0_20491_1929  0.0142751 
iB30_350_v n1_20583_1976 0  0.0142751 
iB30_350_g 0 n0_20491_1976  0.0142751 
iB30_351_v n1_20771_1727 0  0.0142751 
iB30_351_g 0 n0_20679_1713  0.0142751 
iB30_352_v n1_20771_1760 0  0.0142751 
iB30_352_g 0 n0_20679_1746  0.0142751 
iB30_353_v n1_20771_1943 0  0.0142751 
iB30_353_g 0 n0_20679_1929  0.0142751 
iB30_354_v n1_20771_1976 0  0.0142751 
iB30_354_g 0 n0_20679_1976  0.0142751 
iB30_355_v n1_20583_2159 0  0.0142751 
iB30_355_g 0 n0_20491_2145  0.0142751 
iB30_356_v n1_20583_2192 0  0.0142751 
iB30_356_g 0 n0_20491_2178  0.0142751 
iB30_357_v n1_20583_2375 0  0.0142751 
iB30_357_g 0 n0_20491_2361  0.0142751 
iB30_358_v n1_20583_2408 0  0.0142751 
iB30_358_g 0 n0_20491_2394  0.0142751 
iB30_359_v n1_20771_2159 0  0.0142751 
iB30_359_g 0 n0_20679_2145  0.0142751 
iB30_360_v n1_20771_2192 0  0.0142751 
iB30_360_g 0 n0_20679_2178  0.0142751 
iB30_361_v n1_20771_2375 0  0.0142751 
iB30_361_g 0 n0_20679_2361  0.0142751 
iB30_362_v n1_20771_2408 0  0.0142751 
iB30_362_g 0 n0_20679_2394  0.0142751 
iB30_363_v n1_20583_2543 0  0.0142751 
iB30_363_g 0 n0_20491_2577  0.0142751 
iB30_364_v n1_20583_2591 0  0.0142751 
iB30_364_g 0 n0_20491_2577  0.0142751 
iB30_365_v n1_20583_2624 0  0.0142751 
iB30_365_g 0 n0_20491_2610  0.0142751 
iB30_366_v n1_20583_2807 0  0.0142751 
iB30_366_g 0 n0_20491_2793  0.0142751 
iB30_367_v n1_20583_2840 0  0.0142751 
iB30_367_g 0 n0_20491_2826  0.0142751 
iB30_368_v n1_20771_2543 0  0.0142751 
iB30_368_g 0 n0_20679_2577  0.0142751 
iB30_369_v n1_20771_2591 0  0.0142751 
iB30_369_g 0 n0_20679_2577  0.0142751 
iB30_370_v n1_20771_2624 0  0.0142751 
iB30_370_g 0 n0_20679_2610  0.0142751 
iB30_371_v n1_20771_2807 0  0.0142751 
iB30_371_g 0 n0_20679_2826  0.0142751 
iB30_372_v n1_20771_2840 0  0.0142751 
iB30_372_g 0 n0_20679_2826  0.0142751 
iB30_373_v n1_20583_3023 0  0.0142751 
iB30_373_g 0 n0_20491_3009  0.0142751 
iB30_374_v n1_20583_3056 0  0.0142751 
iB30_374_g 0 n0_20491_3042  0.0142751 
iB30_375_v n1_20583_3239 0  0.0142751 
iB30_375_g 0 n0_20491_3225  0.0142751 
iB30_376_v n1_20771_3023 0  0.0142751 
iB30_376_g 0 n0_20679_3009  0.0142751 
iB30_377_v n1_20771_3056 0  0.0142751 
iB30_377_g 0 n0_20679_3042  0.0142751 
iB30_378_v n1_20771_3239 0  0.0142751 
iB30_378_g 0 n0_20679_3225  0.0142751 
iB30_379_v n1_20583_3272 0  0.0142751 
iB30_379_g 0 n0_20491_3258  0.0142751 
iB30_380_v n1_20583_3455 0  0.0142751 
iB30_380_g 0 n0_20491_3441  0.0142751 
iB30_381_v n1_20583_3488 0  0.0142751 
iB30_381_g 0 n0_20491_3474  0.0142751 
iB30_382_v n1_20583_3671 0  0.0142751 
iB30_382_g 0 n0_20491_3657  0.0142751 
iB30_383_v n1_20771_3272 0  0.0142751 
iB30_383_g 0 n0_20679_3258  0.0142751 
iB30_384_v n1_20771_3455 0  0.0142751 
iB30_384_g 0 n0_20679_3441  0.0142751 
iB30_385_v n1_20771_3488 0  0.0142751 
iB30_385_g 0 n0_20679_3474  0.0142751 
iB30_386_v n1_20771_3671 0  0.0142751 
iB30_386_g 0 n0_20679_3657  0.0142751 
iB30_387_v n1_20583_3704 0  0.0142751 
iB30_387_g 0 n0_20491_3690  0.0142751 
iB30_388_v n1_20771_3704 0  0.0142751 
iB30_388_g 0 n0_20679_3690  0.0142751 
iB30_389_v n1_20771_3887 0  0.0142751 
iB30_389_g 0 n0_20679_3873  0.0142751 
iB30_390_v n1_20771_3920 0  0.0142751 
iB30_390_g 0 n0_20679_3906  0.0142751 
iB30_391_v n1_20583_4103 0  0.0142751 
iB30_391_g 0 n0_20491_4089  0.0142751 
iB30_392_v n1_20583_4136 0  0.0142751 
iB30_392_g 0 n0_20491_4122  0.0142751 
iB30_393_v n1_20583_4319 0  0.0142751 
iB30_393_g 0 n0_20491_4305  0.0142751 
iB30_394_v n1_20583_4352 0  0.0142751 
iB30_394_g 0 n0_20491_4338  0.0142751 
iB30_395_v n1_20771_4103 0  0.0142751 
iB30_395_g 0 n0_20679_4089  0.0142751 
iB30_396_v n1_20771_4136 0  0.0142751 
iB30_396_g 0 n0_20679_4122  0.0142751 
iB30_397_v n1_20771_4319 0  0.0142751 
iB30_397_g 0 n0_20679_4305  0.0142751 
iB30_398_v n1_20771_4352 0  0.0142751 
iB30_398_g 0 n0_20679_4338  0.0142751 
iB30_399_v n1_20583_4535 0  0.0142751 
iB30_399_g 0 n0_20491_4521  0.0142751 
iB30_400_v n1_20583_4568 0  0.0142751 
iB30_400_g 0 n0_20491_4554  0.0142751 
iB30_401_v n1_20583_4751 0  0.0142751 
iB30_401_g 0 n0_20491_4737  0.0142751 
iB30_402_v n1_20583_4784 0  0.0142751 
iB30_402_g 0 n0_20491_4770  0.0142751 
iB30_403_v n1_20771_4535 0  0.0142751 
iB30_403_g 0 n0_20679_4521  0.0142751 
iB30_404_v n1_20771_4568 0  0.0142751 
iB30_404_g 0 n0_20679_4554  0.0142751 
iB30_405_v n1_20771_4751 0  0.0142751 
iB30_405_g 0 n0_20679_4737  0.0142751 
iB30_406_v n1_20771_4784 0  0.0142751 
iB30_406_g 0 n0_20679_4770  0.0142751 
iB30_407_v n1_20583_4967 0  0.0142751 
iB30_407_g 0 n0_20491_4953  0.0142751 
iB30_408_v n1_20583_5000 0  0.0142751 
iB30_408_g 0 n0_20491_4986  0.0142751 
iB30_409_v n1_20583_5183 0  0.0142751 
iB30_409_g 0 n0_20491_5169  0.0142751 
iB30_410_v n1_20583_5216 0  0.0142751 
iB30_410_g 0 n0_20491_5202  0.0142751 
iB30_411_v n1_20630_4967 0  0.0142751 
iB30_411_g 0 n0_20491_4953  0.0142751 
iB30_412_v n1_20630_5000 0  0.0142751 
iB30_412_g 0 n0_20491_4986  0.0142751 
iB30_413_v n1_20771_5000 0  0.0142751 
iB30_413_g 0 n0_20679_5169  0.0142751 
iB30_414_v n1_20771_5183 0  0.0142751 
iB30_414_g 0 n0_20679_5169  0.0142751 
iB30_415_v n1_20771_5216 0  0.0142751 
iB30_415_g 0 n0_20679_5202  0.0142751 
iB12_0_v n1_7083_10799 0  0.0328986 
iB12_0_g 0 n0_6991_10785  0.0328986 
iB12_1_v n1_7083_10832 0  0.0328986 
iB12_1_g 0 n0_6991_10818  0.0328986 
iB12_2_v n1_7271_10799 0  0.0328986 
iB12_2_g 0 n0_7179_10785  0.0328986 
iB12_3_v n1_7271_10832 0  0.0328986 
iB12_3_g 0 n0_7179_10818  0.0328986 
iB12_4_v n1_7083_11015 0  0.0328986 
iB12_4_g 0 n0_6991_11001  0.0328986 
iB12_5_v n1_7083_11048 0  0.0328986 
iB12_5_g 0 n0_6991_11048  0.0328986 
iB12_6_v n1_7083_11204 0  0.0328986 
iB12_6_g 0 n0_6991_11217  0.0328986 
iB12_7_v n1_7083_11231 0  0.0328986 
iB12_7_g 0 n0_6991_11217  0.0328986 
iB12_8_v n1_7083_11264 0  0.0328986 
iB12_8_g 0 n0_6991_11250  0.0328986 
iB12_9_v n1_7271_11015 0  0.0328986 
iB12_9_g 0 n0_7179_11001  0.0328986 
iB12_10_v n1_7271_11048 0  0.0328986 
iB12_10_g 0 n0_7179_11048  0.0328986 
iB12_11_v n1_7271_11204 0  0.0328986 
iB12_11_g 0 n0_7179_11217  0.0328986 
iB12_12_v n1_7271_11231 0  0.0328986 
iB12_12_g 0 n0_7179_11217  0.0328986 
iB12_13_v n1_7271_11264 0  0.0328986 
iB12_13_g 0 n0_7179_11250  0.0328986 
iB12_14_v n1_7083_11447 0  0.0328986 
iB12_14_g 0 n0_6991_11433  0.0328986 
iB12_15_v n1_7083_11480 0  0.0328986 
iB12_15_g 0 n0_6991_11466  0.0328986 
iB12_16_v n1_7083_11663 0  0.0328986 
iB12_16_g 0 n0_6991_11649  0.0328986 
iB12_17_v n1_7083_11696 0  0.0328986 
iB12_17_g 0 n0_6991_11682  0.0328986 
iB12_18_v n1_7130_11663 0  0.0328986 
iB12_18_g 0 n0_6991_11649  0.0328986 
iB12_19_v n1_7130_11696 0  0.0328986 
iB12_19_g 0 n0_6991_11682  0.0328986 
iB12_20_v n1_7271_11447 0  0.0328986 
iB12_20_g 0 n0_7179_11433  0.0328986 
iB12_21_v n1_7271_11480 0  0.0328986 
iB12_21_g 0 n0_7179_11466  0.0328986 
iB12_22_v n1_7271_11663 0  0.0328986 
iB12_22_g 0 n0_7179_11466  0.0328986 
iB12_23_v n1_7271_11696 0  0.0328986 
iB12_23_g 0 n0_7179_11865  0.0328986 
iB12_24_v n1_7083_11879 0  0.0328986 
iB12_24_g 0 n0_6991_11865  0.0328986 
iB12_25_v n1_7083_11912 0  0.0328986 
iB12_25_g 0 n0_6991_11898  0.0328986 
iB12_26_v n1_7083_12095 0  0.0328986 
iB12_26_g 0 n0_6991_12081  0.0328986 
iB12_27_v n1_7083_12128 0  0.0328986 
iB12_27_g 0 n0_6991_12128  0.0328986 
iB12_28_v n1_7271_11879 0  0.0328986 
iB12_28_g 0 n0_7179_11865  0.0328986 
iB12_29_v n1_7271_11912 0  0.0328986 
iB12_29_g 0 n0_7179_11898  0.0328986 
iB12_30_v n1_7271_12095 0  0.0328986 
iB12_30_g 0 n0_7179_12081  0.0328986 
iB12_31_v n1_7271_12128 0  0.0328986 
iB12_31_g 0 n0_7179_12128  0.0328986 
iB12_32_v n1_7083_12284 0  0.0328986 
iB12_32_g 0 n0_6991_12297  0.0328986 
iB12_33_v n1_7083_12311 0  0.0328986 
iB12_33_g 0 n0_6991_12297  0.0328986 
iB12_34_v n1_7083_12344 0  0.0328986 
iB12_34_g 0 n0_6991_12330  0.0328986 
iB12_35_v n1_7083_12527 0  0.0328986 
iB12_35_g 0 n0_6991_12513  0.0328986 
iB12_36_v n1_7083_12560 0  0.0328986 
iB12_36_g 0 n0_6991_12546  0.0328986 
iB12_37_v n1_7271_12284 0  0.0328986 
iB12_37_g 0 n0_7179_12297  0.0328986 
iB12_38_v n1_7271_12311 0  0.0328986 
iB12_38_g 0 n0_7179_12297  0.0328986 
iB12_39_v n1_7271_12344 0  0.0328986 
iB12_39_g 0 n0_7179_12330  0.0328986 
iB12_40_v n1_7271_12527 0  0.0328986 
iB12_40_g 0 n0_7179_12513  0.0328986 
iB12_41_v n1_7271_12560 0  0.0328986 
iB12_41_g 0 n0_7179_12546  0.0328986 
iB12_42_v n1_7083_12743 0  0.0328986 
iB12_42_g 0 n0_6991_12729  0.0328986 
iB12_43_v n1_7083_12959 0  0.0328986 
iB12_43_g 0 n0_6991_12945  0.0328986 
iB12_44_v n1_7083_12992 0  0.0328986 
iB12_44_g 0 n0_6991_12978  0.0328986 
iB12_45_v n1_7271_12743 0  0.0328986 
iB12_45_g 0 n0_7179_12729  0.0328986 
iB12_46_v n1_7271_12776 0  0.0328986 
iB12_46_g 0 n0_7179_12762  0.0328986 
iB12_47_v n1_7271_12959 0  0.0328986 
iB12_47_g 0 n0_7179_12945  0.0328986 
iB12_48_v n1_7271_12992 0  0.0328986 
iB12_48_g 0 n0_7179_12978  0.0328986 
iB12_49_v n1_7083_13175 0  0.0328986 
iB12_49_g 0 n0_6991_13161  0.0328986 
iB12_50_v n1_7083_13208 0  0.0328986 
iB12_50_g 0 n0_6991_13194  0.0328986 
iB12_51_v n1_7083_13391 0  0.0328986 
iB12_51_g 0 n0_6991_13377  0.0328986 
iB12_52_v n1_7083_13424 0  0.0328986 
iB12_52_g 0 n0_6991_13424  0.0328986 
iB12_53_v n1_7271_13175 0  0.0328986 
iB12_53_g 0 n0_7179_13161  0.0328986 
iB12_54_v n1_7271_13208 0  0.0328986 
iB12_54_g 0 n0_7179_13194  0.0328986 
iB12_55_v n1_7271_13391 0  0.0328986 
iB12_55_g 0 n0_7179_13377  0.0328986 
iB12_56_v n1_7271_13424 0  0.0328986 
iB12_56_g 0 n0_7179_13424  0.0328986 
iB12_57_v n1_7083_13580 0  0.0328986 
iB12_57_g 0 n0_6991_13593  0.0328986 
iB12_58_v n1_7083_13607 0  0.0328986 
iB12_58_g 0 n0_6991_13593  0.0328986 
iB12_59_v n1_7083_13640 0  0.0328986 
iB12_59_g 0 n0_6991_13626  0.0328986 
iB12_60_v n1_7083_13823 0  0.0328986 
iB12_60_g 0 n0_6991_13809  0.0328986 
iB12_61_v n1_7083_13856 0  0.0328986 
iB12_61_g 0 n0_6991_13842  0.0328986 
iB12_62_v n1_7271_13580 0  0.0328986 
iB12_62_g 0 n0_7179_13593  0.0328986 
iB12_63_v n1_7271_13607 0  0.0328986 
iB12_63_g 0 n0_7179_13593  0.0328986 
iB12_64_v n1_7271_13640 0  0.0328986 
iB12_64_g 0 n0_7179_13626  0.0328986 
iB12_65_v n1_7271_13823 0  0.0328986 
iB12_65_g 0 n0_7179_13809  0.0328986 
iB12_66_v n1_7271_13856 0  0.0328986 
iB12_66_g 0 n0_7179_13842  0.0328986 
iB12_67_v n1_7083_14039 0  0.0328986 
iB12_67_g 0 n0_6991_13842  0.0328986 
iB12_68_v n1_7083_14072 0  0.0328986 
iB12_68_g 0 n0_6991_13842  0.0328986 
iB12_69_v n1_7083_14255 0  0.0328986 
iB12_69_g 0 n0_6991_13842  0.0328986 
iB12_70_v n1_7130_14039 0  0.0328986 
iB12_70_g 0 n0_7179_13842  0.0328986 
iB12_71_v n1_7271_14039 0  0.0328986 
iB12_71_g 0 n0_7179_13842  0.0328986 
iB12_72_v n1_7271_14072 0  0.0328986 
iB12_72_g 0 n0_7179_13842  0.0328986 
iB12_73_v n1_7271_14255 0  0.0328986 
iB12_73_g 0 n0_7179_13842  0.0328986 
iB12_74_v n1_7083_14288 0  0.0328986 
iB12_74_g 0 n0_6991_13842  0.0328986 
iB12_75_v n1_7083_14471 0  0.0328986 
iB12_75_g 0 n0_6991_13842  0.0328986 
iB12_76_v n1_7083_14504 0  0.0328986 
iB12_76_g 0 n0_6991_13842  0.0328986 
iB12_77_v n1_7083_14553 0  0.0328986 
iB12_77_g 0 n0_6991_13842  0.0328986 
iB12_78_v n1_7271_14288 0  0.0328986 
iB12_78_g 0 n0_7179_13842  0.0328986 
iB12_79_v n1_7271_14471 0  0.0328986 
iB12_79_g 0 n0_7179_13842  0.0328986 
iB12_80_v n1_7271_14504 0  0.0328986 
iB12_80_g 0 n0_7179_13842  0.0328986 
iB12_81_v n1_7271_14553 0  0.0328986 
iB12_81_g 0 n0_7179_13842  0.0328986 
iB12_82_v n1_7083_14687 0  0.0328986 
iB12_82_g 0 n0_6991_13842  0.0328986 
iB12_83_v n1_7083_14720 0  0.0328986 
iB12_83_g 0 n0_6991_13842  0.0328986 
iB12_84_v n1_7083_14903 0  0.0328986 
iB12_84_g 0 n0_8116_14889  0.0328986 
iB12_85_v n1_7083_14936 0  0.0328986 
iB12_85_g 0 n0_8116_14922  0.0328986 
iB12_86_v n1_7271_14687 0  0.0328986 
iB12_86_g 0 n0_7179_13842  0.0328986 
iB12_87_v n1_7271_14720 0  0.0328986 
iB12_87_g 0 n0_7179_13842  0.0328986 
iB12_88_v n1_7271_14903 0  0.0328986 
iB12_88_g 0 n0_8116_14889  0.0328986 
iB12_89_v n1_7271_14936 0  0.0328986 
iB12_89_g 0 n0_8116_14922  0.0328986 
iB12_90_v n1_7083_15335 0  0.0328986 
iB12_90_g 0 n0_6146_15321  0.0328986 
iB12_91_v n1_7083_15368 0  0.0328986 
iB12_91_g 0 n0_6146_15354  0.0328986 
iB12_92_v n1_7271_15119 0  0.0328986 
iB12_92_g 0 n0_8116_15138  0.0328986 
iB12_93_v n1_7271_15152 0  0.0328986 
iB12_93_g 0 n0_8116_15138  0.0328986 
iB12_94_v n1_7271_15335 0  0.0328986 
iB12_94_g 0 n0_8116_15321  0.0328986 
iB12_95_v n1_7271_15368 0  0.0328986 
iB12_95_g 0 n0_8116_15354  0.0328986 
iB12_96_v n1_7083_15551 0  0.0328986 
iB12_96_g 0 n0_6146_15537  0.0328986 
iB12_97_v n1_7083_15584 0  0.0328986 
iB12_97_g 0 n0_6146_15584  0.0328986 
iB12_98_v n1_7083_15740 0  0.0328986 
iB12_98_g 0 n0_6146_15753  0.0328986 
iB12_99_v n1_7083_15767 0  0.0328986 
iB12_99_g 0 n0_6146_15753  0.0328986 
iB12_100_v n1_7083_15800 0  0.0328986 
iB12_100_g 0 n0_6146_15800  0.0328986 
iB12_101_v n1_7271_15551 0  0.0328986 
iB12_101_g 0 n0_8116_15537  0.0328986 
iB12_102_v n1_7271_15584 0  0.0328986 
iB12_102_g 0 n0_8116_15584  0.0328986 
iB12_103_v n1_7271_15740 0  0.0328986 
iB12_103_g 0 n0_8116_15753  0.0328986 
iB12_104_v n1_7271_15767 0  0.0328986 
iB12_104_g 0 n0_8116_15753  0.0328986 
iB12_105_v n1_7271_15800 0  0.0328986 
iB12_105_g 0 n0_8116_15800  0.0328986 
iB12_106_v n1_9333_10799 0  0.0328986 
iB12_106_g 0 n0_9241_10785  0.0328986 
iB12_107_v n1_9333_10832 0  0.0328986 
iB12_107_g 0 n0_9241_10818  0.0328986 
iB12_108_v n1_9333_11015 0  0.0328986 
iB12_108_g 0 n0_9241_11001  0.0328986 
iB12_109_v n1_9333_11048 0  0.0328986 
iB12_109_g 0 n0_9241_11034  0.0328986 
iB12_110_v n1_9333_11231 0  0.0328986 
iB12_110_g 0 n0_9241_11217  0.0328986 
iB12_111_v n1_9333_11264 0  0.0328986 
iB12_111_g 0 n0_9241_11250  0.0328986 
iB12_112_v n1_9333_11447 0  0.0328986 
iB12_112_g 0 n0_9241_11433  0.0328986 
iB12_113_v n1_9333_11480 0  0.0328986 
iB12_113_g 0 n0_9241_11466  0.0328986 
iB12_114_v n1_9333_11663 0  0.0328986 
iB12_114_g 0 n0_9241_11649  0.0328986 
iB12_115_v n1_9333_11696 0  0.0328986 
iB12_115_g 0 n0_9241_11682  0.0328986 
iB12_116_v n1_9333_11879 0  0.0328986 
iB12_116_g 0 n0_9241_11682  0.0328986 
iB12_117_v n1_9333_11912 0  0.0328986 
iB12_117_g 0 n0_9241_11682  0.0328986 
iB12_118_v n1_9333_12095 0  0.0328986 
iB12_118_g 0 n0_9241_11682  0.0328986 
iB12_119_v n1_9333_12128 0  0.0328986 
iB12_119_g 0 n0_9241_11682  0.0328986 
iB12_120_v n1_9333_12311 0  0.0328986 
iB12_120_g 0 n0_9241_11682  0.0328986 
iB12_121_v n1_9333_12344 0  0.0328986 
iB12_121_g 0 n0_9241_11682  0.0328986 
iB12_122_v n1_9333_12527 0  0.0328986 
iB12_122_g 0 n0_9241_11682  0.0328986 
iB12_123_v n1_9333_12560 0  0.0328986 
iB12_123_g 0 n0_9241_11682  0.0328986 
iB12_124_v n1_9333_12743 0  0.0328986 
iB12_124_g 0 n0_8304_12729  0.0328986 
iB12_125_v n1_9333_12959 0  0.0328986 
iB12_125_g 0 n0_8396_12945  0.0328986 
iB12_126_v n1_9333_12992 0  0.0328986 
iB12_126_g 0 n0_8396_12978  0.0328986 
iB12_127_v n1_9333_13175 0  0.0328986 
iB12_127_g 0 n0_8396_13161  0.0328986 
iB12_128_v n1_9333_13208 0  0.0328986 
iB12_128_g 0 n0_8396_13194  0.0328986 
iB12_129_v n1_9333_13391 0  0.0328986 
iB12_129_g 0 n0_8396_13377  0.0328986 
iB12_130_v n1_9333_13424 0  0.0328986 
iB12_130_g 0 n0_8396_13424  0.0328986 
iB12_131_v n1_9333_13607 0  0.0328986 
iB12_131_g 0 n0_8396_13593  0.0328986 
iB12_132_v n1_9333_13640 0  0.0328986 
iB12_132_g 0 n0_8396_13640  0.0328986 
iB12_133_v n1_9333_13796 0  0.0328986 
iB12_133_g 0 n0_8396_13809  0.0328986 
iB12_134_v n1_9333_13823 0  0.0328986 
iB12_134_g 0 n0_8396_13809  0.0328986 
iB12_135_v n1_9333_13856 0  0.0328986 
iB12_135_g 0 n0_8396_13856  0.0328986 
iB12_136_v n1_9333_13990 0  0.0328986 
iB12_136_g 0 n0_8396_14025  0.0328986 
iB12_137_v n1_9333_14012 0  0.0328986 
iB12_137_g 0 n0_8396_14025  0.0328986 
iB12_138_v n1_9333_14039 0  0.0328986 
iB12_138_g 0 n0_8396_14025  0.0328986 
iB12_139_v n1_9333_14072 0  0.0328986 
iB12_139_g 0 n0_8396_14072  0.0328986 
iB12_140_v n1_9333_14228 0  0.0328986 
iB12_140_g 0 n0_8396_14241  0.0328986 
iB12_141_v n1_9333_14255 0  0.0328986 
iB12_141_g 0 n0_8396_14241  0.0328986 
iB12_142_v n1_9333_14288 0  0.0328986 
iB12_142_g 0 n0_8396_14274  0.0328986 
iB12_143_v n1_9333_14471 0  0.0328986 
iB12_143_g 0 n0_8396_14457  0.0328986 
iB12_144_v n1_9333_14504 0  0.0328986 
iB12_144_g 0 n0_8396_14504  0.0328986 
iB12_145_v n1_9333_14660 0  0.0328986 
iB12_145_g 0 n0_8396_14673  0.0328986 
iB12_146_v n1_9333_14687 0  0.0328986 
iB12_146_g 0 n0_8396_14673  0.0328986 
iB12_147_v n1_9333_14720 0  0.0328986 
iB12_147_g 0 n0_8396_14706  0.0328986 
iB12_148_v n1_9333_14903 0  0.0328986 
iB12_148_g 0 n0_8396_14889  0.0328986 
iB12_149_v n1_9333_14936 0  0.0328986 
iB12_149_g 0 n0_8396_14922  0.0328986 
iB12_150_v n1_9333_15335 0  0.0328986 
iB12_150_g 0 n0_8396_15321  0.0328986 
iB12_151_v n1_9333_15368 0  0.0328986 
iB12_151_g 0 n0_8396_15354  0.0328986 
iB12_152_v n1_9333_15551 0  0.0328986 
iB12_152_g 0 n0_8396_15537  0.0328986 
iB12_153_v n1_9333_15584 0  0.0328986 
iB12_153_g 0 n0_8396_15584  0.0328986 
iB12_154_v n1_9333_15740 0  0.0328986 
iB12_154_g 0 n0_8396_15753  0.0328986 
iB12_155_v n1_9333_15767 0  0.0328986 
iB12_155_g 0 n0_8396_15753  0.0328986 
iB12_156_v n1_9333_15800 0  0.0328986 
iB12_156_g 0 n0_8396_15800  0.0328986 
iB12_157_v n1_9333_15934 0  0.0328986 
iB12_157_g 0 n0_8396_15969  0.0328986 
iB12_158_v n1_9521_10799 0  0.0328986 
iB12_158_g 0 n0_9429_10785  0.0328986 
iB12_159_v n1_9521_10832 0  0.0328986 
iB12_159_g 0 n0_9429_10818  0.0328986 
iB12_160_v n1_9521_11015 0  0.0328986 
iB12_160_g 0 n0_9429_11001  0.0328986 
iB12_161_v n1_9521_11048 0  0.0328986 
iB12_161_g 0 n0_9429_11034  0.0328986 
iB12_162_v n1_9521_11231 0  0.0328986 
iB12_162_g 0 n0_9429_11217  0.0328986 
iB12_163_v n1_9521_11264 0  0.0328986 
iB12_163_g 0 n0_9429_11250  0.0328986 
iB12_164_v n1_9380_11663 0  0.0328986 
iB12_164_g 0 n0_9241_11649  0.0328986 
iB12_165_v n1_9380_11696 0  0.0328986 
iB12_165_g 0 n0_9241_11682  0.0328986 
iB12_166_v n1_9521_11447 0  0.0328986 
iB12_166_g 0 n0_9429_11433  0.0328986 
iB12_167_v n1_9521_11480 0  0.0328986 
iB12_167_g 0 n0_9429_11466  0.0328986 
iB12_168_v n1_9521_11663 0  0.0328986 
iB12_168_g 0 n0_9429_11466  0.0328986 
iB12_169_v n1_9521_11696 0  0.0328986 
iB12_169_g 0 n0_9241_11682  0.0328986 
iB12_170_v n1_9521_11879 0  0.0328986 
iB12_170_g 0 n0_9241_11682  0.0328986 
iB12_171_v n1_9521_11912 0  0.0328986 
iB12_171_g 0 n0_9241_11682  0.0328986 
iB12_172_v n1_9521_12095 0  0.0328986 
iB12_172_g 0 n0_9241_11682  0.0328986 
iB12_173_v n1_9521_12128 0  0.0328986 
iB12_173_g 0 n0_9241_11682  0.0328986 
iB12_174_v n1_9521_12311 0  0.0328986 
iB12_174_g 0 n0_10366_12297  0.0328986 
iB12_175_v n1_9521_12344 0  0.0328986 
iB12_175_g 0 n0_10366_12330  0.0328986 
iB12_176_v n1_9521_12527 0  0.0328986 
iB12_176_g 0 n0_10366_12513  0.0328986 
iB12_177_v n1_9521_12560 0  0.0328986 
iB12_177_g 0 n0_10366_12566  0.0328986 
iB12_178_v n1_9521_12743 0  0.0328986 
iB12_178_g 0 n0_10366_12729  0.0328986 
iB12_179_v n1_9521_12776 0  0.0328986 
iB12_179_g 0 n0_10366_12762  0.0328986 
iB12_180_v n1_9521_12959 0  0.0328986 
iB12_180_g 0 n0_10366_12945  0.0328986 
iB12_181_v n1_9521_12992 0  0.0328986 
iB12_181_g 0 n0_10366_12978  0.0328986 
iB12_182_v n1_9521_13175 0  0.0328986 
iB12_182_g 0 n0_10366_13161  0.0328986 
iB12_183_v n1_9521_13208 0  0.0328986 
iB12_183_g 0 n0_10366_13194  0.0328986 
iB12_184_v n1_9521_13391 0  0.0328986 
iB12_184_g 0 n0_10366_13377  0.0328986 
iB12_185_v n1_9521_13424 0  0.0328986 
iB12_185_g 0 n0_10366_13410  0.0328986 
iB12_186_v n1_9521_13607 0  0.0328986 
iB12_186_g 0 n0_10366_13593  0.0328986 
iB12_187_v n1_9521_13640 0  0.0328986 
iB12_187_g 0 n0_10366_13640  0.0328986 
iB12_188_v n1_9521_13796 0  0.0328986 
iB12_188_g 0 n0_10366_13809  0.0328986 
iB12_189_v n1_9521_13823 0  0.0328986 
iB12_189_g 0 n0_10366_13809  0.0328986 
iB12_190_v n1_9521_13856 0  0.0328986 
iB12_190_g 0 n0_10366_13856  0.0328986 
iB12_191_v n1_9380_13990 0  0.0328986 
iB12_191_g 0 n0_8396_14025  0.0328986 
iB12_192_v n1_9380_14012 0  0.0328986 
iB12_192_g 0 n0_8396_14025  0.0328986 
iB12_193_v n1_9380_14039 0  0.0328986 
iB12_193_g 0 n0_8396_14025  0.0328986 
iB12_194_v n1_9521_13990 0  0.0328986 
iB12_194_g 0 n0_10366_14025  0.0328986 
iB12_195_v n1_9521_14012 0  0.0328986 
iB12_195_g 0 n0_10366_14025  0.0328986 
iB12_196_v n1_9521_14039 0  0.0328986 
iB12_196_g 0 n0_10366_14025  0.0328986 
iB12_197_v n1_9521_14072 0  0.0328986 
iB12_197_g 0 n0_10366_14072  0.0328986 
iB12_198_v n1_9521_14228 0  0.0328986 
iB12_198_g 0 n0_10366_14241  0.0328986 
iB12_199_v n1_9521_14255 0  0.0328986 
iB12_199_g 0 n0_10366_14241  0.0328986 
iB12_200_v n1_9521_14288 0  0.0328986 
iB12_200_g 0 n0_10366_14274  0.0328986 
iB12_201_v n1_9521_14471 0  0.0328986 
iB12_201_g 0 n0_10366_14457  0.0328986 
iB12_202_v n1_9521_14504 0  0.0328986 
iB12_202_g 0 n0_10366_14504  0.0328986 
iB12_203_v n1_9521_14660 0  0.0328986 
iB12_203_g 0 n0_10366_14673  0.0328986 
iB12_204_v n1_9521_14687 0  0.0328986 
iB12_204_g 0 n0_10366_14673  0.0328986 
iB12_205_v n1_9521_14720 0  0.0328986 
iB12_205_g 0 n0_10366_14706  0.0328986 
iB12_206_v n1_9521_14903 0  0.0328986 
iB12_206_g 0 n0_10366_14889  0.0328986 
iB12_207_v n1_9521_14936 0  0.0328986 
iB12_207_g 0 n0_10366_14922  0.0328986 
iB12_208_v n1_9521_15119 0  0.0328986 
iB12_208_g 0 n0_10366_15138  0.0328986 
iB12_209_v n1_9521_15152 0  0.0328986 
iB12_209_g 0 n0_10366_15138  0.0328986 
iB12_210_v n1_9521_15335 0  0.0328986 
iB12_210_g 0 n0_10366_15321  0.0328986 
iB12_211_v n1_9521_15368 0  0.0328986 
iB12_211_g 0 n0_10366_15354  0.0328986 
iB12_212_v n1_9521_15551 0  0.0328986 
iB12_212_g 0 n0_10366_15537  0.0328986 
iB12_213_v n1_9521_15584 0  0.0328986 
iB12_213_g 0 n0_10366_15584  0.0328986 
iB12_214_v n1_9521_15740 0  0.0328986 
iB12_214_g 0 n0_10366_15753  0.0328986 
iB12_215_v n1_9521_15767 0  0.0328986 
iB12_215_g 0 n0_10366_15753  0.0328986 
iB12_216_v n1_9521_15800 0  0.0328986 
iB12_216_g 0 n0_10366_15800  0.0328986 
iB12_217_v n1_9521_15934 0  0.0328986 
iB12_217_g 0 n0_10366_15969  0.0328986 
iB31_0_v n1_16083_5350 0  0.0218109 
iB31_0_g 0 n0_15991_5385  0.0218109 
iB31_1_v n1_16083_5399 0  0.0218109 
iB31_1_g 0 n0_15991_5385  0.0218109 
iB31_2_v n1_16083_5432 0  0.0218109 
iB31_2_g 0 n0_15991_5418  0.0218109 
iB31_3_v n1_16083_5566 0  0.0218109 
iB31_3_g 0 n0_15991_5601  0.0218109 
iB31_4_v n1_16083_5615 0  0.0218109 
iB31_4_g 0 n0_15991_5601  0.0218109 
iB31_5_v n1_16083_5648 0  0.0218109 
iB31_5_g 0 n0_15991_5634  0.0218109 
iB31_6_v n1_16083_5831 0  0.0218109 
iB31_6_g 0 n0_15991_5817  0.0218109 
iB31_7_v n1_16083_5864 0  0.0218109 
iB31_7_g 0 n0_15991_5850  0.0218109 
iB31_8_v n1_16083_6263 0  0.0218109 
iB31_8_g 0 n0_15991_6249  0.0218109 
iB31_9_v n1_16083_6296 0  0.0218109 
iB31_9_g 0 n0_15991_6282  0.0218109 
iB31_10_v n1_16083_6333 0  0.0218109 
iB31_10_g 0 n0_15991_6319  0.0218109 
iB31_11_v n1_16083_6430 0  0.0218109 
iB31_11_g 0 n0_15991_6465  0.0218109 
iB31_12_v n1_16083_6479 0  0.0218109 
iB31_12_g 0 n0_15991_6465  0.0218109 
iB31_13_v n1_16083_6512 0  0.0218109 
iB31_13_g 0 n0_15991_6498  0.0218109 
iB31_14_v n1_16083_6695 0  0.0218109 
iB31_14_g 0 n0_15991_6681  0.0218109 
iB31_15_v n1_16083_6728 0  0.0218109 
iB31_15_g 0 n0_15991_6714  0.0218109 
iB31_16_v n1_16083_6911 0  0.0218109 
iB31_16_g 0 n0_15991_6897  0.0218109 
iB31_17_v n1_16083_6944 0  0.0218109 
iB31_17_g 0 n0_15991_6930  0.0218109 
iB31_18_v n1_16083_7127 0  0.0218109 
iB31_18_g 0 n0_15991_7113  0.0218109 
iB31_19_v n1_16083_7160 0  0.0218109 
iB31_19_g 0 n0_15991_7146  0.0218109 
iB31_20_v n1_16130_7160 0  0.0218109 
iB31_20_g 0 n0_16179_7113  0.0218109 
iB31_21_v n1_16083_7343 0  0.0218109 
iB31_21_g 0 n0_15991_7329  0.0218109 
iB31_22_v n1_16083_7376 0  0.0218109 
iB31_22_g 0 n0_15991_7362  0.0218109 
iB31_23_v n1_16083_7559 0  0.0218109 
iB31_23_g 0 n0_15991_7545  0.0218109 
iB31_24_v n1_16083_7592 0  0.0218109 
iB31_24_g 0 n0_15991_7578  0.0218109 
iB31_25_v n1_16083_7775 0  0.0218109 
iB31_25_g 0 n0_15991_7761  0.0218109 
iB31_26_v n1_16083_7808 0  0.0218109 
iB31_26_g 0 n0_15991_7794  0.0218109 
iB31_27_v n1_16083_7845 0  0.0218109 
iB31_27_g 0 n0_15991_7831  0.0218109 
iB31_28_v n1_16083_7942 0  0.0218109 
iB31_28_g 0 n0_15991_7977  0.0218109 
iB31_29_v n1_16083_7991 0  0.0218109 
iB31_29_g 0 n0_15991_7977  0.0218109 
iB31_30_v n1_16083_8024 0  0.0218109 
iB31_30_g 0 n0_15991_8010  0.0218109 
iB31_31_v n1_16083_8207 0  0.0218109 
iB31_31_g 0 n0_15991_8193  0.0218109 
iB31_32_v n1_16083_8240 0  0.0218109 
iB31_32_g 0 n0_15991_8226  0.0218109 
iB31_33_v n1_16083_8456 0  0.0218109 
iB31_33_g 0 n0_16130_8409  0.0218109 
iB31_34_v n1_16083_8639 0  0.0218109 
iB31_34_g 0 n0_15991_8625  0.0218109 
iB31_35_v n1_16083_8672 0  0.0218109 
iB31_35_g 0 n0_15991_8658  0.0218109 
iB31_36_v n1_16083_8855 0  0.0218109 
iB31_36_g 0 n0_15991_8841  0.0218109 
iB31_37_v n1_16083_8888 0  0.0218109 
iB31_37_g 0 n0_15991_8874  0.0218109 
iB31_38_v n1_16083_8925 0  0.0218109 
iB31_38_g 0 n0_15991_8911  0.0218109 
iB31_39_v n1_16083_9022 0  0.0218109 
iB31_39_g 0 n0_15991_9057  0.0218109 
iB31_40_v n1_16083_9071 0  0.0218109 
iB31_40_g 0 n0_15991_9057  0.0218109 
iB31_41_v n1_16083_9104 0  0.0218109 
iB31_41_g 0 n0_15991_9090  0.0218109 
iB31_42_v n1_16083_9287 0  0.0218109 
iB31_42_g 0 n0_15991_9273  0.0218109 
iB31_43_v n1_16083_9320 0  0.0218109 
iB31_43_g 0 n0_15991_9306  0.0218109 
iB31_44_v n1_16083_9503 0  0.0218109 
iB31_44_g 0 n0_15991_9489  0.0218109 
iB31_45_v n1_16083_9536 0  0.0218109 
iB31_45_g 0 n0_15991_9522  0.0218109 
iB31_46_v n1_16083_9719 0  0.0218109 
iB31_46_g 0 n0_15991_9705  0.0218109 
iB31_47_v n1_16083_9752 0  0.0218109 
iB31_47_g 0 n0_15991_9738  0.0218109 
iB31_48_v n1_16130_9503 0  0.0218109 
iB31_48_g 0 n0_15991_9489  0.0218109 
iB31_49_v n1_16130_9536 0  0.0218109 
iB31_49_g 0 n0_15991_9522  0.0218109 
iB31_50_v n1_16083_9935 0  0.0218109 
iB31_50_g 0 n0_15991_9921  0.0218109 
iB31_51_v n1_16083_9968 0  0.0218109 
iB31_51_g 0 n0_15991_9954  0.0218109 
iB31_52_v n1_16083_10005 0  0.0218109 
iB31_52_g 0 n0_15991_9991  0.0218109 
iB31_53_v n1_16083_10102 0  0.0218109 
iB31_53_g 0 n0_15991_10137  0.0218109 
iB31_54_v n1_16083_10151 0  0.0218109 
iB31_54_g 0 n0_15991_10137  0.0218109 
iB31_55_v n1_16083_10184 0  0.0218109 
iB31_55_g 0 n0_15991_10170  0.0218109 
iB31_56_v n1_16083_10367 0  0.0218109 
iB31_56_g 0 n0_15991_10353  0.0218109 
iB31_57_v n1_16083_10400 0  0.0218109 
iB31_57_g 0 n0_15991_10386  0.0218109 
iB31_58_v n1_16271_5350 0  0.0218109 
iB31_58_g 0 n0_16179_5385  0.0218109 
iB31_59_v n1_16271_5399 0  0.0218109 
iB31_59_g 0 n0_16179_5385  0.0218109 
iB31_60_v n1_16271_5432 0  0.0218109 
iB31_60_g 0 n0_16179_5418  0.0218109 
iB31_61_v n1_16271_5566 0  0.0218109 
iB31_61_g 0 n0_16179_5601  0.0218109 
iB31_62_v n1_16271_5615 0  0.0218109 
iB31_62_g 0 n0_16179_5601  0.0218109 
iB31_63_v n1_16271_5648 0  0.0218109 
iB31_63_g 0 n0_16179_5634  0.0218109 
iB31_64_v n1_16271_5831 0  0.0218109 
iB31_64_g 0 n0_16179_5817  0.0218109 
iB31_65_v n1_16271_5864 0  0.0218109 
iB31_65_g 0 n0_16179_5850  0.0218109 
iB31_66_v n1_16271_6047 0  0.0218109 
iB31_66_g 0 n0_16179_6033  0.0218109 
iB31_67_v n1_16271_6080 0  0.0218109 
iB31_67_g 0 n0_16179_6066  0.0218109 
iB31_68_v n1_16271_6263 0  0.0218109 
iB31_68_g 0 n0_16179_6249  0.0218109 
iB31_69_v n1_16271_6296 0  0.0218109 
iB31_69_g 0 n0_16179_6282  0.0218109 
iB31_70_v n1_16271_6333 0  0.0218109 
iB31_70_g 0 n0_16179_6319  0.0218109 
iB31_71_v n1_16271_6430 0  0.0218109 
iB31_71_g 0 n0_16179_6465  0.0218109 
iB31_72_v n1_16271_6479 0  0.0218109 
iB31_72_g 0 n0_16179_6465  0.0218109 
iB31_73_v n1_16271_6512 0  0.0218109 
iB31_73_g 0 n0_16179_6498  0.0218109 
iB31_74_v n1_16271_6695 0  0.0218109 
iB31_74_g 0 n0_16179_6681  0.0218109 
iB31_75_v n1_16271_6728 0  0.0218109 
iB31_75_g 0 n0_16179_6714  0.0218109 
iB31_76_v n1_16271_6911 0  0.0218109 
iB31_76_g 0 n0_16179_6897  0.0218109 
iB31_77_v n1_16271_6944 0  0.0218109 
iB31_77_g 0 n0_16179_6930  0.0218109 
iB31_78_v n1_16271_7127 0  0.0218109 
iB31_78_g 0 n0_16179_7113  0.0218109 
iB31_79_v n1_16271_7160 0  0.0218109 
iB31_79_g 0 n0_16179_7113  0.0218109 
iB31_80_v n1_16271_7343 0  0.0218109 
iB31_80_g 0 n0_16179_7329  0.0218109 
iB31_81_v n1_16271_7376 0  0.0218109 
iB31_81_g 0 n0_16179_7362  0.0218109 
iB31_82_v n1_16271_7559 0  0.0218109 
iB31_82_g 0 n0_16179_7545  0.0218109 
iB31_83_v n1_16271_7592 0  0.0218109 
iB31_83_g 0 n0_16179_7578  0.0218109 
iB31_84_v n1_16271_7775 0  0.0218109 
iB31_84_g 0 n0_16179_7761  0.0218109 
iB31_85_v n1_16271_7808 0  0.0218109 
iB31_85_g 0 n0_16179_7794  0.0218109 
iB31_86_v n1_16271_7845 0  0.0218109 
iB31_86_g 0 n0_16179_7831  0.0218109 
iB31_87_v n1_16271_7942 0  0.0218109 
iB31_87_g 0 n0_16179_7977  0.0218109 
iB31_88_v n1_16271_7991 0  0.0218109 
iB31_88_g 0 n0_16179_7977  0.0218109 
iB31_89_v n1_16271_8024 0  0.0218109 
iB31_89_g 0 n0_16179_8010  0.0218109 
iB31_90_v n1_16271_8207 0  0.0218109 
iB31_90_g 0 n0_16179_8193  0.0218109 
iB31_91_v n1_16271_8240 0  0.0218109 
iB31_91_g 0 n0_16179_8226  0.0218109 
iB31_92_v n1_16271_8423 0  0.0218109 
iB31_92_g 0 n0_16179_8409  0.0218109 
iB31_93_v n1_16271_8456 0  0.0218109 
iB31_93_g 0 n0_16179_8442  0.0218109 
iB31_94_v n1_16271_8639 0  0.0218109 
iB31_94_g 0 n0_16179_8625  0.0218109 
iB31_95_v n1_16271_8672 0  0.0218109 
iB31_95_g 0 n0_16179_8658  0.0218109 
iB31_96_v n1_16271_8855 0  0.0218109 
iB31_96_g 0 n0_16179_8841  0.0218109 
iB31_97_v n1_16271_8888 0  0.0218109 
iB31_97_g 0 n0_16179_8874  0.0218109 
iB31_98_v n1_16271_8925 0  0.0218109 
iB31_98_g 0 n0_16179_8911  0.0218109 
iB31_99_v n1_16271_9022 0  0.0218109 
iB31_99_g 0 n0_16179_9057  0.0218109 
iB31_100_v n1_16271_9071 0  0.0218109 
iB31_100_g 0 n0_16179_9057  0.0218109 
iB31_101_v n1_16271_9104 0  0.0218109 
iB31_101_g 0 n0_16179_9090  0.0218109 
iB31_102_v n1_16271_9287 0  0.0218109 
iB31_102_g 0 n0_16179_9273  0.0218109 
iB31_103_v n1_16271_9320 0  0.0218109 
iB31_103_g 0 n0_16179_9306  0.0218109 
iB31_104_v n1_16271_9503 0  0.0218109 
iB31_104_g 0 n0_16179_9306  0.0218109 
iB31_105_v n1_16271_9536 0  0.0218109 
iB31_105_g 0 n0_16179_9705  0.0218109 
iB31_106_v n1_16271_9719 0  0.0218109 
iB31_106_g 0 n0_16179_9705  0.0218109 
iB31_107_v n1_16271_9752 0  0.0218109 
iB31_107_g 0 n0_16179_9738  0.0218109 
iB31_108_v n1_16271_9935 0  0.0218109 
iB31_108_g 0 n0_16179_9921  0.0218109 
iB31_109_v n1_16271_9968 0  0.0218109 
iB31_109_g 0 n0_16179_9954  0.0218109 
iB31_110_v n1_16271_10005 0  0.0218109 
iB31_110_g 0 n0_16179_9991  0.0218109 
iB31_111_v n1_16271_10102 0  0.0218109 
iB31_111_g 0 n0_16179_10137  0.0218109 
iB31_112_v n1_16271_10151 0  0.0218109 
iB31_112_g 0 n0_16179_10137  0.0218109 
iB31_113_v n1_16271_10184 0  0.0218109 
iB31_113_g 0 n0_16179_10170  0.0218109 
iB31_114_v n1_16271_10367 0  0.0218109 
iB31_114_g 0 n0_16179_10353  0.0218109 
iB31_115_v n1_16271_10400 0  0.0218109 
iB31_115_g 0 n0_16179_10386  0.0218109 
iB31_116_v n1_16271_10616 0  0.0218109 
iB31_116_g 0 n0_16179_10602  0.0218109 
iB31_117_v n1_18333_5350 0  0.0218109 
iB31_117_g 0 n0_18241_5385  0.0218109 
iB31_118_v n1_18333_5399 0  0.0218109 
iB31_118_g 0 n0_18241_5385  0.0218109 
iB31_119_v n1_18333_5432 0  0.0218109 
iB31_119_g 0 n0_18241_5418  0.0218109 
iB31_120_v n1_18333_5566 0  0.0218109 
iB31_120_g 0 n0_18241_5601  0.0218109 
iB31_121_v n1_18333_5615 0  0.0218109 
iB31_121_g 0 n0_18241_5601  0.0218109 
iB31_122_v n1_18333_5648 0  0.0218109 
iB31_122_g 0 n0_18241_5634  0.0218109 
iB31_123_v n1_18521_5350 0  0.0218109 
iB31_123_g 0 n0_18429_5385  0.0218109 
iB31_124_v n1_18521_5399 0  0.0218109 
iB31_124_g 0 n0_18429_5385  0.0218109 
iB31_125_v n1_18521_5432 0  0.0218109 
iB31_125_g 0 n0_18429_5418  0.0218109 
iB31_126_v n1_18521_5566 0  0.0218109 
iB31_126_g 0 n0_18429_5601  0.0218109 
iB31_127_v n1_18521_5615 0  0.0218109 
iB31_127_g 0 n0_18429_5601  0.0218109 
iB31_128_v n1_18521_5648 0  0.0218109 
iB31_128_g 0 n0_18429_5634  0.0218109 
iB31_129_v n1_18333_5831 0  0.0218109 
iB31_129_g 0 n0_18241_5817  0.0218109 
iB31_130_v n1_18333_5864 0  0.0218109 
iB31_130_g 0 n0_18241_5850  0.0218109 
iB31_131_v n1_18521_5831 0  0.0218109 
iB31_131_g 0 n0_18429_5817  0.0218109 
iB31_132_v n1_18521_5864 0  0.0218109 
iB31_132_g 0 n0_18429_5850  0.0218109 
iB31_133_v n1_18521_6047 0  0.0218109 
iB31_133_g 0 n0_18429_6033  0.0218109 
iB31_134_v n1_18521_6080 0  0.0218109 
iB31_134_g 0 n0_18429_6066  0.0218109 
iB31_135_v n1_18333_6263 0  0.0218109 
iB31_135_g 0 n0_18241_6249  0.0218109 
iB31_136_v n1_18333_6296 0  0.0218109 
iB31_136_g 0 n0_18241_6282  0.0218109 
iB31_137_v n1_18333_6333 0  0.0218109 
iB31_137_g 0 n0_18241_6319  0.0218109 
iB31_138_v n1_18333_6430 0  0.0218109 
iB31_138_g 0 n0_18241_6465  0.0218109 
iB31_139_v n1_18333_6479 0  0.0218109 
iB31_139_g 0 n0_18241_6465  0.0218109 
iB31_140_v n1_18333_6512 0  0.0218109 
iB31_140_g 0 n0_18241_6498  0.0218109 
iB31_141_v n1_18521_6263 0  0.0218109 
iB31_141_g 0 n0_18429_6249  0.0218109 
iB31_142_v n1_18521_6296 0  0.0218109 
iB31_142_g 0 n0_18429_6282  0.0218109 
iB31_143_v n1_18521_6333 0  0.0218109 
iB31_143_g 0 n0_18429_6319  0.0218109 
iB31_144_v n1_18521_6430 0  0.0218109 
iB31_144_g 0 n0_18429_6465  0.0218109 
iB31_145_v n1_18521_6479 0  0.0218109 
iB31_145_g 0 n0_18429_6465  0.0218109 
iB31_146_v n1_18521_6512 0  0.0218109 
iB31_146_g 0 n0_18429_6498  0.0218109 
iB31_147_v n1_18333_6695 0  0.0218109 
iB31_147_g 0 n0_18241_6681  0.0218109 
iB31_148_v n1_18333_6728 0  0.0218109 
iB31_148_g 0 n0_18241_6714  0.0218109 
iB31_149_v n1_18333_6911 0  0.0218109 
iB31_149_g 0 n0_18241_6897  0.0218109 
iB31_150_v n1_18521_6695 0  0.0218109 
iB31_150_g 0 n0_18429_6681  0.0218109 
iB31_151_v n1_18521_6728 0  0.0218109 
iB31_151_g 0 n0_18429_6714  0.0218109 
iB31_152_v n1_18521_6911 0  0.0218109 
iB31_152_g 0 n0_18429_6897  0.0218109 
iB31_153_v n1_18333_6944 0  0.0218109 
iB31_153_g 0 n0_18241_6930  0.0218109 
iB31_154_v n1_18333_7127 0  0.0218109 
iB31_154_g 0 n0_18241_7113  0.0218109 
iB31_155_v n1_18333_7160 0  0.0218109 
iB31_155_g 0 n0_18241_7146  0.0218109 
iB31_156_v n1_18380_7160 0  0.0218109 
iB31_156_g 0 n0_18429_7113  0.0218109 
iB31_157_v n1_18521_6944 0  0.0218109 
iB31_157_g 0 n0_18429_6930  0.0218109 
iB31_158_v n1_18521_7127 0  0.0218109 
iB31_158_g 0 n0_18429_7113  0.0218109 
iB31_159_v n1_18521_7160 0  0.0218109 
iB31_159_g 0 n0_18429_7113  0.0218109 
iB31_160_v n1_18333_7343 0  0.0218109 
iB31_160_g 0 n0_18241_7329  0.0218109 
iB31_161_v n1_18333_7376 0  0.0218109 
iB31_161_g 0 n0_18241_7362  0.0218109 
iB31_162_v n1_18333_7559 0  0.0218109 
iB31_162_g 0 n0_18241_7545  0.0218109 
iB31_163_v n1_18333_7592 0  0.0218109 
iB31_163_g 0 n0_18241_7578  0.0218109 
iB31_164_v n1_18521_7343 0  0.0218109 
iB31_164_g 0 n0_18429_7329  0.0218109 
iB31_165_v n1_18521_7376 0  0.0218109 
iB31_165_g 0 n0_18429_7362  0.0218109 
iB31_166_v n1_18521_7559 0  0.0218109 
iB31_166_g 0 n0_18429_7545  0.0218109 
iB31_167_v n1_18521_7592 0  0.0218109 
iB31_167_g 0 n0_18429_7578  0.0218109 
iB31_168_v n1_18333_7775 0  0.0218109 
iB31_168_g 0 n0_18241_7761  0.0218109 
iB31_169_v n1_18333_7808 0  0.0218109 
iB31_169_g 0 n0_18241_7794  0.0218109 
iB31_170_v n1_18333_7845 0  0.0218109 
iB31_170_g 0 n0_18241_7831  0.0218109 
iB31_171_v n1_18333_7942 0  0.0218109 
iB31_171_g 0 n0_18241_7977  0.0218109 
iB31_172_v n1_18333_7991 0  0.0218109 
iB31_172_g 0 n0_18241_7977  0.0218109 
iB31_173_v n1_18333_8024 0  0.0218109 
iB31_173_g 0 n0_18241_8010  0.0218109 
iB31_174_v n1_18521_7775 0  0.0218109 
iB31_174_g 0 n0_18429_7761  0.0218109 
iB31_175_v n1_18521_7808 0  0.0218109 
iB31_175_g 0 n0_18429_7794  0.0218109 
iB31_176_v n1_18521_7845 0  0.0218109 
iB31_176_g 0 n0_18429_7831  0.0218109 
iB31_177_v n1_18521_7942 0  0.0218109 
iB31_177_g 0 n0_18429_7977  0.0218109 
iB31_178_v n1_18521_7991 0  0.0218109 
iB31_178_g 0 n0_18429_7977  0.0218109 
iB31_179_v n1_18521_8024 0  0.0218109 
iB31_179_g 0 n0_18429_8010  0.0218109 
iB31_180_v n1_18333_8207 0  0.0218109 
iB31_180_g 0 n0_18241_8193  0.0218109 
iB31_181_v n1_18333_8240 0  0.0218109 
iB31_181_g 0 n0_18241_8226  0.0218109 
iB31_182_v n1_18333_8456 0  0.0218109 
iB31_182_g 0 n0_18380_8409  0.0218109 
iB31_183_v n1_18521_8207 0  0.0218109 
iB31_183_g 0 n0_18429_8193  0.0218109 
iB31_184_v n1_18521_8240 0  0.0218109 
iB31_184_g 0 n0_18429_8226  0.0218109 
iB31_185_v n1_18521_8423 0  0.0218109 
iB31_185_g 0 n0_18429_8409  0.0218109 
iB31_186_v n1_18521_8456 0  0.0218109 
iB31_186_g 0 n0_18429_8442  0.0218109 
iB31_187_v n1_18333_8639 0  0.0218109 
iB31_187_g 0 n0_18241_8625  0.0218109 
iB31_188_v n1_18333_8672 0  0.0218109 
iB31_188_g 0 n0_18241_8658  0.0218109 
iB31_189_v n1_18333_8855 0  0.0218109 
iB31_189_g 0 n0_18241_8841  0.0218109 
iB31_190_v n1_18333_8888 0  0.0218109 
iB31_190_g 0 n0_18241_8874  0.0218109 
iB31_191_v n1_18333_8925 0  0.0218109 
iB31_191_g 0 n0_18241_8911  0.0218109 
iB31_192_v n1_18521_8639 0  0.0218109 
iB31_192_g 0 n0_18429_8625  0.0218109 
iB31_193_v n1_18521_8672 0  0.0218109 
iB31_193_g 0 n0_18429_8658  0.0218109 
iB31_194_v n1_18521_8855 0  0.0218109 
iB31_194_g 0 n0_18429_8841  0.0218109 
iB31_195_v n1_18521_8888 0  0.0218109 
iB31_195_g 0 n0_18429_8874  0.0218109 
iB31_196_v n1_18521_8925 0  0.0218109 
iB31_196_g 0 n0_18429_8911  0.0218109 
iB31_197_v n1_18333_9022 0  0.0218109 
iB31_197_g 0 n0_18241_9057  0.0218109 
iB31_198_v n1_18333_9071 0  0.0218109 
iB31_198_g 0 n0_18241_9057  0.0218109 
iB31_199_v n1_18333_9104 0  0.0218109 
iB31_199_g 0 n0_18241_9090  0.0218109 
iB31_200_v n1_18333_9287 0  0.0218109 
iB31_200_g 0 n0_18241_9273  0.0218109 
iB31_201_v n1_18333_9320 0  0.0218109 
iB31_201_g 0 n0_18241_9306  0.0218109 
iB31_202_v n1_18521_9022 0  0.0218109 
iB31_202_g 0 n0_18429_9057  0.0218109 
iB31_203_v n1_18521_9071 0  0.0218109 
iB31_203_g 0 n0_18429_9057  0.0218109 
iB31_204_v n1_18521_9104 0  0.0218109 
iB31_204_g 0 n0_18429_9090  0.0218109 
iB31_205_v n1_18521_9287 0  0.0218109 
iB31_205_g 0 n0_18429_9273  0.0218109 
iB31_206_v n1_18521_9320 0  0.0218109 
iB31_206_g 0 n0_18429_9306  0.0218109 
iB31_207_v n1_18333_9503 0  0.0218109 
iB31_207_g 0 n0_18241_9489  0.0218109 
iB31_208_v n1_18333_9536 0  0.0218109 
iB31_208_g 0 n0_18241_9522  0.0218109 
iB31_209_v n1_18333_9719 0  0.0218109 
iB31_209_g 0 n0_18241_9705  0.0218109 
iB31_210_v n1_18333_9752 0  0.0218109 
iB31_210_g 0 n0_18241_9738  0.0218109 
iB31_211_v n1_18380_9503 0  0.0218109 
iB31_211_g 0 n0_18241_9489  0.0218109 
iB31_212_v n1_18380_9536 0  0.0218109 
iB31_212_g 0 n0_18241_9522  0.0218109 
iB31_213_v n1_18521_9503 0  0.0218109 
iB31_213_g 0 n0_18429_9306  0.0218109 
iB31_214_v n1_18521_9536 0  0.0218109 
iB31_214_g 0 n0_18429_9705  0.0218109 
iB31_215_v n1_18521_9719 0  0.0218109 
iB31_215_g 0 n0_18429_9705  0.0218109 
iB31_216_v n1_18521_9752 0  0.0218109 
iB31_216_g 0 n0_18429_9738  0.0218109 
iB31_217_v n1_18333_9935 0  0.0218109 
iB31_217_g 0 n0_18241_9921  0.0218109 
iB31_218_v n1_18333_9968 0  0.0218109 
iB31_218_g 0 n0_18241_9954  0.0218109 
iB31_219_v n1_18333_10005 0  0.0218109 
iB31_219_g 0 n0_18241_9991  0.0218109 
iB31_220_v n1_18333_10102 0  0.0218109 
iB31_220_g 0 n0_18241_10137  0.0218109 
iB31_221_v n1_18333_10151 0  0.0218109 
iB31_221_g 0 n0_18241_10137  0.0218109 
iB31_222_v n1_18333_10184 0  0.0218109 
iB31_222_g 0 n0_18241_10170  0.0218109 
iB31_223_v n1_18521_9935 0  0.0218109 
iB31_223_g 0 n0_18429_9921  0.0218109 
iB31_224_v n1_18521_9968 0  0.0218109 
iB31_224_g 0 n0_18429_9954  0.0218109 
iB31_225_v n1_18521_10005 0  0.0218109 
iB31_225_g 0 n0_18429_9991  0.0218109 
iB31_226_v n1_18521_10102 0  0.0218109 
iB31_226_g 0 n0_18429_10137  0.0218109 
iB31_227_v n1_18521_10151 0  0.0218109 
iB31_227_g 0 n0_18429_10137  0.0218109 
iB31_228_v n1_18521_10184 0  0.0218109 
iB31_228_g 0 n0_18429_10170  0.0218109 
iB31_229_v n1_18333_10367 0  0.0218109 
iB31_229_g 0 n0_18241_10353  0.0218109 
iB31_230_v n1_18333_10400 0  0.0218109 
iB31_230_g 0 n0_18241_10386  0.0218109 
iB31_231_v n1_18521_10367 0  0.0218109 
iB31_231_g 0 n0_18429_10353  0.0218109 
iB31_232_v n1_18521_10400 0  0.0218109 
iB31_232_g 0 n0_18429_10386  0.0218109 
iB31_233_v n1_18521_10616 0  0.0218109 
iB31_233_g 0 n0_18429_10602  0.0218109 
iB31_234_v n1_20583_5399 0  0.0218109 
iB31_234_g 0 n0_20491_5385  0.0218109 
iB31_235_v n1_20583_5432 0  0.0218109 
iB31_235_g 0 n0_20491_5418  0.0218109 
iB31_236_v n1_20583_5615 0  0.0218109 
iB31_236_g 0 n0_20491_5601  0.0218109 
iB31_237_v n1_20583_5648 0  0.0218109 
iB31_237_g 0 n0_20491_5634  0.0218109 
iB31_238_v n1_20771_5399 0  0.0218109 
iB31_238_g 0 n0_20679_5385  0.0218109 
iB31_239_v n1_20771_5432 0  0.0218109 
iB31_239_g 0 n0_20679_5418  0.0218109 
iB31_240_v n1_20771_5615 0  0.0218109 
iB31_240_g 0 n0_20679_5601  0.0218109 
iB31_241_v n1_20771_5648 0  0.0218109 
iB31_241_g 0 n0_20679_5634  0.0218109 
iB31_242_v n1_20583_5782 0  0.0218109 
iB31_242_g 0 n0_20491_5817  0.0218109 
iB31_243_v n1_20583_5831 0  0.0218109 
iB31_243_g 0 n0_20491_5817  0.0218109 
iB31_244_v n1_20583_5864 0  0.0218109 
iB31_244_g 0 n0_20491_5850  0.0218109 
iB31_245_v n1_20771_5782 0  0.0218109 
iB31_245_g 0 n0_20679_5817  0.0218109 
iB31_246_v n1_20771_5831 0  0.0218109 
iB31_246_g 0 n0_20679_5817  0.0218109 
iB31_247_v n1_20771_5864 0  0.0218109 
iB31_247_g 0 n0_20679_5850  0.0218109 
iB31_248_v n1_20771_6047 0  0.0218109 
iB31_248_g 0 n0_20679_6033  0.0218109 
iB31_249_v n1_20771_6080 0  0.0218109 
iB31_249_g 0 n0_20679_6066  0.0218109 
iB31_250_v n1_20583_6263 0  0.0218109 
iB31_250_g 0 n0_20491_6249  0.0218109 
iB31_251_v n1_20583_6296 0  0.0218109 
iB31_251_g 0 n0_20491_6282  0.0218109 
iB31_252_v n1_20583_6333 0  0.0218109 
iB31_252_g 0 n0_20491_6319  0.0218109 
iB31_253_v n1_20583_6479 0  0.0218109 
iB31_253_g 0 n0_20491_6465  0.0218109 
iB31_254_v n1_20583_6512 0  0.0218109 
iB31_254_g 0 n0_20491_6498  0.0218109 
iB31_255_v n1_20771_6263 0  0.0218109 
iB31_255_g 0 n0_20679_6249  0.0218109 
iB31_256_v n1_20771_6296 0  0.0218109 
iB31_256_g 0 n0_20679_6282  0.0218109 
iB31_257_v n1_20771_6479 0  0.0218109 
iB31_257_g 0 n0_20679_6465  0.0218109 
iB31_258_v n1_20771_6512 0  0.0218109 
iB31_258_g 0 n0_20679_6498  0.0218109 
iB31_259_v n1_20583_6695 0  0.0218109 
iB31_259_g 0 n0_20491_6681  0.0218109 
iB31_260_v n1_20583_6728 0  0.0218109 
iB31_260_g 0 n0_20491_6714  0.0218109 
iB31_261_v n1_20583_6911 0  0.0218109 
iB31_261_g 0 n0_20491_6897  0.0218109 
iB31_262_v n1_20771_6695 0  0.0218109 
iB31_262_g 0 n0_20679_6681  0.0218109 
iB31_263_v n1_20771_6728 0  0.0218109 
iB31_263_g 0 n0_20679_6714  0.0218109 
iB31_264_v n1_20771_6911 0  0.0218109 
iB31_264_g 0 n0_20679_6897  0.0218109 
iB31_265_v n1_20583_6944 0  0.0218109 
iB31_265_g 0 n0_20491_6930  0.0218109 
iB31_266_v n1_20583_7127 0  0.0218109 
iB31_266_g 0 n0_20491_7113  0.0218109 
iB31_267_v n1_20583_7160 0  0.0218109 
iB31_267_g 0 n0_20491_7146  0.0218109 
iB31_268_v n1_20630_7160 0  0.0218109 
iB31_268_g 0 n0_20679_7113  0.0218109 
iB31_269_v n1_20771_6944 0  0.0218109 
iB31_269_g 0 n0_20679_6930  0.0218109 
iB31_270_v n1_20771_7127 0  0.0218109 
iB31_270_g 0 n0_20679_7113  0.0218109 
iB31_271_v n1_20771_7160 0  0.0218109 
iB31_271_g 0 n0_20679_7113  0.0218109 
iB31_272_v n1_20583_7343 0  0.0218109 
iB31_272_g 0 n0_20491_7329  0.0218109 
iB31_273_v n1_20583_7376 0  0.0218109 
iB31_273_g 0 n0_20491_7362  0.0218109 
iB31_274_v n1_20583_7559 0  0.0218109 
iB31_274_g 0 n0_20491_7545  0.0218109 
iB31_275_v n1_20583_7592 0  0.0218109 
iB31_275_g 0 n0_20491_7578  0.0218109 
iB31_276_v n1_20771_7343 0  0.0218109 
iB31_276_g 0 n0_20679_7329  0.0218109 
iB31_277_v n1_20771_7376 0  0.0218109 
iB31_277_g 0 n0_20679_7362  0.0218109 
iB31_278_v n1_20771_7559 0  0.0218109 
iB31_278_g 0 n0_20679_7545  0.0218109 
iB31_279_v n1_20771_7592 0  0.0218109 
iB31_279_g 0 n0_20679_7578  0.0218109 
iB31_280_v n1_20583_7775 0  0.0218109 
iB31_280_g 0 n0_20491_7761  0.0218109 
iB31_281_v n1_20583_7808 0  0.0218109 
iB31_281_g 0 n0_20491_7794  0.0218109 
iB31_282_v n1_20583_7991 0  0.0218109 
iB31_282_g 0 n0_20491_7977  0.0218109 
iB31_283_v n1_20583_8024 0  0.0218109 
iB31_283_g 0 n0_20491_8010  0.0218109 
iB31_284_v n1_20771_7775 0  0.0218109 
iB31_284_g 0 n0_20679_7761  0.0218109 
iB31_285_v n1_20771_7808 0  0.0218109 
iB31_285_g 0 n0_20679_7794  0.0218109 
iB31_286_v n1_20771_7991 0  0.0218109 
iB31_286_g 0 n0_20679_7977  0.0218109 
iB31_287_v n1_20771_8024 0  0.0218109 
iB31_287_g 0 n0_20679_8010  0.0218109 
iB31_288_v n1_20583_8207 0  0.0218109 
iB31_288_g 0 n0_20491_8193  0.0218109 
iB31_289_v n1_20583_8240 0  0.0218109 
iB31_289_g 0 n0_20491_8226  0.0218109 
iB31_290_v n1_20583_8456 0  0.0218109 
iB31_290_g 0 n0_20630_8409  0.0218109 
iB31_291_v n1_20771_8207 0  0.0218109 
iB31_291_g 0 n0_20679_8193  0.0218109 
iB31_292_v n1_20771_8240 0  0.0218109 
iB31_292_g 0 n0_20679_8226  0.0218109 
iB31_293_v n1_20771_8423 0  0.0218109 
iB31_293_g 0 n0_20679_8409  0.0218109 
iB31_294_v n1_20771_8456 0  0.0218109 
iB31_294_g 0 n0_20679_8442  0.0218109 
iB31_295_v n1_20583_8639 0  0.0218109 
iB31_295_g 0 n0_20491_8625  0.0218109 
iB31_296_v n1_20583_8672 0  0.0218109 
iB31_296_g 0 n0_20491_8658  0.0218109 
iB31_297_v n1_20583_8855 0  0.0218109 
iB31_297_g 0 n0_20491_8841  0.0218109 
iB31_298_v n1_20583_8888 0  0.0218109 
iB31_298_g 0 n0_20491_8874  0.0218109 
iB31_299_v n1_20771_8639 0  0.0218109 
iB31_299_g 0 n0_20679_8625  0.0218109 
iB31_300_v n1_20771_8672 0  0.0218109 
iB31_300_g 0 n0_20679_8658  0.0218109 
iB31_301_v n1_20771_8855 0  0.0218109 
iB31_301_g 0 n0_20679_8841  0.0218109 
iB31_302_v n1_20771_8888 0  0.0218109 
iB31_302_g 0 n0_20679_8874  0.0218109 
iB31_303_v n1_20583_9071 0  0.0218109 
iB31_303_g 0 n0_20491_9057  0.0218109 
iB31_304_v n1_20583_9104 0  0.0218109 
iB31_304_g 0 n0_20491_9090  0.0218109 
iB31_305_v n1_20583_9287 0  0.0218109 
iB31_305_g 0 n0_20491_9213  0.0218109 
iB31_306_v n1_20583_9320 0  0.0218109 
iB31_306_g 0 n0_20491_9213  0.0218109 
iB31_307_v n1_20771_9071 0  0.0218109 
iB31_307_g 0 n0_20679_9057  0.0218109 
iB31_308_v n1_20771_9104 0  0.0218109 
iB31_308_g 0 n0_20679_9090  0.0218109 
iB31_309_v n1_20771_9287 0  0.0218109 
iB31_309_g 0 n0_20679_9213  0.0218109 
iB31_310_v n1_20771_9320 0  0.0218109 
iB31_310_g 0 n0_20679_9213  0.0218109 
iB31_311_v n1_20583_9503 0  0.0218109 
iB31_311_g 0 n0_20491_9213  0.0218109 
iB31_312_v n1_20583_9536 0  0.0218109 
iB31_312_g 0 n0_20491_9213  0.0218109 
iB31_313_v n1_20583_9719 0  0.0218109 
iB31_313_g 0 n0_20491_9213  0.0218109 
iB31_314_v n1_20583_9752 0  0.0218109 
iB31_314_g 0 n0_20491_9213  0.0218109 
iB31_315_v n1_20630_9503 0  0.0218109 
iB31_315_g 0 n0_20679_9213  0.0218109 
iB31_316_v n1_20630_9536 0  0.0218109 
iB31_316_g 0 n0_20679_9213  0.0218109 
iB31_317_v n1_20771_9503 0  0.0218109 
iB31_317_g 0 n0_20679_9213  0.0218109 
iB31_318_v n1_20771_9536 0  0.0218109 
iB31_318_g 0 n0_20679_9213  0.0218109 
iB31_319_v n1_20771_9719 0  0.0218109 
iB31_319_g 0 n0_20679_9213  0.0218109 
iB31_320_v n1_20771_9752 0  0.0218109 
iB31_320_g 0 n0_20679_9213  0.0218109 
iB31_321_v n1_20583_9935 0  0.0218109 
iB31_321_g 0 n0_20491_9213  0.0218109 
iB31_322_v n1_20583_9968 0  0.0218109 
iB31_322_g 0 n0_20491_9213  0.0218109 
iB31_323_v n1_20583_10151 0  0.0218109 
iB31_323_g 0 n0_20491_9213  0.0218109 
iB31_324_v n1_20583_10184 0  0.0218109 
iB31_324_g 0 n0_20491_9213  0.0218109 
iB31_325_v n1_20771_9935 0  0.0218109 
iB31_325_g 0 n0_20679_9213  0.0218109 
iB31_326_v n1_20771_9968 0  0.0218109 
iB31_326_g 0 n0_20679_9213  0.0218109 
iB31_327_v n1_20771_10151 0  0.0218109 
iB31_327_g 0 n0_20679_9213  0.0218109 
iB31_328_v n1_20771_10184 0  0.0218109 
iB31_328_g 0 n0_20679_9213  0.0218109 
iB31_329_v n1_20583_10367 0  0.0218109 
iB31_329_g 0 n0_19554_10353  0.0218109 
iB31_330_v n1_20583_10400 0  0.0218109 
iB31_330_g 0 n0_19554_10386  0.0218109 
iB31_331_v n1_20771_10367 0  0.0218109 
iB31_331_g 0 n0_19554_10353  0.0218109 
iB31_332_v n1_20771_10400 0  0.0218109 
iB31_332_g 0 n0_19554_10386  0.0218109 
iB31_333_v n1_20771_10616 0  0.0218109 
iB31_333_g 0 n0_19554_10602  0.0218109 
iB13_0_v n1_6900_18527 0  0.0272331 
iB13_0_g 0 n0_6146_18561  0.0272331 
iB13_1_v n1_6900_18548 0  0.0272331 
iB13_1_g 0 n0_6146_18561  0.0272331 
iB13_2_v n1_6900_18575 0  0.0272331 
iB13_2_g 0 n0_6146_18561  0.0272331 
iB13_3_v n1_6900_18608 0  0.0272331 
iB13_3_g 0 n0_6146_18608  0.0272331 
iB13_4_v n1_6900_18764 0  0.0272331 
iB13_4_g 0 n0_6146_18777  0.0272331 
iB13_5_v n1_6900_18791 0  0.0272331 
iB13_5_g 0 n0_6146_18777  0.0272331 
iB13_6_v n1_6900_18824 0  0.0272331 
iB13_6_g 0 n0_6146_18824  0.0272331 
iB13_7_v n1_6900_19007 0  0.0272331 
iB13_7_g 0 n0_6146_18993  0.0272331 
iB13_8_v n1_6900_19040 0  0.0272331 
iB13_8_g 0 n0_6146_19040  0.0272331 
iB13_9_v n1_6900_19196 0  0.0272331 
iB13_9_g 0 n0_6146_19209  0.0272331 
iB13_10_v n1_6900_19223 0  0.0272331 
iB13_10_g 0 n0_6146_19209  0.0272331 
iB13_11_v n1_6900_19256 0  0.0272331 
iB13_11_g 0 n0_6146_19242  0.0272331 
iB13_12_v n1_6900_19439 0  0.0272331 
iB13_12_g 0 n0_6146_19425  0.0272331 
iB13_13_v n1_6900_19472 0  0.0272331 
iB13_13_g 0 n0_6146_19472  0.0272331 
iB13_14_v n1_6900_19655 0  0.0272331 
iB13_14_g 0 n0_6146_19641  0.0272331 
iB13_15_v n1_6900_19688 0  0.0272331 
iB13_15_g 0 n0_6146_19674  0.0272331 
iB13_16_v n1_6900_19871 0  0.0272331 
iB13_16_g 0 n0_6146_19857  0.0272331 
iB13_17_v n1_6900_19904 0  0.0272331 
iB13_17_g 0 n0_6146_19890  0.0272331 
iB13_18_v n1_6900_20087 0  0.0272331 
iB13_18_g 0 n0_6146_20073  0.0272331 
iB13_19_v n1_6900_20120 0  0.0272331 
iB13_19_g 0 n0_6146_20106  0.0272331 
iB13_20_v n1_6900_20303 0  0.0272331 
iB13_20_g 0 n0_6146_20289  0.0272331 
iB13_21_v n1_6900_20336 0  0.0272331 
iB13_21_g 0 n0_6146_20322  0.0272331 
iB13_22_v n1_6900_20519 0  0.0272331 
iB13_22_g 0 n0_6146_20505  0.0272331 
iB13_23_v n1_6900_20552 0  0.0272331 
iB13_23_g 0 n0_6146_20538  0.0272331 
iB13_24_v n1_6900_20687 0  0.0272331 
iB13_24_g 0 n0_6146_20754  0.0272331 
iB13_25_v n1_6900_20735 0  0.0272331 
iB13_25_g 0 n0_6146_20754  0.0272331 
iB13_26_v n1_6900_20768 0  0.0272331 
iB13_26_g 0 n0_6146_20754  0.0272331 
iB13_27_v n1_6900_20951 0  0.0272331 
iB13_27_g 0 n0_6146_20937  0.0272331 
iB13_28_v n1_6900_20984 0  0.0272331 
iB13_28_g 0 n0_6146_20970  0.0272331 
iB13_29_v n1_7083_15956 0  0.0272331 
iB13_29_g 0 n0_6146_15969  0.0272331 
iB13_30_v n1_7083_15983 0  0.0272331 
iB13_30_g 0 n0_6146_15969  0.0272331 
iB13_31_v n1_7083_16016 0  0.0272331 
iB13_31_g 0 n0_6146_16016  0.0272331 
iB13_32_v n1_7083_16172 0  0.0272331 
iB13_32_g 0 n0_6146_16185  0.0272331 
iB13_33_v n1_7083_16199 0  0.0272331 
iB13_33_g 0 n0_6146_16185  0.0272331 
iB13_34_v n1_7083_16232 0  0.0272331 
iB13_34_g 0 n0_6146_16185  0.0272331 
iB13_35_v n1_7130_16172 0  0.0272331 
iB13_35_g 0 n0_6146_16185  0.0272331 
iB13_36_v n1_7130_16199 0  0.0272331 
iB13_36_g 0 n0_6146_16185  0.0272331 
iB13_37_v n1_7130_16232 0  0.0272331 
iB13_37_g 0 n0_6146_16185  0.0272331 
iB13_38_v n1_7271_15956 0  0.0272331 
iB13_38_g 0 n0_8116_15969  0.0272331 
iB13_39_v n1_7271_15983 0  0.0272331 
iB13_39_g 0 n0_8116_15969  0.0272331 
iB13_40_v n1_7271_16016 0  0.0272331 
iB13_40_g 0 n0_8116_16016  0.0272331 
iB13_41_v n1_7271_16172 0  0.0272331 
iB13_41_g 0 n0_8116_16185  0.0272331 
iB13_42_v n1_7271_16199 0  0.0272331 
iB13_42_g 0 n0_8116_16185  0.0272331 
iB13_43_v n1_7083_16415 0  0.0272331 
iB13_43_g 0 n0_6146_16401  0.0272331 
iB13_44_v n1_7083_16448 0  0.0272331 
iB13_44_g 0 n0_6146_16434  0.0272331 
iB13_45_v n1_7083_16631 0  0.0272331 
iB13_45_g 0 n0_6146_16617  0.0272331 
iB13_46_v n1_7083_16664 0  0.0272331 
iB13_46_g 0 n0_6146_16650  0.0272331 
iB13_47_v n1_7271_16415 0  0.0272331 
iB13_47_g 0 n0_8116_16401  0.0272331 
iB13_48_v n1_7271_16448 0  0.0272331 
iB13_48_g 0 n0_8116_16434  0.0272331 
iB13_49_v n1_7271_16631 0  0.0272331 
iB13_49_g 0 n0_8116_16617  0.0272331 
iB13_50_v n1_7271_16664 0  0.0272331 
iB13_50_g 0 n0_8116_16650  0.0272331 
iB13_51_v n1_7083_16847 0  0.0272331 
iB13_51_g 0 n0_6146_16833  0.0272331 
iB13_52_v n1_7083_16880 0  0.0272331 
iB13_52_g 0 n0_6146_16866  0.0272331 
iB13_53_v n1_7083_17063 0  0.0272331 
iB13_53_g 0 n0_6146_17049  0.0272331 
iB13_54_v n1_7083_17096 0  0.0272331 
iB13_54_g 0 n0_6146_17096  0.0272331 
iB13_55_v n1_7271_16847 0  0.0272331 
iB13_55_g 0 n0_8116_16833  0.0272331 
iB13_56_v n1_7271_16880 0  0.0272331 
iB13_56_g 0 n0_8116_16866  0.0272331 
iB13_57_v n1_7271_17063 0  0.0272331 
iB13_57_g 0 n0_8116_17049  0.0272331 
iB13_58_v n1_7271_17096 0  0.0272331 
iB13_58_g 0 n0_8116_17096  0.0272331 
iB13_59_v n1_7083_17230 0  0.0272331 
iB13_59_g 0 n0_6146_17265  0.0272331 
iB13_60_v n1_7083_17468 0  0.0272331 
iB13_60_g 0 n0_6146_17481  0.0272331 
iB13_61_v n1_7083_17495 0  0.0272331 
iB13_61_g 0 n0_6146_17481  0.0272331 
iB13_62_v n1_7271_17230 0  0.0272331 
iB13_62_g 0 n0_8116_17265  0.0272331 
iB13_63_v n1_7271_17252 0  0.0272331 
iB13_63_g 0 n0_8116_17265  0.0272331 
iB13_64_v n1_7271_17279 0  0.0272331 
iB13_64_g 0 n0_8116_17265  0.0272331 
iB13_65_v n1_7271_17312 0  0.0272331 
iB13_65_g 0 n0_8116_17312  0.0272331 
iB13_66_v n1_7271_17468 0  0.0272331 
iB13_66_g 0 n0_8116_17481  0.0272331 
iB13_67_v n1_7271_17495 0  0.0272331 
iB13_67_g 0 n0_8116_17481  0.0272331 
iB13_68_v n1_7083_17528 0  0.0272331 
iB13_68_g 0 n0_6146_17528  0.0272331 
iB13_69_v n1_7083_17711 0  0.0272331 
iB13_69_g 0 n0_6146_17697  0.0272331 
iB13_70_v n1_7083_17744 0  0.0272331 
iB13_70_g 0 n0_6146_17730  0.0272331 
iB13_71_v n1_7083_17927 0  0.0272331 
iB13_71_g 0 n0_6146_17913  0.0272331 
iB13_72_v n1_7271_17528 0  0.0272331 
iB13_72_g 0 n0_8116_17514  0.0272331 
iB13_73_v n1_7271_17711 0  0.0272331 
iB13_73_g 0 n0_8116_17697  0.0272331 
iB13_74_v n1_7271_17744 0  0.0272331 
iB13_74_g 0 n0_8116_17730  0.0272331 
iB13_75_v n1_7271_17927 0  0.0272331 
iB13_75_g 0 n0_8116_17913  0.0272331 
iB13_76_v n1_7083_17960 0  0.0272331 
iB13_76_g 0 n0_6146_17946  0.0272331 
iB13_77_v n1_7083_18143 0  0.0272331 
iB13_77_g 0 n0_6146_18129  0.0272331 
iB13_78_v n1_7083_18176 0  0.0272331 
iB13_78_g 0 n0_6146_18162  0.0272331 
iB13_79_v n1_7271_17960 0  0.0272331 
iB13_79_g 0 n0_8116_17946  0.0272331 
iB13_80_v n1_7271_18143 0  0.0272331 
iB13_80_g 0 n0_8116_18129  0.0272331 
iB13_81_v n1_7271_18176 0  0.0272331 
iB13_81_g 0 n0_8116_18162  0.0272331 
iB13_82_v n1_7083_18359 0  0.0272331 
iB13_82_g 0 n0_6146_18345  0.0272331 
iB13_83_v n1_7083_18392 0  0.0272331 
iB13_83_g 0 n0_6146_18392  0.0272331 
iB13_84_v n1_7083_18526 0  0.0272331 
iB13_84_g 0 n0_6146_18561  0.0272331 
iB13_85_v n1_7083_18527 0  0.0272331 
iB13_85_g 0 n0_6146_18561  0.0272331 
iB13_86_v n1_7083_18548 0  0.0272331 
iB13_86_g 0 n0_6146_18561  0.0272331 
iB13_87_v n1_7083_18575 0  0.0272331 
iB13_87_g 0 n0_6146_18561  0.0272331 
iB13_88_v n1_7083_18608 0  0.0272331 
iB13_88_g 0 n0_6146_18608  0.0272331 
iB13_89_v n1_7130_18392 0  0.0272331 
iB13_89_g 0 n0_6146_18392  0.0272331 
iB13_90_v n1_7130_18526 0  0.0272331 
iB13_90_g 0 n0_6146_18561  0.0272331 
iB13_91_v n1_7130_18527 0  0.0272331 
iB13_91_g 0 n0_6146_18561  0.0272331 
iB13_92_v n1_7130_18548 0  0.0272331 
iB13_92_g 0 n0_6146_18561  0.0272331 
iB13_93_v n1_7271_18359 0  0.0272331 
iB13_93_g 0 n0_8116_18345  0.0272331 
iB13_94_v n1_7271_18392 0  0.0272331 
iB13_94_g 0 n0_8116_18392  0.0272331 
iB13_95_v n1_7271_18526 0  0.0272331 
iB13_95_g 0 n0_8116_18561  0.0272331 
iB13_96_v n1_7271_18527 0  0.0272331 
iB13_96_g 0 n0_8116_18561  0.0272331 
iB13_97_v n1_7271_18548 0  0.0272331 
iB13_97_g 0 n0_8116_18561  0.0272331 
iB13_98_v n1_7271_18575 0  0.0272331 
iB13_98_g 0 n0_8116_18561  0.0272331 
iB13_99_v n1_7271_18608 0  0.0272331 
iB13_99_g 0 n0_8116_18608  0.0272331 
iB13_100_v n1_7083_18764 0  0.0272331 
iB13_100_g 0 n0_6146_18777  0.0272331 
iB13_101_v n1_7083_18791 0  0.0272331 
iB13_101_g 0 n0_6146_18777  0.0272331 
iB13_102_v n1_7083_18824 0  0.0272331 
iB13_102_g 0 n0_6146_18824  0.0272331 
iB13_103_v n1_7083_19007 0  0.0272331 
iB13_103_g 0 n0_6146_18993  0.0272331 
iB13_104_v n1_7083_19040 0  0.0272331 
iB13_104_g 0 n0_6146_19040  0.0272331 
iB13_105_v n1_7271_18764 0  0.0272331 
iB13_105_g 0 n0_8116_18777  0.0272331 
iB13_106_v n1_7271_18791 0  0.0272331 
iB13_106_g 0 n0_8116_18777  0.0272331 
iB13_107_v n1_7271_18824 0  0.0272331 
iB13_107_g 0 n0_8116_18810  0.0272331 
iB13_108_v n1_7271_19007 0  0.0272331 
iB13_108_g 0 n0_8116_18993  0.0272331 
iB13_109_v n1_7271_19040 0  0.0272331 
iB13_109_g 0 n0_8116_19026  0.0272331 
iB13_110_v n1_7083_19196 0  0.0272331 
iB13_110_g 0 n0_6146_19209  0.0272331 
iB13_111_v n1_7083_19223 0  0.0272331 
iB13_111_g 0 n0_6146_19209  0.0272331 
iB13_112_v n1_7083_19256 0  0.0272331 
iB13_112_g 0 n0_6146_19242  0.0272331 
iB13_113_v n1_7083_19390 0  0.0272331 
iB13_113_g 0 n0_6146_19425  0.0272331 
iB13_114_v n1_7083_19439 0  0.0272331 
iB13_114_g 0 n0_6146_19425  0.0272331 
iB13_115_v n1_7083_19472 0  0.0272331 
iB13_115_g 0 n0_6146_19472  0.0272331 
iB13_116_v n1_7271_19196 0  0.0272331 
iB13_116_g 0 n0_8116_19209  0.0272331 
iB13_117_v n1_7271_19223 0  0.0272331 
iB13_117_g 0 n0_8116_19209  0.0272331 
iB13_118_v n1_7271_19256 0  0.0272331 
iB13_118_g 0 n0_8116_19256  0.0272331 
iB13_119_v n1_7271_19390 0  0.0272331 
iB13_119_g 0 n0_8116_19425  0.0272331 
iB13_120_v n1_7271_19439 0  0.0272331 
iB13_120_g 0 n0_8116_19425  0.0272331 
iB13_121_v n1_7271_19472 0  0.0272331 
iB13_121_g 0 n0_8116_19458  0.0272331 
iB13_122_v n1_7083_19871 0  0.0272331 
iB13_122_g 0 n0_6146_19857  0.0272331 
iB13_123_v n1_7083_19904 0  0.0272331 
iB13_123_g 0 n0_6146_19890  0.0272331 
iB13_124_v n1_7271_19655 0  0.0272331 
iB13_124_g 0 n0_8116_19641  0.0272331 
iB13_125_v n1_7271_19688 0  0.0272331 
iB13_125_g 0 n0_8116_19674  0.0272331 
iB13_126_v n1_7271_19871 0  0.0272331 
iB13_126_g 0 n0_8116_19857  0.0272331 
iB13_127_v n1_7271_19904 0  0.0272331 
iB13_127_g 0 n0_8116_19890  0.0272331 
iB13_128_v n1_7083_20087 0  0.0272331 
iB13_128_g 0 n0_6146_20073  0.0272331 
iB13_129_v n1_7083_20120 0  0.0272331 
iB13_129_g 0 n0_6146_20106  0.0272331 
iB13_130_v n1_7083_20303 0  0.0272331 
iB13_130_g 0 n0_6146_20289  0.0272331 
iB13_131_v n1_7083_20336 0  0.0272331 
iB13_131_g 0 n0_6146_20322  0.0272331 
iB13_132_v n1_7271_20087 0  0.0272331 
iB13_132_g 0 n0_8116_20073  0.0272331 
iB13_133_v n1_7271_20120 0  0.0272331 
iB13_133_g 0 n0_8116_20106  0.0272331 
iB13_134_v n1_7271_20303 0  0.0272331 
iB13_134_g 0 n0_8116_20289  0.0272331 
iB13_135_v n1_7271_20336 0  0.0272331 
iB13_135_g 0 n0_8116_20322  0.0272331 
iB13_136_v n1_7083_20519 0  0.0272331 
iB13_136_g 0 n0_6146_20505  0.0272331 
iB13_137_v n1_7083_20552 0  0.0272331 
iB13_137_g 0 n0_6146_20538  0.0272331 
iB13_138_v n1_7083_20687 0  0.0272331 
iB13_138_g 0 n0_6146_20754  0.0272331 
iB13_139_v n1_7083_20735 0  0.0272331 
iB13_139_g 0 n0_6146_20754  0.0272331 
iB13_140_v n1_7083_20768 0  0.0272331 
iB13_140_g 0 n0_6146_20754  0.0272331 
iB13_141_v n1_7130_20687 0  0.0272331 
iB13_141_g 0 n0_6146_20754  0.0272331 
iB13_142_v n1_7130_20735 0  0.0272331 
iB13_142_g 0 n0_6146_20754  0.0272331 
iB13_143_v n1_7130_20768 0  0.0272331 
iB13_143_g 0 n0_6146_20754  0.0272331 
iB13_144_v n1_7271_20519 0  0.0272331 
iB13_144_g 0 n0_8116_20505  0.0272331 
iB13_145_v n1_7271_20552 0  0.0272331 
iB13_145_g 0 n0_8116_20538  0.0272331 
iB13_146_v n1_7271_20687 0  0.0272331 
iB13_146_g 0 n0_8116_20754  0.0272331 
iB13_147_v n1_7271_20768 0  0.0272331 
iB13_147_g 0 n0_8116_20754  0.0272331 
iB13_148_v n1_7083_20951 0  0.0272331 
iB13_148_g 0 n0_6146_20937  0.0272331 
iB13_149_v n1_7083_20984 0  0.0272331 
iB13_149_g 0 n0_6146_20970  0.0272331 
iB13_150_v n1_7271_20951 0  0.0272331 
iB13_150_g 0 n0_8116_20937  0.0272331 
iB13_151_v n1_7271_20984 0  0.0272331 
iB13_151_g 0 n0_8116_20970  0.0272331 
iB13_152_v n1_7364_18526 0  0.0272331 
iB13_152_g 0 n0_8116_18561  0.0272331 
iB13_153_v n1_7364_18527 0  0.0272331 
iB13_153_g 0 n0_8116_18561  0.0272331 
iB13_154_v n1_7364_18575 0  0.0272331 
iB13_154_g 0 n0_8116_18561  0.0272331 
iB13_155_v n1_7364_18608 0  0.0272331 
iB13_155_g 0 n0_8116_18608  0.0272331 
iB13_156_v n1_7364_18764 0  0.0272331 
iB13_156_g 0 n0_8116_18777  0.0272331 
iB13_157_v n1_7364_18791 0  0.0272331 
iB13_157_g 0 n0_8116_18777  0.0272331 
iB13_158_v n1_7364_18824 0  0.0272331 
iB13_158_g 0 n0_8116_18810  0.0272331 
iB13_159_v n1_7364_19007 0  0.0272331 
iB13_159_g 0 n0_8116_18993  0.0272331 
iB13_160_v n1_7364_19040 0  0.0272331 
iB13_160_g 0 n0_8116_19026  0.0272331 
iB13_161_v n1_7364_19223 0  0.0272331 
iB13_161_g 0 n0_8116_19209  0.0272331 
iB13_162_v n1_7364_19256 0  0.0272331 
iB13_162_g 0 n0_8116_19256  0.0272331 
iB13_163_v n1_7364_19390 0  0.0272331 
iB13_163_g 0 n0_8116_19425  0.0272331 
iB13_164_v n1_7364_19439 0  0.0272331 
iB13_164_g 0 n0_8116_19425  0.0272331 
iB13_165_v n1_7364_19472 0  0.0272331 
iB13_165_g 0 n0_8116_19458  0.0272331 
iB13_166_v n1_7364_19655 0  0.0272331 
iB13_166_g 0 n0_8116_19641  0.0272331 
iB13_167_v n1_7364_19688 0  0.0272331 
iB13_167_g 0 n0_8116_19674  0.0272331 
iB13_168_v n1_7364_19871 0  0.0272331 
iB13_168_g 0 n0_8116_19857  0.0272331 
iB13_169_v n1_7364_19904 0  0.0272331 
iB13_169_g 0 n0_8116_19890  0.0272331 
iB13_170_v n1_7364_20087 0  0.0272331 
iB13_170_g 0 n0_8116_20073  0.0272331 
iB13_171_v n1_7364_20120 0  0.0272331 
iB13_171_g 0 n0_8116_20106  0.0272331 
iB13_172_v n1_7364_20303 0  0.0272331 
iB13_172_g 0 n0_8116_20289  0.0272331 
iB13_173_v n1_7364_20336 0  0.0272331 
iB13_173_g 0 n0_8116_20322  0.0272331 
iB13_174_v n1_7364_20519 0  0.0272331 
iB13_174_g 0 n0_8116_20505  0.0272331 
iB13_175_v n1_7364_20552 0  0.0272331 
iB13_175_g 0 n0_8116_20538  0.0272331 
iB13_176_v n1_7364_20687 0  0.0272331 
iB13_176_g 0 n0_8116_20754  0.0272331 
iB13_177_v n1_7364_20735 0  0.0272331 
iB13_177_g 0 n0_8116_20754  0.0272331 
iB13_178_v n1_7364_20768 0  0.0272331 
iB13_178_g 0 n0_8116_20754  0.0272331 
iB13_179_v n1_7364_20951 0  0.0272331 
iB13_179_g 0 n0_8116_20937  0.0272331 
iB13_180_v n1_7364_20984 0  0.0272331 
iB13_180_g 0 n0_8116_20970  0.0272331 
iB13_181_v n1_9333_15956 0  0.0272331 
iB13_181_g 0 n0_8396_15969  0.0272331 
iB13_182_v n1_9333_15983 0  0.0272331 
iB13_182_g 0 n0_8396_15969  0.0272331 
iB13_183_v n1_9333_16016 0  0.0272331 
iB13_183_g 0 n0_8396_16016  0.0272331 
iB13_184_v n1_9333_16172 0  0.0272331 
iB13_184_g 0 n0_8396_16185  0.0272331 
iB13_185_v n1_9333_16199 0  0.0272331 
iB13_185_g 0 n0_8396_16185  0.0272331 
iB13_186_v n1_9333_16232 0  0.0272331 
iB13_186_g 0 n0_8396_16185  0.0272331 
iB13_187_v n1_9333_16415 0  0.0272331 
iB13_187_g 0 n0_8396_16401  0.0272331 
iB13_188_v n1_9333_16448 0  0.0272331 
iB13_188_g 0 n0_8396_16434  0.0272331 
iB13_189_v n1_9333_16631 0  0.0272331 
iB13_189_g 0 n0_8396_16617  0.0272331 
iB13_190_v n1_9333_16664 0  0.0272331 
iB13_190_g 0 n0_8396_16650  0.0272331 
iB13_191_v n1_9333_16847 0  0.0272331 
iB13_191_g 0 n0_8396_16833  0.0272331 
iB13_192_v n1_9333_16880 0  0.0272331 
iB13_192_g 0 n0_8396_16866  0.0272331 
iB13_193_v n1_9333_17063 0  0.0272331 
iB13_193_g 0 n0_8396_17049  0.0272331 
iB13_194_v n1_9333_17096 0  0.0272331 
iB13_194_g 0 n0_8396_17096  0.0272331 
iB13_195_v n1_9333_17230 0  0.0272331 
iB13_195_g 0 n0_8396_17265  0.0272331 
iB13_196_v n1_9333_17468 0  0.0272331 
iB13_196_g 0 n0_8396_17481  0.0272331 
iB13_197_v n1_9333_17495 0  0.0272331 
iB13_197_g 0 n0_8396_17481  0.0272331 
iB13_198_v n1_9333_17528 0  0.0272331 
iB13_198_g 0 n0_8396_17514  0.0272331 
iB13_199_v n1_9333_17711 0  0.0272331 
iB13_199_g 0 n0_8396_17697  0.0272331 
iB13_200_v n1_9333_17744 0  0.0272331 
iB13_200_g 0 n0_8396_17730  0.0272331 
iB13_201_v n1_9333_17927 0  0.0272331 
iB13_201_g 0 n0_8396_17913  0.0272331 
iB13_202_v n1_9333_17960 0  0.0272331 
iB13_202_g 0 n0_8396_17946  0.0272331 
iB13_203_v n1_9333_18143 0  0.0272331 
iB13_203_g 0 n0_8396_18129  0.0272331 
iB13_204_v n1_9333_18176 0  0.0272331 
iB13_204_g 0 n0_8396_18162  0.0272331 
iB13_205_v n1_9150_18527 0  0.0272331 
iB13_205_g 0 n0_8396_18561  0.0272331 
iB13_206_v n1_9150_18548 0  0.0272331 
iB13_206_g 0 n0_8396_18561  0.0272331 
iB13_207_v n1_9150_18575 0  0.0272331 
iB13_207_g 0 n0_8396_18561  0.0272331 
iB13_208_v n1_9150_18608 0  0.0272331 
iB13_208_g 0 n0_8396_18608  0.0272331 
iB13_209_v n1_9333_18359 0  0.0272331 
iB13_209_g 0 n0_8396_18345  0.0272331 
iB13_210_v n1_9333_18392 0  0.0272331 
iB13_210_g 0 n0_8396_18392  0.0272331 
iB13_211_v n1_9333_18527 0  0.0272331 
iB13_211_g 0 n0_8396_18561  0.0272331 
iB13_212_v n1_9333_18548 0  0.0272331 
iB13_212_g 0 n0_8396_18561  0.0272331 
iB13_213_v n1_9333_18575 0  0.0272331 
iB13_213_g 0 n0_8396_18561  0.0272331 
iB13_214_v n1_9333_18608 0  0.0272331 
iB13_214_g 0 n0_8396_18608  0.0272331 
iB13_215_v n1_9150_18764 0  0.0272331 
iB13_215_g 0 n0_8396_18777  0.0272331 
iB13_216_v n1_9150_18791 0  0.0272331 
iB13_216_g 0 n0_8396_18777  0.0272331 
iB13_217_v n1_9150_18824 0  0.0272331 
iB13_217_g 0 n0_8396_18810  0.0272331 
iB13_218_v n1_9150_19007 0  0.0272331 
iB13_218_g 0 n0_8396_18993  0.0272331 
iB13_219_v n1_9150_19040 0  0.0272331 
iB13_219_g 0 n0_8396_19026  0.0272331 
iB13_220_v n1_9333_18764 0  0.0272331 
iB13_220_g 0 n0_8396_18777  0.0272331 
iB13_221_v n1_9333_18791 0  0.0272331 
iB13_221_g 0 n0_8396_18777  0.0272331 
iB13_222_v n1_9333_18824 0  0.0272331 
iB13_222_g 0 n0_8396_18810  0.0272331 
iB13_223_v n1_9333_19007 0  0.0272331 
iB13_223_g 0 n0_8396_18993  0.0272331 
iB13_224_v n1_9333_19040 0  0.0272331 
iB13_224_g 0 n0_8396_19026  0.0272331 
iB13_225_v n1_9150_19223 0  0.0272331 
iB13_225_g 0 n0_8396_19209  0.0272331 
iB13_226_v n1_9150_19256 0  0.0272331 
iB13_226_g 0 n0_8396_19256  0.0272331 
iB13_227_v n1_9150_19412 0  0.0272331 
iB13_227_g 0 n0_8396_19425  0.0272331 
iB13_228_v n1_9150_19439 0  0.0272331 
iB13_228_g 0 n0_8396_19425  0.0272331 
iB13_229_v n1_9150_19472 0  0.0272331 
iB13_229_g 0 n0_8396_19458  0.0272331 
iB13_230_v n1_9333_19223 0  0.0272331 
iB13_230_g 0 n0_8396_19209  0.0272331 
iB13_231_v n1_9333_19256 0  0.0272331 
iB13_231_g 0 n0_8396_19256  0.0272331 
iB13_232_v n1_9333_19412 0  0.0272331 
iB13_232_g 0 n0_8396_19425  0.0272331 
iB13_233_v n1_9333_19439 0  0.0272331 
iB13_233_g 0 n0_8396_19425  0.0272331 
iB13_234_v n1_9333_19472 0  0.0272331 
iB13_234_g 0 n0_8396_19458  0.0272331 
iB13_235_v n1_9150_19655 0  0.0272331 
iB13_235_g 0 n0_8396_19641  0.0272331 
iB13_236_v n1_9150_19688 0  0.0272331 
iB13_236_g 0 n0_8396_19674  0.0272331 
iB13_237_v n1_9150_19871 0  0.0272331 
iB13_237_g 0 n0_8396_19857  0.0272331 
iB13_238_v n1_9150_19904 0  0.0272331 
iB13_238_g 0 n0_8396_19890  0.0272331 
iB13_239_v n1_9333_19871 0  0.0272331 
iB13_239_g 0 n0_8396_19857  0.0272331 
iB13_240_v n1_9333_19904 0  0.0272331 
iB13_240_g 0 n0_8396_19890  0.0272331 
iB13_241_v n1_9150_20087 0  0.0272331 
iB13_241_g 0 n0_8396_20073  0.0272331 
iB13_242_v n1_9150_20120 0  0.0272331 
iB13_242_g 0 n0_8396_20106  0.0272331 
iB13_243_v n1_9150_20303 0  0.0272331 
iB13_243_g 0 n0_8396_20289  0.0272331 
iB13_244_v n1_9150_20336 0  0.0272331 
iB13_244_g 0 n0_8396_20322  0.0272331 
iB13_245_v n1_9333_20087 0  0.0272331 
iB13_245_g 0 n0_8396_20073  0.0272331 
iB13_246_v n1_9333_20120 0  0.0272331 
iB13_246_g 0 n0_8396_20106  0.0272331 
iB13_247_v n1_9333_20303 0  0.0272331 
iB13_247_g 0 n0_8396_20289  0.0272331 
iB13_248_v n1_9333_20336 0  0.0272331 
iB13_248_g 0 n0_8396_20322  0.0272331 
iB13_249_v n1_9150_20519 0  0.0272331 
iB13_249_g 0 n0_8396_20505  0.0272331 
iB13_250_v n1_9150_20552 0  0.0272331 
iB13_250_g 0 n0_8396_20538  0.0272331 
iB13_251_v n1_9150_20687 0  0.0272331 
iB13_251_g 0 n0_8396_20754  0.0272331 
iB13_252_v n1_9150_20735 0  0.0272331 
iB13_252_g 0 n0_8396_20754  0.0272331 
iB13_253_v n1_9150_20768 0  0.0272331 
iB13_253_g 0 n0_8396_20754  0.0272331 
iB13_254_v n1_9333_20519 0  0.0272331 
iB13_254_g 0 n0_8396_20505  0.0272331 
iB13_255_v n1_9333_20552 0  0.0272331 
iB13_255_g 0 n0_8396_20538  0.0272331 
iB13_256_v n1_9333_20687 0  0.0272331 
iB13_256_g 0 n0_8396_20754  0.0272331 
iB13_257_v n1_9333_20735 0  0.0272331 
iB13_257_g 0 n0_8396_20754  0.0272331 
iB13_258_v n1_9333_20768 0  0.0272331 
iB13_258_g 0 n0_8396_20754  0.0272331 
iB13_259_v n1_9150_20951 0  0.0272331 
iB13_259_g 0 n0_8396_20937  0.0272331 
iB13_260_v n1_9150_20984 0  0.0272331 
iB13_260_g 0 n0_8396_20970  0.0272331 
iB13_261_v n1_9333_20951 0  0.0272331 
iB13_261_g 0 n0_8396_20937  0.0272331 
iB13_262_v n1_9333_20984 0  0.0272331 
iB13_262_g 0 n0_8396_20970  0.0272331 
iB13_263_v n1_9380_16172 0  0.0272331 
iB13_263_g 0 n0_8396_16185  0.0272331 
iB13_264_v n1_9380_16199 0  0.0272331 
iB13_264_g 0 n0_8396_16185  0.0272331 
iB13_265_v n1_9380_16232 0  0.0272331 
iB13_265_g 0 n0_8396_16185  0.0272331 
iB13_266_v n1_9521_15956 0  0.0272331 
iB13_266_g 0 n0_10366_15969  0.0272331 
iB13_267_v n1_9521_15983 0  0.0272331 
iB13_267_g 0 n0_10366_15969  0.0272331 
iB13_268_v n1_9521_16016 0  0.0272331 
iB13_268_g 0 n0_10366_16016  0.0272331 
iB13_269_v n1_9521_16172 0  0.0272331 
iB13_269_g 0 n0_10366_16185  0.0272331 
iB13_270_v n1_9521_16199 0  0.0272331 
iB13_270_g 0 n0_10366_16185  0.0272331 
iB13_271_v n1_9521_16415 0  0.0272331 
iB13_271_g 0 n0_10366_16401  0.0272331 
iB13_272_v n1_9521_16448 0  0.0272331 
iB13_272_g 0 n0_10366_16434  0.0272331 
iB13_273_v n1_9521_16631 0  0.0272331 
iB13_273_g 0 n0_10366_16617  0.0272331 
iB13_274_v n1_9521_16664 0  0.0272331 
iB13_274_g 0 n0_10366_16650  0.0272331 
iB13_275_v n1_9521_16847 0  0.0272331 
iB13_275_g 0 n0_10366_16833  0.0272331 
iB13_276_v n1_9521_16880 0  0.0272331 
iB13_276_g 0 n0_10366_16866  0.0272331 
iB13_277_v n1_9521_17063 0  0.0272331 
iB13_277_g 0 n0_10366_17049  0.0272331 
iB13_278_v n1_9521_17096 0  0.0272331 
iB13_278_g 0 n0_10366_17096  0.0272331 
iB13_279_v n1_9521_17230 0  0.0272331 
iB13_279_g 0 n0_10366_17265  0.0272331 
iB13_280_v n1_9521_17252 0  0.0272331 
iB13_280_g 0 n0_10366_17265  0.0272331 
iB13_281_v n1_9521_17279 0  0.0272331 
iB13_281_g 0 n0_10366_17265  0.0272331 
iB13_282_v n1_9521_17312 0  0.0272331 
iB13_282_g 0 n0_10366_17312  0.0272331 
iB13_283_v n1_9521_17468 0  0.0272331 
iB13_283_g 0 n0_10366_17481  0.0272331 
iB13_284_v n1_9521_17495 0  0.0272331 
iB13_284_g 0 n0_10366_17481  0.0272331 
iB13_285_v n1_9521_17528 0  0.0272331 
iB13_285_g 0 n0_10366_17514  0.0272331 
iB13_286_v n1_9521_17711 0  0.0272331 
iB13_286_g 0 n0_10366_17697  0.0272331 
iB13_287_v n1_9521_17744 0  0.0272331 
iB13_287_g 0 n0_10366_17730  0.0272331 
iB13_288_v n1_9521_17927 0  0.0272331 
iB13_288_g 0 n0_10366_17913  0.0272331 
iB13_289_v n1_9521_17960 0  0.0272331 
iB13_289_g 0 n0_10366_17946  0.0272331 
iB13_290_v n1_9521_18143 0  0.0272331 
iB13_290_g 0 n0_10366_18129  0.0272331 
iB13_291_v n1_9521_18176 0  0.0272331 
iB13_291_g 0 n0_10366_18162  0.0272331 
iB13_292_v n1_9380_18392 0  0.0272331 
iB13_292_g 0 n0_8396_18392  0.0272331 
iB13_293_v n1_9380_18527 0  0.0272331 
iB13_293_g 0 n0_8396_18561  0.0272331 
iB13_294_v n1_9380_18548 0  0.0272331 
iB13_294_g 0 n0_8396_18561  0.0272331 
iB13_295_v n1_9521_18359 0  0.0272331 
iB13_295_g 0 n0_10366_18345  0.0272331 
iB13_296_v n1_9521_18392 0  0.0272331 
iB13_296_g 0 n0_10366_18392  0.0272331 
iB13_297_v n1_9521_18527 0  0.0272331 
iB13_297_g 0 n0_10366_18561  0.0272331 
iB13_298_v n1_9521_18548 0  0.0272331 
iB13_298_g 0 n0_10366_18561  0.0272331 
iB13_299_v n1_9521_18575 0  0.0272331 
iB13_299_g 0 n0_10366_18561  0.0272331 
iB13_300_v n1_9521_18608 0  0.0272331 
iB13_300_g 0 n0_10366_18608  0.0272331 
iB13_301_v n1_9614_18527 0  0.0272331 
iB13_301_g 0 n0_10366_18561  0.0272331 
iB13_302_v n1_9614_18548 0  0.0272331 
iB13_302_g 0 n0_10366_18561  0.0272331 
iB13_303_v n1_9614_18575 0  0.0272331 
iB13_303_g 0 n0_10366_18561  0.0272331 
iB13_304_v n1_9614_18608 0  0.0272331 
iB13_304_g 0 n0_10366_18608  0.0272331 
iB13_305_v n1_9521_18764 0  0.0272331 
iB13_305_g 0 n0_10366_18777  0.0272331 
iB13_306_v n1_9521_18791 0  0.0272331 
iB13_306_g 0 n0_10366_18777  0.0272331 
iB13_307_v n1_9521_18824 0  0.0272331 
iB13_307_g 0 n0_10366_18810  0.0272331 
iB13_308_v n1_9521_19007 0  0.0272331 
iB13_308_g 0 n0_10366_18993  0.0272331 
iB13_309_v n1_9521_19040 0  0.0272331 
iB13_309_g 0 n0_10366_19026  0.0272331 
iB13_310_v n1_9614_18764 0  0.0272331 
iB13_310_g 0 n0_10366_18777  0.0272331 
iB13_311_v n1_9614_18791 0  0.0272331 
iB13_311_g 0 n0_10366_18777  0.0272331 
iB13_312_v n1_9614_18824 0  0.0272331 
iB13_312_g 0 n0_10366_18810  0.0272331 
iB13_313_v n1_9614_19007 0  0.0272331 
iB13_313_g 0 n0_10366_18993  0.0272331 
iB13_314_v n1_9614_19040 0  0.0272331 
iB13_314_g 0 n0_10366_19026  0.0272331 
iB13_315_v n1_9521_19223 0  0.0272331 
iB13_315_g 0 n0_10366_19209  0.0272331 
iB13_316_v n1_9521_19256 0  0.0272331 
iB13_316_g 0 n0_10366_19256  0.0272331 
iB13_317_v n1_9521_19412 0  0.0272331 
iB13_317_g 0 n0_10366_19425  0.0272331 
iB13_318_v n1_9521_19439 0  0.0272331 
iB13_318_g 0 n0_10366_19425  0.0272331 
iB13_319_v n1_9521_19472 0  0.0272331 
iB13_319_g 0 n0_10366_19458  0.0272331 
iB13_320_v n1_9614_19223 0  0.0272331 
iB13_320_g 0 n0_10366_19209  0.0272331 
iB13_321_v n1_9614_19256 0  0.0272331 
iB13_321_g 0 n0_10366_19256  0.0272331 
iB13_322_v n1_9614_19412 0  0.0272331 
iB13_322_g 0 n0_10366_19425  0.0272331 
iB13_323_v n1_9614_19439 0  0.0272331 
iB13_323_g 0 n0_10366_19425  0.0272331 
iB13_324_v n1_9614_19472 0  0.0272331 
iB13_324_g 0 n0_10366_19458  0.0272331 
iB13_325_v n1_9521_19655 0  0.0272331 
iB13_325_g 0 n0_10366_19641  0.0272331 
iB13_326_v n1_9521_19688 0  0.0272331 
iB13_326_g 0 n0_10366_19674  0.0272331 
iB13_327_v n1_9521_19871 0  0.0272331 
iB13_327_g 0 n0_10366_19857  0.0272331 
iB13_328_v n1_9521_19904 0  0.0272331 
iB13_328_g 0 n0_10366_19890  0.0272331 
iB13_329_v n1_9614_19655 0  0.0272331 
iB13_329_g 0 n0_10366_19641  0.0272331 
iB13_330_v n1_9614_19688 0  0.0272331 
iB13_330_g 0 n0_10366_19674  0.0272331 
iB13_331_v n1_9614_19871 0  0.0272331 
iB13_331_g 0 n0_10366_19857  0.0272331 
iB13_332_v n1_9614_19904 0  0.0272331 
iB13_332_g 0 n0_10366_19890  0.0272331 
iB13_333_v n1_9521_20087 0  0.0272331 
iB13_333_g 0 n0_10366_20073  0.0272331 
iB13_334_v n1_9521_20120 0  0.0272331 
iB13_334_g 0 n0_10366_20106  0.0272331 
iB13_335_v n1_9521_20303 0  0.0272331 
iB13_335_g 0 n0_10366_20289  0.0272331 
iB13_336_v n1_9521_20336 0  0.0272331 
iB13_336_g 0 n0_10366_20322  0.0272331 
iB13_337_v n1_9614_20087 0  0.0272331 
iB13_337_g 0 n0_10366_20073  0.0272331 
iB13_338_v n1_9614_20120 0  0.0272331 
iB13_338_g 0 n0_10366_20106  0.0272331 
iB13_339_v n1_9614_20303 0  0.0272331 
iB13_339_g 0 n0_10366_20289  0.0272331 
iB13_340_v n1_9614_20336 0  0.0272331 
iB13_340_g 0 n0_10366_20322  0.0272331 
iB13_341_v n1_9380_20687 0  0.0272331 
iB13_341_g 0 n0_8396_20754  0.0272331 
iB13_342_v n1_9380_20735 0  0.0272331 
iB13_342_g 0 n0_8396_20754  0.0272331 
iB13_343_v n1_9380_20768 0  0.0272331 
iB13_343_g 0 n0_8396_20754  0.0272331 
iB13_344_v n1_9521_20519 0  0.0272331 
iB13_344_g 0 n0_10366_20505  0.0272331 
iB13_345_v n1_9521_20552 0  0.0272331 
iB13_345_g 0 n0_10366_20538  0.0272331 
iB13_346_v n1_9521_20687 0  0.0272331 
iB13_346_g 0 n0_10366_20754  0.0272331 
iB13_347_v n1_9521_20768 0  0.0272331 
iB13_347_g 0 n0_10366_20754  0.0272331 
iB13_348_v n1_9614_20519 0  0.0272331 
iB13_348_g 0 n0_10366_20505  0.0272331 
iB13_349_v n1_9614_20552 0  0.0272331 
iB13_349_g 0 n0_10366_20538  0.0272331 
iB13_350_v n1_9614_20687 0  0.0272331 
iB13_350_g 0 n0_10366_20754  0.0272331 
iB13_351_v n1_9614_20735 0  0.0272331 
iB13_351_g 0 n0_10366_20754  0.0272331 
iB13_352_v n1_9614_20768 0  0.0272331 
iB13_352_g 0 n0_10366_20754  0.0272331 
iB13_353_v n1_9521_20951 0  0.0272331 
iB13_353_g 0 n0_10366_20937  0.0272331 
iB13_354_v n1_9521_20984 0  0.0272331 
iB13_354_g 0 n0_10366_20970  0.0272331 
iB13_355_v n1_9614_20951 0  0.0272331 
iB13_355_g 0 n0_10366_20937  0.0272331 
iB13_356_v n1_9614_20984 0  0.0272331 
iB13_356_g 0 n0_10366_20970  0.0272331 
iB32_0_v n1_16083_10799 0  0.025099 
iB32_0_g 0 n0_15991_10785  0.025099 
iB32_1_v n1_16083_10832 0  0.025099 
iB32_1_g 0 n0_15991_10818  0.025099 
iB32_2_v n1_16083_11015 0  0.025099 
iB32_2_g 0 n0_15991_11001  0.025099 
iB32_3_v n1_16083_11048 0  0.025099 
iB32_3_g 0 n0_15991_11048  0.025099 
iB32_4_v n1_16083_11196 0  0.025099 
iB32_4_g 0 n0_15991_11217  0.025099 
iB32_5_v n1_16083_11204 0  0.025099 
iB32_5_g 0 n0_15991_11217  0.025099 
iB32_6_v n1_16083_11231 0  0.025099 
iB32_6_g 0 n0_15991_11217  0.025099 
iB32_7_v n1_16083_11264 0  0.025099 
iB32_7_g 0 n0_15991_11250  0.025099 
iB32_8_v n1_16083_11447 0  0.025099 
iB32_8_g 0 n0_15991_11433  0.025099 
iB32_9_v n1_16083_11480 0  0.025099 
iB32_9_g 0 n0_15991_11466  0.025099 
iB32_10_v n1_16083_11663 0  0.025099 
iB32_10_g 0 n0_15991_11649  0.025099 
iB32_11_v n1_16083_11696 0  0.025099 
iB32_11_g 0 n0_15991_11682  0.025099 
iB32_12_v n1_16130_11663 0  0.025099 
iB32_12_g 0 n0_15991_11649  0.025099 
iB32_13_v n1_16130_11696 0  0.025099 
iB32_13_g 0 n0_15991_11682  0.025099 
iB32_14_v n1_16083_11879 0  0.025099 
iB32_14_g 0 n0_15991_11865  0.025099 
iB32_15_v n1_16083_11912 0  0.025099 
iB32_15_g 0 n0_15991_11898  0.025099 
iB32_16_v n1_16083_12095 0  0.025099 
iB32_16_g 0 n0_15991_12081  0.025099 
iB32_17_v n1_16083_12128 0  0.025099 
iB32_17_g 0 n0_15991_12128  0.025099 
iB32_18_v n1_16083_12276 0  0.025099 
iB32_18_g 0 n0_15991_12297  0.025099 
iB32_19_v n1_16083_12284 0  0.025099 
iB32_19_g 0 n0_15991_12297  0.025099 
iB32_20_v n1_16083_12311 0  0.025099 
iB32_20_g 0 n0_15991_12297  0.025099 
iB32_21_v n1_16083_12344 0  0.025099 
iB32_21_g 0 n0_15991_12330  0.025099 
iB32_22_v n1_16083_12527 0  0.025099 
iB32_22_g 0 n0_15991_12513  0.025099 
iB32_23_v n1_16083_12560 0  0.025099 
iB32_23_g 0 n0_15991_12546  0.025099 
iB32_24_v n1_16083_12743 0  0.025099 
iB32_24_g 0 n0_16130_12776  0.025099 
iB32_25_v n1_16083_12959 0  0.025099 
iB32_25_g 0 n0_15991_12945  0.025099 
iB32_26_v n1_16083_12992 0  0.025099 
iB32_26_g 0 n0_15991_12992  0.025099 
iB32_27_v n1_16083_13175 0  0.025099 
iB32_27_g 0 n0_15991_13161  0.025099 
iB32_28_v n1_16083_13208 0  0.025099 
iB32_28_g 0 n0_15991_13194  0.025099 
iB32_29_v n1_16083_13391 0  0.025099 
iB32_29_g 0 n0_15991_13377  0.025099 
iB32_30_v n1_16083_13424 0  0.025099 
iB32_30_g 0 n0_15991_13423  0.025099 
iB32_31_v n1_16083_13607 0  0.025099 
iB32_31_g 0 n0_15991_13593  0.025099 
iB32_32_v n1_16083_13640 0  0.025099 
iB32_32_g 0 n0_15991_13647  0.025099 
iB32_33_v n1_16083_13788 0  0.025099 
iB32_33_g 0 n0_15991_13809  0.025099 
iB32_34_v n1_16083_13823 0  0.025099 
iB32_34_g 0 n0_15991_13809  0.025099 
iB32_35_v n1_16083_13856 0  0.025099 
iB32_35_g 0 n0_15991_13842  0.025099 
iB32_36_v n1_16083_14039 0  0.025099 
iB32_36_g 0 n0_15991_14025  0.025099 
iB32_37_v n1_16083_14072 0  0.025099 
iB32_37_g 0 n0_15991_14058  0.025099 
iB32_38_v n1_16083_14255 0  0.025099 
iB32_38_g 0 n0_15991_14241  0.025099 
iB32_39_v n1_16130_14039 0  0.025099 
iB32_39_g 0 n0_15991_14025  0.025099 
iB32_40_v n1_16083_14288 0  0.025099 
iB32_40_g 0 n0_15991_14274  0.025099 
iB32_41_v n1_16083_14471 0  0.025099 
iB32_41_g 0 n0_15991_14457  0.025099 
iB32_42_v n1_16083_14504 0  0.025099 
iB32_42_g 0 n0_15991_14511  0.025099 
iB32_43_v n1_16083_14652 0  0.025099 
iB32_43_g 0 n0_15991_14673  0.025099 
iB32_44_v n1_16083_14687 0  0.025099 
iB32_44_g 0 n0_15991_14673  0.025099 
iB32_45_v n1_16083_14720 0  0.025099 
iB32_45_g 0 n0_15991_14706  0.025099 
iB32_46_v n1_16083_14903 0  0.025099 
iB32_46_g 0 n0_15991_14889  0.025099 
iB32_47_v n1_16083_14936 0  0.025099 
iB32_47_g 0 n0_15991_14943  0.025099 
iB32_48_v n1_16083_15300 0  0.025099 
iB32_48_g 0 n0_15991_15321  0.025099 
iB32_49_v n1_16083_15335 0  0.025099 
iB32_49_g 0 n0_15991_15321  0.025099 
iB32_50_v n1_16083_15368 0  0.025099 
iB32_50_g 0 n0_15991_15354  0.025099 
iB32_51_v n1_16083_15551 0  0.025099 
iB32_51_g 0 n0_15991_15537  0.025099 
iB32_52_v n1_16083_15584 0  0.025099 
iB32_52_g 0 n0_15991_15584  0.025099 
iB32_53_v n1_16083_15740 0  0.025099 
iB32_53_g 0 n0_15991_15753  0.025099 
iB32_54_v n1_16083_15767 0  0.025099 
iB32_54_g 0 n0_15991_15753  0.025099 
iB32_55_v n1_16083_15800 0  0.025099 
iB32_55_g 0 n0_15991_15786  0.025099 
iB32_56_v n1_16271_10799 0  0.025099 
iB32_56_g 0 n0_16179_10785  0.025099 
iB32_57_v n1_16271_10832 0  0.025099 
iB32_57_g 0 n0_16179_10818  0.025099 
iB32_58_v n1_16271_11015 0  0.025099 
iB32_58_g 0 n0_16179_11001  0.025099 
iB32_59_v n1_16271_11048 0  0.025099 
iB32_59_g 0 n0_16179_11048  0.025099 
iB32_60_v n1_16271_11196 0  0.025099 
iB32_60_g 0 n0_16179_11217  0.025099 
iB32_61_v n1_16271_11204 0  0.025099 
iB32_61_g 0 n0_16179_11217  0.025099 
iB32_62_v n1_16271_11231 0  0.025099 
iB32_62_g 0 n0_16179_11217  0.025099 
iB32_63_v n1_16271_11264 0  0.025099 
iB32_63_g 0 n0_16179_11250  0.025099 
iB32_64_v n1_16271_11447 0  0.025099 
iB32_64_g 0 n0_16179_11433  0.025099 
iB32_65_v n1_16271_11480 0  0.025099 
iB32_65_g 0 n0_16179_11466  0.025099 
iB32_66_v n1_16271_11663 0  0.025099 
iB32_66_g 0 n0_16179_11466  0.025099 
iB32_67_v n1_16271_11696 0  0.025099 
iB32_67_g 0 n0_16179_11865  0.025099 
iB32_68_v n1_16271_11879 0  0.025099 
iB32_68_g 0 n0_16179_11865  0.025099 
iB32_69_v n1_16271_11912 0  0.025099 
iB32_69_g 0 n0_16179_11898  0.025099 
iB32_70_v n1_16271_12095 0  0.025099 
iB32_70_g 0 n0_16179_12081  0.025099 
iB32_71_v n1_16271_12128 0  0.025099 
iB32_71_g 0 n0_16179_12128  0.025099 
iB32_72_v n1_16271_12276 0  0.025099 
iB32_72_g 0 n0_16179_12297  0.025099 
iB32_73_v n1_16271_12284 0  0.025099 
iB32_73_g 0 n0_16179_12297  0.025099 
iB32_74_v n1_16271_12311 0  0.025099 
iB32_74_g 0 n0_16179_12297  0.025099 
iB32_75_v n1_16271_12344 0  0.025099 
iB32_75_g 0 n0_16179_12330  0.025099 
iB32_76_v n1_16271_12527 0  0.025099 
iB32_76_g 0 n0_16179_12513  0.025099 
iB32_77_v n1_16271_12560 0  0.025099 
iB32_77_g 0 n0_16179_12546  0.025099 
iB32_78_v n1_16271_12743 0  0.025099 
iB32_78_g 0 n0_16179_12729  0.025099 
iB32_79_v n1_16271_12776 0  0.025099 
iB32_79_g 0 n0_16179_12776  0.025099 
iB32_80_v n1_16271_12959 0  0.025099 
iB32_80_g 0 n0_16179_12945  0.025099 
iB32_81_v n1_16271_12992 0  0.025099 
iB32_81_g 0 n0_16179_12992  0.025099 
iB32_82_v n1_16271_13175 0  0.025099 
iB32_82_g 0 n0_16179_13161  0.025099 
iB32_83_v n1_16271_13208 0  0.025099 
iB32_83_g 0 n0_16179_13194  0.025099 
iB32_84_v n1_16271_13391 0  0.025099 
iB32_84_g 0 n0_16179_13377  0.025099 
iB32_85_v n1_16271_13424 0  0.025099 
iB32_85_g 0 n0_16179_13423  0.025099 
iB32_86_v n1_16271_13607 0  0.025099 
iB32_86_g 0 n0_16179_13593  0.025099 
iB32_87_v n1_16271_13640 0  0.025099 
iB32_87_g 0 n0_16179_13647  0.025099 
iB32_88_v n1_16271_13788 0  0.025099 
iB32_88_g 0 n0_16179_13809  0.025099 
iB32_89_v n1_16271_13823 0  0.025099 
iB32_89_g 0 n0_16179_13809  0.025099 
iB32_90_v n1_16271_13856 0  0.025099 
iB32_90_g 0 n0_16179_13842  0.025099 
iB32_91_v n1_16271_14039 0  0.025099 
iB32_91_g 0 n0_16179_13842  0.025099 
iB32_92_v n1_16271_14072 0  0.025099 
iB32_92_g 0 n0_16179_14241  0.025099 
iB32_93_v n1_16271_14255 0  0.025099 
iB32_93_g 0 n0_16179_14241  0.025099 
iB32_94_v n1_16271_14288 0  0.025099 
iB32_94_g 0 n0_16179_14274  0.025099 
iB32_95_v n1_16271_14471 0  0.025099 
iB32_95_g 0 n0_16179_14457  0.025099 
iB32_96_v n1_16271_14504 0  0.025099 
iB32_96_g 0 n0_16179_14511  0.025099 
iB32_97_v n1_16271_14652 0  0.025099 
iB32_97_g 0 n0_16179_14673  0.025099 
iB32_98_v n1_16271_14687 0  0.025099 
iB32_98_g 0 n0_16179_14673  0.025099 
iB32_99_v n1_16271_14720 0  0.025099 
iB32_99_g 0 n0_16179_14706  0.025099 
iB32_100_v n1_16271_14903 0  0.025099 
iB32_100_g 0 n0_16179_14889  0.025099 
iB32_101_v n1_16271_14936 0  0.025099 
iB32_101_g 0 n0_16179_14943  0.025099 
iB32_102_v n1_16271_15084 0  0.025099 
iB32_102_g 0 n0_16179_15105  0.025099 
iB32_103_v n1_16271_15119 0  0.025099 
iB32_103_g 0 n0_16179_15105  0.025099 
iB32_104_v n1_16271_15152 0  0.025099 
iB32_104_g 0 n0_16179_15159  0.025099 
iB32_105_v n1_16271_15300 0  0.025099 
iB32_105_g 0 n0_16179_15321  0.025099 
iB32_106_v n1_16271_15335 0  0.025099 
iB32_106_g 0 n0_16179_15321  0.025099 
iB32_107_v n1_16271_15368 0  0.025099 
iB32_107_g 0 n0_16179_15354  0.025099 
iB32_108_v n1_16271_15551 0  0.025099 
iB32_108_g 0 n0_16179_15537  0.025099 
iB32_109_v n1_16271_15584 0  0.025099 
iB32_109_g 0 n0_16179_15584  0.025099 
iB32_110_v n1_16271_15740 0  0.025099 
iB32_110_g 0 n0_16179_15753  0.025099 
iB32_111_v n1_16271_15767 0  0.025099 
iB32_111_g 0 n0_16179_15753  0.025099 
iB32_112_v n1_16271_15800 0  0.025099 
iB32_112_g 0 n0_16179_15786  0.025099 
iB32_113_v n1_18333_10799 0  0.025099 
iB32_113_g 0 n0_18241_10785  0.025099 
iB32_114_v n1_18333_10832 0  0.025099 
iB32_114_g 0 n0_18241_10818  0.025099 
iB32_115_v n1_18521_10799 0  0.025099 
iB32_115_g 0 n0_18429_10785  0.025099 
iB32_116_v n1_18521_10832 0  0.025099 
iB32_116_g 0 n0_18429_10818  0.025099 
iB32_117_v n1_18333_11015 0  0.025099 
iB32_117_g 0 n0_18241_11001  0.025099 
iB32_118_v n1_18333_11048 0  0.025099 
iB32_118_g 0 n0_18241_11055  0.025099 
iB32_119_v n1_18333_11196 0  0.025099 
iB32_119_g 0 n0_18241_11217  0.025099 
iB32_120_v n1_18333_11231 0  0.025099 
iB32_120_g 0 n0_18241_11217  0.025099 
iB32_121_v n1_18333_11264 0  0.025099 
iB32_121_g 0 n0_18241_11250  0.025099 
iB32_122_v n1_18521_11015 0  0.025099 
iB32_122_g 0 n0_18429_11001  0.025099 
iB32_123_v n1_18521_11048 0  0.025099 
iB32_123_g 0 n0_18429_11055  0.025099 
iB32_124_v n1_18521_11196 0  0.025099 
iB32_124_g 0 n0_18429_11217  0.025099 
iB32_125_v n1_18521_11231 0  0.025099 
iB32_125_g 0 n0_18429_11217  0.025099 
iB32_126_v n1_18521_11264 0  0.025099 
iB32_126_g 0 n0_18429_11250  0.025099 
iB32_127_v n1_18333_11447 0  0.025099 
iB32_127_g 0 n0_18241_11433  0.025099 
iB32_128_v n1_18333_11480 0  0.025099 
iB32_128_g 0 n0_18241_11466  0.025099 
iB32_129_v n1_18333_11663 0  0.025099 
iB32_129_g 0 n0_18241_11649  0.025099 
iB32_130_v n1_18333_11696 0  0.025099 
iB32_130_g 0 n0_18241_11682  0.025099 
iB32_131_v n1_18380_11663 0  0.025099 
iB32_131_g 0 n0_18241_11649  0.025099 
iB32_132_v n1_18380_11696 0  0.025099 
iB32_132_g 0 n0_18241_11682  0.025099 
iB32_133_v n1_18521_11447 0  0.025099 
iB32_133_g 0 n0_18429_11433  0.025099 
iB32_134_v n1_18521_11480 0  0.025099 
iB32_134_g 0 n0_18429_11466  0.025099 
iB32_135_v n1_18521_11663 0  0.025099 
iB32_135_g 0 n0_18429_11466  0.025099 
iB32_136_v n1_18521_11696 0  0.025099 
iB32_136_g 0 n0_18429_11865  0.025099 
iB32_137_v n1_18333_11879 0  0.025099 
iB32_137_g 0 n0_18241_11865  0.025099 
iB32_138_v n1_18333_11912 0  0.025099 
iB32_138_g 0 n0_18241_11898  0.025099 
iB32_139_v n1_18333_12095 0  0.025099 
iB32_139_g 0 n0_18241_12081  0.025099 
iB32_140_v n1_18333_12128 0  0.025099 
iB32_140_g 0 n0_18241_12128  0.025099 
iB32_141_v n1_18521_11879 0  0.025099 
iB32_141_g 0 n0_18429_11865  0.025099 
iB32_142_v n1_18521_11912 0  0.025099 
iB32_142_g 0 n0_18429_11898  0.025099 
iB32_143_v n1_18521_12095 0  0.025099 
iB32_143_g 0 n0_18429_12081  0.025099 
iB32_144_v n1_18521_12128 0  0.025099 
iB32_144_g 0 n0_18429_12128  0.025099 
iB32_145_v n1_18333_12284 0  0.025099 
iB32_145_g 0 n0_18241_12297  0.025099 
iB32_146_v n1_18333_12311 0  0.025099 
iB32_146_g 0 n0_18241_12297  0.025099 
iB32_147_v n1_18333_12344 0  0.025099 
iB32_147_g 0 n0_18241_12330  0.025099 
iB32_148_v n1_18333_12527 0  0.025099 
iB32_148_g 0 n0_18241_12513  0.025099 
iB32_149_v n1_18333_12560 0  0.025099 
iB32_149_g 0 n0_18241_12546  0.025099 
iB32_150_v n1_18521_12284 0  0.025099 
iB32_150_g 0 n0_18429_12297  0.025099 
iB32_151_v n1_18521_12311 0  0.025099 
iB32_151_g 0 n0_18429_12297  0.025099 
iB32_152_v n1_18521_12344 0  0.025099 
iB32_152_g 0 n0_18429_12330  0.025099 
iB32_153_v n1_18521_12527 0  0.025099 
iB32_153_g 0 n0_18429_12513  0.025099 
iB32_154_v n1_18521_12560 0  0.025099 
iB32_154_g 0 n0_18429_12546  0.025099 
iB32_155_v n1_18333_12743 0  0.025099 
iB32_155_g 0 n0_18241_12729  0.025099 
iB32_156_v n1_18333_12959 0  0.025099 
iB32_156_g 0 n0_18241_12945  0.025099 
iB32_157_v n1_18333_12992 0  0.025099 
iB32_157_g 0 n0_18241_12978  0.025099 
iB32_158_v n1_18521_12743 0  0.025099 
iB32_158_g 0 n0_18429_12729  0.025099 
iB32_159_v n1_18521_12776 0  0.025099 
iB32_159_g 0 n0_18429_12762  0.025099 
iB32_160_v n1_18521_12959 0  0.025099 
iB32_160_g 0 n0_18429_12945  0.025099 
iB32_161_v n1_18521_12992 0  0.025099 
iB32_161_g 0 n0_18429_12978  0.025099 
iB32_162_v n1_18333_13175 0  0.025099 
iB32_162_g 0 n0_18241_13161  0.025099 
iB32_163_v n1_18333_13208 0  0.025099 
iB32_163_g 0 n0_18241_13194  0.025099 
iB32_164_v n1_18333_13391 0  0.025099 
iB32_164_g 0 n0_18241_13377  0.025099 
iB32_165_v n1_18333_13424 0  0.025099 
iB32_165_g 0 n0_18429_13423  0.025099 
iB32_166_v n1_18521_13175 0  0.025099 
iB32_166_g 0 n0_18429_13161  0.025099 
iB32_167_v n1_18521_13208 0  0.025099 
iB32_167_g 0 n0_18429_13194  0.025099 
iB32_168_v n1_18521_13391 0  0.025099 
iB32_168_g 0 n0_18429_13377  0.025099 
iB32_169_v n1_18521_13424 0  0.025099 
iB32_169_g 0 n0_18429_13423  0.025099 
iB32_170_v n1_18333_13607 0  0.025099 
iB32_170_g 0 n0_18241_13593  0.025099 
iB32_171_v n1_18333_13640 0  0.025099 
iB32_171_g 0 n0_18241_13640  0.025099 
iB32_172_v n1_18333_13788 0  0.025099 
iB32_172_g 0 n0_18241_13809  0.025099 
iB32_173_v n1_18333_13796 0  0.025099 
iB32_173_g 0 n0_18241_13809  0.025099 
iB32_174_v n1_18333_13823 0  0.025099 
iB32_174_g 0 n0_18241_13809  0.025099 
iB32_175_v n1_18333_13856 0  0.025099 
iB32_175_g 0 n0_18241_13842  0.025099 
iB32_176_v n1_18521_13607 0  0.025099 
iB32_176_g 0 n0_18429_13593  0.025099 
iB32_177_v n1_18521_13640 0  0.025099 
iB32_177_g 0 n0_18429_13640  0.025099 
iB32_178_v n1_18521_13788 0  0.025099 
iB32_178_g 0 n0_18429_13809  0.025099 
iB32_179_v n1_18521_13796 0  0.025099 
iB32_179_g 0 n0_18429_13809  0.025099 
iB32_180_v n1_18521_13823 0  0.025099 
iB32_180_g 0 n0_18429_13809  0.025099 
iB32_181_v n1_18521_13856 0  0.025099 
iB32_181_g 0 n0_18429_13842  0.025099 
iB32_182_v n1_18333_14039 0  0.025099 
iB32_182_g 0 n0_18241_14025  0.025099 
iB32_183_v n1_18333_14072 0  0.025099 
iB32_183_g 0 n0_18241_14058  0.025099 
iB32_184_v n1_18333_14255 0  0.025099 
iB32_184_g 0 n0_18241_14241  0.025099 
iB32_185_v n1_18380_14039 0  0.025099 
iB32_185_g 0 n0_18241_14025  0.025099 
iB32_186_v n1_18521_14039 0  0.025099 
iB32_186_g 0 n0_18429_13842  0.025099 
iB32_187_v n1_18521_14072 0  0.025099 
iB32_187_g 0 n0_18429_14241  0.025099 
iB32_188_v n1_18521_14255 0  0.025099 
iB32_188_g 0 n0_18429_14241  0.025099 
iB32_189_v n1_18333_14288 0  0.025099 
iB32_189_g 0 n0_18241_14274  0.025099 
iB32_190_v n1_18333_14471 0  0.025099 
iB32_190_g 0 n0_18241_14457  0.025099 
iB32_191_v n1_18333_14504 0  0.025099 
iB32_191_g 0 n0_18241_14504  0.025099 
iB32_192_v n1_18333_14652 0  0.025099 
iB32_192_g 0 n0_18241_14673  0.025099 
iB32_193_v n1_18333_14660 0  0.025099 
iB32_193_g 0 n0_18241_14673  0.025099 
iB32_194_v n1_18521_14288 0  0.025099 
iB32_194_g 0 n0_18429_14274  0.025099 
iB32_195_v n1_18521_14471 0  0.025099 
iB32_195_g 0 n0_18429_14457  0.025099 
iB32_196_v n1_18521_14504 0  0.025099 
iB32_196_g 0 n0_18429_14504  0.025099 
iB32_197_v n1_18521_14652 0  0.025099 
iB32_197_g 0 n0_18429_14673  0.025099 
iB32_198_v n1_18521_14660 0  0.025099 
iB32_198_g 0 n0_18429_14673  0.025099 
iB32_199_v n1_18333_14687 0  0.025099 
iB32_199_g 0 n0_18241_14673  0.025099 
iB32_200_v n1_18333_14720 0  0.025099 
iB32_200_g 0 n0_18241_14706  0.025099 
iB32_201_v n1_18333_14903 0  0.025099 
iB32_201_g 0 n0_18241_14889  0.025099 
iB32_202_v n1_18333_14936 0  0.025099 
iB32_202_g 0 n0_18241_14936  0.025099 
iB32_203_v n1_18521_14687 0  0.025099 
iB32_203_g 0 n0_18429_14673  0.025099 
iB32_204_v n1_18521_14720 0  0.025099 
iB32_204_g 0 n0_18429_14706  0.025099 
iB32_205_v n1_18521_14903 0  0.025099 
iB32_205_g 0 n0_18429_14889  0.025099 
iB32_206_v n1_18521_14936 0  0.025099 
iB32_206_g 0 n0_18429_14936  0.025099 
iB32_207_v n1_18333_15308 0  0.025099 
iB32_207_g 0 n0_18241_15321  0.025099 
iB32_208_v n1_18333_15335 0  0.025099 
iB32_208_g 0 n0_18241_15321  0.025099 
iB32_209_v n1_18333_15368 0  0.025099 
iB32_209_g 0 n0_18241_15354  0.025099 
iB32_210_v n1_18521_15092 0  0.025099 
iB32_210_g 0 n0_18429_15105  0.025099 
iB32_211_v n1_18521_15119 0  0.025099 
iB32_211_g 0 n0_18429_15105  0.025099 
iB32_212_v n1_18521_15152 0  0.025099 
iB32_212_g 0 n0_18429_15152  0.025099 
iB32_213_v n1_18521_15308 0  0.025099 
iB32_213_g 0 n0_18429_15321  0.025099 
iB32_214_v n1_18521_15335 0  0.025099 
iB32_214_g 0 n0_18429_15321  0.025099 
iB32_215_v n1_18521_15368 0  0.025099 
iB32_215_g 0 n0_18429_15354  0.025099 
iB32_216_v n1_18333_15551 0  0.025099 
iB32_216_g 0 n0_18241_15537  0.025099 
iB32_217_v n1_18333_15584 0  0.025099 
iB32_217_g 0 n0_18241_15584  0.025099 
iB32_218_v n1_18333_15740 0  0.025099 
iB32_218_g 0 n0_18241_15753  0.025099 
iB32_219_v n1_18333_15767 0  0.025099 
iB32_219_g 0 n0_18241_15753  0.025099 
iB32_220_v n1_18333_15800 0  0.025099 
iB32_220_g 0 n0_18241_15786  0.025099 
iB32_221_v n1_18521_15551 0  0.025099 
iB32_221_g 0 n0_18429_15537  0.025099 
iB32_222_v n1_18521_15584 0  0.025099 
iB32_222_g 0 n0_18429_15584  0.025099 
iB32_223_v n1_18521_15740 0  0.025099 
iB32_223_g 0 n0_18429_15753  0.025099 
iB32_224_v n1_18521_15767 0  0.025099 
iB32_224_g 0 n0_18429_15753  0.025099 
iB32_225_v n1_18521_15800 0  0.025099 
iB32_225_g 0 n0_18429_15786  0.025099 
iB32_226_v n1_20583_10799 0  0.025099 
iB32_226_g 0 n0_19554_10785  0.025099 
iB32_227_v n1_20583_10832 0  0.025099 
iB32_227_g 0 n0_19554_10818  0.025099 
iB32_228_v n1_20771_10799 0  0.025099 
iB32_228_g 0 n0_19554_10785  0.025099 
iB32_229_v n1_20771_10832 0  0.025099 
iB32_229_g 0 n0_20679_11956  0.025099 
iB32_230_v n1_20583_11015 0  0.025099 
iB32_230_g 0 n0_20491_11956  0.025099 
iB32_231_v n1_20583_11048 0  0.025099 
iB32_231_g 0 n0_20491_11956  0.025099 
iB32_232_v n1_20583_11231 0  0.025099 
iB32_232_g 0 n0_20491_11956  0.025099 
iB32_233_v n1_20583_11264 0  0.025099 
iB32_233_g 0 n0_20491_11956  0.025099 
iB32_234_v n1_20771_11015 0  0.025099 
iB32_234_g 0 n0_20679_11956  0.025099 
iB32_235_v n1_20771_11048 0  0.025099 
iB32_235_g 0 n0_20679_11956  0.025099 
iB32_236_v n1_20771_11231 0  0.025099 
iB32_236_g 0 n0_20679_11956  0.025099 
iB32_237_v n1_20771_11264 0  0.025099 
iB32_237_g 0 n0_20679_11956  0.025099 
iB32_238_v n1_20583_11447 0  0.025099 
iB32_238_g 0 n0_20491_11956  0.025099 
iB32_239_v n1_20583_11480 0  0.025099 
iB32_239_g 0 n0_20491_11956  0.025099 
iB32_240_v n1_20583_11663 0  0.025099 
iB32_240_g 0 n0_20491_11956  0.025099 
iB32_241_v n1_20583_11696 0  0.025099 
iB32_241_g 0 n0_20491_11956  0.025099 
iB32_242_v n1_20630_11663 0  0.025099 
iB32_242_g 0 n0_20679_11956  0.025099 
iB32_243_v n1_20630_11696 0  0.025099 
iB32_243_g 0 n0_20679_11956  0.025099 
iB32_244_v n1_20771_11447 0  0.025099 
iB32_244_g 0 n0_20679_11956  0.025099 
iB32_245_v n1_20771_11480 0  0.025099 
iB32_245_g 0 n0_20679_11956  0.025099 
iB32_246_v n1_20771_11663 0  0.025099 
iB32_246_g 0 n0_20679_11956  0.025099 
iB32_247_v n1_20771_11696 0  0.025099 
iB32_247_g 0 n0_20679_11956  0.025099 
iB32_248_v n1_20583_11879 0  0.025099 
iB32_248_g 0 n0_20491_11956  0.025099 
iB32_249_v n1_20583_11912 0  0.025099 
iB32_249_g 0 n0_20491_11956  0.025099 
iB32_250_v n1_20583_12095 0  0.025099 
iB32_250_g 0 n0_20491_12081  0.025099 
iB32_251_v n1_20583_12128 0  0.025099 
iB32_251_g 0 n0_20491_12114  0.025099 
iB32_252_v n1_20771_11879 0  0.025099 
iB32_252_g 0 n0_20679_11956  0.025099 
iB32_253_v n1_20771_11912 0  0.025099 
iB32_253_g 0 n0_20679_11956  0.025099 
iB32_254_v n1_20771_12095 0  0.025099 
iB32_254_g 0 n0_20679_12081  0.025099 
iB32_255_v n1_20771_12128 0  0.025099 
iB32_255_g 0 n0_20679_12114  0.025099 
iB32_256_v n1_20583_12311 0  0.025099 
iB32_256_g 0 n0_20491_12297  0.025099 
iB32_257_v n1_20583_12344 0  0.025099 
iB32_257_g 0 n0_20491_12330  0.025099 
iB32_258_v n1_20583_12527 0  0.025099 
iB32_258_g 0 n0_20491_12513  0.025099 
iB32_259_v n1_20583_12560 0  0.025099 
iB32_259_g 0 n0_20491_12546  0.025099 
iB32_260_v n1_20771_12311 0  0.025099 
iB32_260_g 0 n0_20679_12297  0.025099 
iB32_261_v n1_20771_12344 0  0.025099 
iB32_261_g 0 n0_20679_12330  0.025099 
iB32_262_v n1_20771_12527 0  0.025099 
iB32_262_g 0 n0_20679_12513  0.025099 
iB32_263_v n1_20771_12560 0  0.025099 
iB32_263_g 0 n0_20679_12546  0.025099 
iB32_264_v n1_20583_12743 0  0.025099 
iB32_264_g 0 n0_20491_12729  0.025099 
iB32_265_v n1_20583_12959 0  0.025099 
iB32_265_g 0 n0_20491_12945  0.025099 
iB32_266_v n1_20583_12992 0  0.025099 
iB32_266_g 0 n0_20491_12978  0.025099 
iB32_267_v n1_20771_12743 0  0.025099 
iB32_267_g 0 n0_20679_12729  0.025099 
iB32_268_v n1_20771_12776 0  0.025099 
iB32_268_g 0 n0_20679_12762  0.025099 
iB32_269_v n1_20771_12959 0  0.025099 
iB32_269_g 0 n0_20679_12945  0.025099 
iB32_270_v n1_20771_12992 0  0.025099 
iB32_270_g 0 n0_20679_12978  0.025099 
iB32_271_v n1_20583_13175 0  0.025099 
iB32_271_g 0 n0_20491_13161  0.025099 
iB32_272_v n1_20583_13208 0  0.025099 
iB32_272_g 0 n0_20491_13194  0.025099 
iB32_273_v n1_20583_13391 0  0.025099 
iB32_273_g 0 n0_20491_13377  0.025099 
iB32_274_v n1_20583_13424 0  0.025099 
iB32_274_g 0 n0_20491_13410  0.025099 
iB32_275_v n1_20771_13175 0  0.025099 
iB32_275_g 0 n0_20679_13161  0.025099 
iB32_276_v n1_20771_13208 0  0.025099 
iB32_276_g 0 n0_20679_13194  0.025099 
iB32_277_v n1_20771_13391 0  0.025099 
iB32_277_g 0 n0_20679_13377  0.025099 
iB32_278_v n1_20771_13424 0  0.025099 
iB32_278_g 0 n0_20679_13410  0.025099 
iB32_279_v n1_20583_13607 0  0.025099 
iB32_279_g 0 n0_20491_13593  0.025099 
iB32_280_v n1_20583_13640 0  0.025099 
iB32_280_g 0 n0_20491_13626  0.025099 
iB32_281_v n1_20583_13823 0  0.025099 
iB32_281_g 0 n0_20491_13809  0.025099 
iB32_282_v n1_20583_13856 0  0.025099 
iB32_282_g 0 n0_20491_13842  0.025099 
iB32_283_v n1_20771_13607 0  0.025099 
iB32_283_g 0 n0_20679_13593  0.025099 
iB32_284_v n1_20771_13640 0  0.025099 
iB32_284_g 0 n0_20679_13626  0.025099 
iB32_285_v n1_20771_13823 0  0.025099 
iB32_285_g 0 n0_20679_13809  0.025099 
iB32_286_v n1_20771_13856 0  0.025099 
iB32_286_g 0 n0_20679_13842  0.025099 
iB32_287_v n1_20583_14039 0  0.025099 
iB32_287_g 0 n0_20491_14025  0.025099 
iB32_288_v n1_20583_14072 0  0.025099 
iB32_288_g 0 n0_20491_14058  0.025099 
iB32_289_v n1_20583_14255 0  0.025099 
iB32_289_g 0 n0_20491_14241  0.025099 
iB32_290_v n1_20630_14039 0  0.025099 
iB32_290_g 0 n0_20491_14025  0.025099 
iB32_291_v n1_20771_14039 0  0.025099 
iB32_291_g 0 n0_20679_13842  0.025099 
iB32_292_v n1_20771_14072 0  0.025099 
iB32_292_g 0 n0_20679_14241  0.025099 
iB32_293_v n1_20771_14255 0  0.025099 
iB32_293_g 0 n0_20679_14241  0.025099 
iB32_294_v n1_20583_14288 0  0.025099 
iB32_294_g 0 n0_20491_14274  0.025099 
iB32_295_v n1_20583_14471 0  0.025099 
iB32_295_g 0 n0_20491_14457  0.025099 
iB32_296_v n1_20583_14504 0  0.025099 
iB32_296_g 0 n0_20491_14490  0.025099 
iB32_297_v n1_20771_14288 0  0.025099 
iB32_297_g 0 n0_20679_14274  0.025099 
iB32_298_v n1_20771_14471 0  0.025099 
iB32_298_g 0 n0_20679_14457  0.025099 
iB32_299_v n1_20771_14504 0  0.025099 
iB32_299_g 0 n0_20679_14490  0.025099 
iB32_300_v n1_20583_14687 0  0.025099 
iB32_300_g 0 n0_20491_14673  0.025099 
iB32_301_v n1_20583_14720 0  0.025099 
iB32_301_g 0 n0_20491_14706  0.025099 
iB32_302_v n1_20583_14903 0  0.025099 
iB32_302_g 0 n0_20491_14889  0.025099 
iB32_303_v n1_20583_14936 0  0.025099 
iB32_303_g 0 n0_20491_14936  0.025099 
iB32_304_v n1_20771_14687 0  0.025099 
iB32_304_g 0 n0_20679_14673  0.025099 
iB32_305_v n1_20771_14720 0  0.025099 
iB32_305_g 0 n0_20679_14706  0.025099 
iB32_306_v n1_20771_14903 0  0.025099 
iB32_306_g 0 n0_20679_14889  0.025099 
iB32_307_v n1_20771_14936 0  0.025099 
iB32_307_g 0 n0_20679_14936  0.025099 
iB32_308_v n1_20583_15308 0  0.025099 
iB32_308_g 0 n0_20491_15321  0.025099 
iB32_309_v n1_20583_15335 0  0.025099 
iB32_309_g 0 n0_20491_15321  0.025099 
iB32_310_v n1_20583_15368 0  0.025099 
iB32_310_g 0 n0_20491_15354  0.025099 
iB32_311_v n1_20771_15092 0  0.025099 
iB32_311_g 0 n0_20679_15105  0.025099 
iB32_312_v n1_20771_15119 0  0.025099 
iB32_312_g 0 n0_20679_15105  0.025099 
iB32_313_v n1_20771_15152 0  0.025099 
iB32_313_g 0 n0_20679_15152  0.025099 
iB32_314_v n1_20771_15308 0  0.025099 
iB32_314_g 0 n0_20679_15321  0.025099 
iB32_315_v n1_20771_15335 0  0.025099 
iB32_315_g 0 n0_20679_15321  0.025099 
iB32_316_v n1_20771_15368 0  0.025099 
iB32_316_g 0 n0_20679_15354  0.025099 
iB32_317_v n1_20583_15551 0  0.025099 
iB32_317_g 0 n0_20491_15537  0.025099 
iB32_318_v n1_20583_15584 0  0.025099 
iB32_318_g 0 n0_20491_15570  0.025099 
iB32_319_v n1_20583_15767 0  0.025099 
iB32_319_g 0 n0_20491_15753  0.025099 
iB32_320_v n1_20583_15800 0  0.025099 
iB32_320_g 0 n0_20491_15786  0.025099 
iB32_321_v n1_20771_15551 0  0.025099 
iB32_321_g 0 n0_20679_15537  0.025099 
iB32_322_v n1_20771_15584 0  0.025099 
iB32_322_g 0 n0_20679_15570  0.025099 
iB32_323_v n1_20771_15767 0  0.025099 
iB32_323_g 0 n0_20679_15753  0.025099 
iB32_324_v n1_20771_15800 0  0.025099 
iB32_324_g 0 n0_20679_15786  0.025099 
v189 _X_n3_7130_13971 0 1.8
v13f _X_n2_10505_9471 0 0
rrb4 n2_12755_2721 _X_n2_12755_2721 2.500000e-01
v201 _X_n3_20630_13971 0 1.8
v191 _X_n3_7130_11721 0 1.8
v9b _X_n2_7130_12846 0 0
rrb6 n2_12755_3846 _X_n2_12755_3846 2.500000e-01
v203 _X_n3_18380_13971 0 1.8
v193 _X_n3_9380_11721 0 1.8
v9d _X_n2_8255_12846 0 0
rr1a0 n3_7130_471 _X_n3_7130_471 2.500000e-01
rrb8 n2_12755_4971 _X_n2_12755_4971 2.500000e-01
v205 _X_n3_16130_13971 0 1.8
v195 _X_n3_380_471 0 1.8
v14b _X_n2_4880_8346 0 0
rrc0 n2_15005_1596 _X_n2_15005_1596 2.500000e-01
v9f _X_n2_380_10596 0 0
rr1a2 n3_7130_2721 _X_n3_7130_2721 2.500000e-01
v207 _X_n3_20630_16221 0 1.8
v197 _X_n3_2630_471 0 1.8
v14d _X_n2_6005_8346 0 0
rrc2 n2_15005_2721 _X_n2_15005_2721 2.500000e-01
rr1a4 n3_7130_4971 _X_n3_7130_4971 2.500000e-01
v209 _X_n3_18380_16221 0 1.8
v199 _X_n3_2630_2721 0 1.8
v14f _X_n2_7130_8346 0 0
rrc4 n2_15005_3846 _X_n2_15005_3846 2.500000e-01
v211 _X_n3_18380_18471 0 1.8
rr1a6 n3_7130_7221 _X_n3_7130_7221 2.500000e-01
rrc6 n2_15005_4971 _X_n2_15005_4971 2.500000e-01
v213 _X_n3_16130_20721 0 1.8
rr1a8 n3_9380_471 _X_n3_9380_471 2.500000e-01
rr1b0 n3_9380_9471 _X_n3_9380_9471 2.500000e-01
rrc8 n2_17255_471 _X_n2_17255_471 2.500000e-01
v215 _X_n3_16130_18471 0 1.8
v15b _X_n2_380_3846 0 0
rrd0 n2_20630_1596 _X_n2_20630_1596 2.500000e-01
rr1b2 n3_380_9471 _X_n3_380_9471 2.500000e-01
v217 _X_n3_16130_16221 0 1.8
v15d _X_n2_1505_3846 0 0
rrd2 n2_20630_3846 _X_n2_20630_3846 2.500000e-01
* vias from: 1 to 3
V24643 n1_333_383 n3_333_383 0.0
V24644 n1_333_431 n3_333_431 0.0
V24645 n1_333_464 n3_333_464 0.0
V24646 n1_333_647 n3_333_647 0.0
V24647 n1_333_680 n3_333_680 0.0
V24648 n1_333_863 n3_333_863 0.0
V24649 n1_333_896 n3_333_896 0.0
V24650 n1_333_1079 n3_333_1079 0.0
V24651 n1_333_1112 n3_333_1112 0.0
V24652 n1_333_1295 n3_333_1295 0.0
V24653 n1_333_1328 n3_333_1328 0.0
V24654 n1_333_1727 n3_333_1727 0.0
V24655 n1_333_1760 n3_333_1760 0.0
V24656 n1_333_1943 n3_333_1943 0.0
V24657 n1_333_1976 n3_333_1976 0.0
V24658 n1_333_2159 n3_333_2159 0.0
V24659 n1_333_2192 n3_333_2192 0.0
V24660 n1_333_2375 n3_333_2375 0.0
V24661 n1_333_2408 n3_333_2408 0.0
V24662 n1_333_2543 n3_333_2543 0.0
V24663 n1_333_2591 n3_333_2591 0.0
V24664 n1_333_2624 n3_333_2624 0.0
V24665 n1_333_2807 n3_333_2807 0.0
V24666 n1_333_2840 n3_333_2840 0.0
V24667 n1_333_3023 n3_333_3023 0.0
V24668 n1_333_3056 n3_333_3056 0.0
V24669 n1_333_3239 n3_333_3239 0.0
V24670 n1_333_3272 n3_333_3272 0.0
V24671 n1_333_3455 n3_333_3455 0.0
V24672 n1_333_3488 n3_333_3488 0.0
V24673 n1_333_3671 n3_333_3671 0.0
V24674 n1_333_3704 n3_333_3704 0.0
V24675 n1_333_4103 n3_333_4103 0.0
V24676 n1_333_4136 n3_333_4136 0.0
V24677 n1_333_4319 n3_333_4319 0.0
V24678 n1_333_4352 n3_333_4352 0.0
V24679 n1_333_4486 n3_333_4486 0.0
V24680 n1_333_4535 n3_333_4535 0.0
V24681 n1_333_4568 n3_333_4568 0.0
V24682 n1_333_4751 n3_333_4751 0.0
V24683 n1_333_4784 n3_333_4784 0.0
V24684 n1_333_4967 n3_333_4967 0.0
V24685 n1_333_5000 n3_333_5000 0.0
V24686 n1_333_5183 n3_333_5183 0.0
V24687 n1_333_5216 n3_333_5216 0.0
V24688 n1_333_5399 n3_333_5399 0.0
V24689 n1_333_5432 n3_333_5432 0.0
V24690 n1_333_5615 n3_333_5615 0.0
V24691 n1_333_5648 n3_333_5648 0.0
V24692 n1_333_5831 n3_333_5831 0.0
V24693 n1_333_5864 n3_333_5864 0.0
V24694 n1_333_6263 n3_333_6263 0.0
V24695 n1_333_6296 n3_333_6296 0.0
V24696 n1_333_6479 n3_333_6479 0.0
V24697 n1_333_6512 n3_333_6512 0.0
V24698 n1_333_6695 n3_333_6695 0.0
V24699 n1_333_6728 n3_333_6728 0.0
V24700 n1_333_6911 n3_333_6911 0.0
V24701 n1_333_6944 n3_333_6944 0.0
V24702 n1_333_7127 n3_333_7127 0.0
V24703 n1_333_7160 n3_333_7160 0.0
V24704 n1_333_7343 n3_333_7343 0.0
V24705 n1_333_7376 n3_333_7376 0.0
V24706 n1_333_7559 n3_333_7559 0.0
V24707 n1_333_7592 n3_333_7592 0.0
V24708 n1_333_7775 n3_333_7775 0.0
V24709 n1_333_7808 n3_333_7808 0.0
V24710 n1_333_7991 n3_333_7991 0.0
V24711 n1_333_8024 n3_333_8024 0.0
V24712 n1_333_8207 n3_333_8207 0.0
V24713 n1_333_8240 n3_333_8240 0.0
V24714 n1_333_8456 n3_333_8456 0.0
V24715 n1_333_8639 n3_333_8639 0.0
V24716 n1_333_8672 n3_333_8672 0.0
V24717 n1_333_8855 n3_333_8855 0.0
V24718 n1_333_8888 n3_333_8888 0.0
V24719 n1_333_9071 n3_333_9071 0.0
V24720 n1_333_9104 n3_333_9104 0.0
V24721 n1_333_9287 n3_333_9287 0.0
V24722 n1_333_9320 n3_333_9320 0.0
V24723 n1_333_9503 n3_333_9503 0.0
V24724 n1_333_9536 n3_333_9536 0.0
V24725 n1_333_9719 n3_333_9719 0.0
V24726 n1_333_9752 n3_333_9752 0.0
V24727 n1_333_9935 n3_333_9935 0.0
V24728 n1_333_9968 n3_333_9968 0.0
V24729 n1_333_10151 n3_333_10151 0.0
V24730 n1_333_10184 n3_333_10184 0.0
V24731 n1_333_10367 n3_333_10367 0.0
V24732 n1_333_10400 n3_333_10400 0.0
V24733 n1_333_10799 n3_333_10799 0.0
V24734 n1_333_10832 n3_333_10832 0.0
V24735 n1_333_11015 n3_333_11015 0.0
V24736 n1_333_11048 n3_333_11048 0.0
V24737 n1_333_11231 n3_333_11231 0.0
V24738 n1_333_11264 n3_333_11264 0.0
V24739 n1_333_11447 n3_333_11447 0.0
V24740 n1_333_11480 n3_333_11480 0.0
V24741 n1_333_11663 n3_333_11663 0.0
V24742 n1_333_11696 n3_333_11696 0.0
V24743 n1_333_11879 n3_333_11879 0.0
V24744 n1_333_11912 n3_333_11912 0.0
V24745 n1_333_12095 n3_333_12095 0.0
V24746 n1_333_12128 n3_333_12128 0.0
V24747 n1_333_12311 n3_333_12311 0.0
V24748 n1_333_12344 n3_333_12344 0.0
V24749 n1_333_12527 n3_333_12527 0.0
V24750 n1_333_12560 n3_333_12560 0.0
V24751 n1_333_12743 n3_333_12743 0.0
V24752 n1_333_12959 n3_333_12959 0.0
V24753 n1_333_12992 n3_333_12992 0.0
V24754 n1_333_13175 n3_333_13175 0.0
V24755 n1_333_13208 n3_333_13208 0.0
V24756 n1_333_13391 n3_333_13391 0.0
V24757 n1_333_13424 n3_333_13424 0.0
V24758 n1_333_13607 n3_333_13607 0.0
V24759 n1_333_13640 n3_333_13640 0.0
V24760 n1_333_13774 n3_333_13774 0.0
V24761 n1_333_13823 n3_333_13823 0.0
V24762 n1_333_13856 n3_333_13856 0.0
V24763 n1_333_14039 n3_333_14039 0.0
V24764 n1_333_14072 n3_333_14072 0.0
V24765 n1_333_14255 n3_333_14255 0.0
V24766 n1_333_14288 n3_333_14288 0.0
V24767 n1_333_14471 n3_333_14471 0.0
V24768 n1_333_14504 n3_333_14504 0.0
V24769 n1_333_14687 n3_333_14687 0.0
V24770 n1_333_14720 n3_333_14720 0.0
V24771 n1_333_14903 n3_333_14903 0.0
V24772 n1_333_14936 n3_333_14936 0.0
V24773 n1_333_15335 n3_333_15335 0.0
V24774 n1_333_15368 n3_333_15368 0.0
V24775 n1_333_15551 n3_333_15551 0.0
V24776 n1_333_15584 n3_333_15584 0.0
V24777 n1_333_15767 n3_333_15767 0.0
V24778 n1_333_15800 n3_333_15800 0.0
V24779 n1_333_15983 n3_333_15983 0.0
V24780 n1_333_16016 n3_333_16016 0.0
V24781 n1_333_16199 n3_333_16199 0.0
V24782 n1_333_16232 n3_333_16232 0.0
V24783 n1_333_16415 n3_333_16415 0.0
V24784 n1_333_16448 n3_333_16448 0.0
V24785 n1_333_16631 n3_333_16631 0.0
V24786 n1_333_16664 n3_333_16664 0.0
V24787 n1_333_16847 n3_333_16847 0.0
V24788 n1_333_16880 n3_333_16880 0.0
V24789 n1_333_17063 n3_333_17063 0.0
V24790 n1_333_17096 n3_333_17096 0.0
V24791 n1_333_17495 n3_333_17495 0.0
V24792 n1_333_17528 n3_333_17528 0.0
V24793 n1_333_17711 n3_333_17711 0.0
V24794 n1_333_17744 n3_333_17744 0.0
V24795 n1_333_17927 n3_333_17927 0.0
V24796 n1_333_17960 n3_333_17960 0.0
V24797 n1_333_18116 n3_333_18116 0.0
V24798 n1_333_18143 n3_333_18143 0.0
V24799 n1_333_18176 n3_333_18176 0.0
V24800 n1_333_18359 n3_333_18359 0.0
V24801 n1_333_18392 n3_333_18392 0.0
V24802 n1_333_18527 n3_333_18527 0.0
V24803 n1_333_18575 n3_333_18575 0.0
V24804 n1_333_18608 n3_333_18608 0.0
V24805 n1_333_18791 n3_333_18791 0.0
V24806 n1_333_18824 n3_333_18824 0.0
V24807 n1_333_19007 n3_333_19007 0.0
V24808 n1_333_19040 n3_333_19040 0.0
V24809 n1_333_19196 n3_333_19196 0.0
V24810 n1_333_19223 n3_333_19223 0.0
V24811 n1_333_19256 n3_333_19256 0.0
V24812 n1_333_19412 n3_333_19412 0.0
V24813 n1_333_19439 n3_333_19439 0.0
V24814 n1_333_19472 n3_333_19472 0.0
V24815 n1_333_19871 n3_333_19871 0.0
V24816 n1_333_19904 n3_333_19904 0.0
V24817 n1_333_20087 n3_333_20087 0.0
V24818 n1_333_20120 n3_333_20120 0.0
V24819 n1_333_20303 n3_333_20303 0.0
V24820 n1_333_20336 n3_333_20336 0.0
V24821 n1_333_20519 n3_333_20519 0.0
V24822 n1_333_20552 n3_333_20552 0.0
V24823 n1_333_20687 n3_333_20687 0.0
V24824 n1_333_20735 n3_333_20735 0.0
V24825 n1_333_20768 n3_333_20768 0.0
V24826 n1_380_431 n3_380_431 0.0
V24827 n1_380_464 n3_380_464 0.0
V24828 n1_380_4967 n3_380_4967 0.0
V24829 n1_380_5000 n3_380_5000 0.0
V24830 n1_380_7160 n3_380_7160 0.0
V24831 n1_380_9503 n3_380_9503 0.0
V24832 n1_380_9536 n3_380_9536 0.0
V24833 n1_380_11663 n3_380_11663 0.0
V24834 n1_380_11696 n3_380_11696 0.0
V24835 n1_380_14039 n3_380_14039 0.0
V24836 n1_380_16199 n3_380_16199 0.0
V24837 n1_380_16232 n3_380_16232 0.0
V24838 n1_380_18392 n3_380_18392 0.0
V24839 n1_380_18527 n3_380_18527 0.0
V24840 n1_380_20687 n3_380_20687 0.0
V24841 n1_380_20735 n3_380_20735 0.0
V24842 n1_380_20768 n3_380_20768 0.0
V24843 n1_521_215 n3_521_215 0.0
V24844 n1_521_248 n3_521_248 0.0
V24845 n1_521_383 n3_521_383 0.0
V24846 n1_521_431 n3_521_431 0.0
V24847 n1_521_647 n3_521_647 0.0
V24848 n1_521_680 n3_521_680 0.0
V24849 n1_521_863 n3_521_863 0.0
V24850 n1_521_896 n3_521_896 0.0
V24851 n1_521_1079 n3_521_1079 0.0
V24852 n1_521_1112 n3_521_1112 0.0
V24853 n1_521_1295 n3_521_1295 0.0
V24854 n1_521_1328 n3_521_1328 0.0
V24855 n1_521_1511 n3_521_1511 0.0
V24856 n1_521_1544 n3_521_1544 0.0
V24857 n1_521_1727 n3_521_1727 0.0
V24858 n1_521_1760 n3_521_1760 0.0
V24859 n1_521_1943 n3_521_1943 0.0
V24860 n1_521_1976 n3_521_1976 0.0
V24861 n1_521_2159 n3_521_2159 0.0
V24862 n1_521_2192 n3_521_2192 0.0
V24863 n1_521_2375 n3_521_2375 0.0
V24864 n1_521_2408 n3_521_2408 0.0
V24865 n1_521_2543 n3_521_2543 0.0
V24866 n1_521_2591 n3_521_2591 0.0
V24867 n1_521_2624 n3_521_2624 0.0
V24868 n1_521_2807 n3_521_2807 0.0
V24869 n1_521_2840 n3_521_2840 0.0
V24870 n1_521_3023 n3_521_3023 0.0
V24871 n1_521_3056 n3_521_3056 0.0
V24872 n1_521_3239 n3_521_3239 0.0
V24873 n1_521_3272 n3_521_3272 0.0
V24874 n1_521_3455 n3_521_3455 0.0
V24875 n1_521_3488 n3_521_3488 0.0
V24876 n1_521_3671 n3_521_3671 0.0
V24877 n1_521_3704 n3_521_3704 0.0
V24878 n1_521_3887 n3_521_3887 0.0
V24879 n1_521_3920 n3_521_3920 0.0
V24880 n1_521_4103 n3_521_4103 0.0
V24881 n1_521_4136 n3_521_4136 0.0
V24882 n1_521_4319 n3_521_4319 0.0
V24883 n1_521_4352 n3_521_4352 0.0
V24884 n1_521_4486 n3_521_4486 0.0
V24885 n1_521_4535 n3_521_4535 0.0
V24886 n1_521_4568 n3_521_4568 0.0
V24887 n1_521_4751 n3_521_4751 0.0
V24888 n1_521_4784 n3_521_4784 0.0
V24889 n1_521_5000 n3_521_5000 0.0
V24890 n1_521_5183 n3_521_5183 0.0
V24891 n1_521_5216 n3_521_5216 0.0
V24892 n1_521_5399 n3_521_5399 0.0
V24893 n1_521_5432 n3_521_5432 0.0
V24894 n1_521_5615 n3_521_5615 0.0
V24895 n1_521_5648 n3_521_5648 0.0
V24896 n1_521_5831 n3_521_5831 0.0
V24897 n1_521_5864 n3_521_5864 0.0
V24898 n1_521_6047 n3_521_6047 0.0
V24899 n1_521_6080 n3_521_6080 0.0
V24900 n1_521_6263 n3_521_6263 0.0
V24901 n1_521_6296 n3_521_6296 0.0
V24902 n1_521_6479 n3_521_6479 0.0
V24903 n1_521_6512 n3_521_6512 0.0
V24904 n1_521_6695 n3_521_6695 0.0
V24905 n1_521_6728 n3_521_6728 0.0
V24906 n1_521_6911 n3_521_6911 0.0
V24907 n1_521_6944 n3_521_6944 0.0
V24908 n1_521_7127 n3_521_7127 0.0
V24909 n1_521_7160 n3_521_7160 0.0
V24910 n1_521_7343 n3_521_7343 0.0
V24911 n1_521_7376 n3_521_7376 0.0
V24912 n1_521_7559 n3_521_7559 0.0
V24913 n1_521_7592 n3_521_7592 0.0
V24914 n1_521_7775 n3_521_7775 0.0
V24915 n1_521_7808 n3_521_7808 0.0
V24916 n1_521_7991 n3_521_7991 0.0
V24917 n1_521_8024 n3_521_8024 0.0
V24918 n1_521_8207 n3_521_8207 0.0
V24919 n1_521_8240 n3_521_8240 0.0
V24920 n1_521_8423 n3_521_8423 0.0
V24921 n1_521_8456 n3_521_8456 0.0
V24922 n1_521_8639 n3_521_8639 0.0
V24923 n1_521_8672 n3_521_8672 0.0
V24924 n1_521_8855 n3_521_8855 0.0
V24925 n1_521_8888 n3_521_8888 0.0
V24926 n1_521_9071 n3_521_9071 0.0
V24927 n1_521_9104 n3_521_9104 0.0
V24928 n1_521_9287 n3_521_9287 0.0
V24929 n1_521_9320 n3_521_9320 0.0
V24930 n1_521_9503 n3_521_9503 0.0
V24931 n1_521_9536 n3_521_9536 0.0
V24932 n1_521_9719 n3_521_9719 0.0
V24933 n1_521_9752 n3_521_9752 0.0
V24934 n1_521_9935 n3_521_9935 0.0
V24935 n1_521_9968 n3_521_9968 0.0
V24936 n1_521_10151 n3_521_10151 0.0
V24937 n1_521_10184 n3_521_10184 0.0
V24938 n1_521_10367 n3_521_10367 0.0
V24939 n1_521_10400 n3_521_10400 0.0
V24940 n1_521_10616 n3_521_10616 0.0
V24941 n1_521_10799 n3_521_10799 0.0
V24942 n1_521_10832 n3_521_10832 0.0
V24943 n1_521_11015 n3_521_11015 0.0
V24944 n1_521_11048 n3_521_11048 0.0
V24945 n1_521_11231 n3_521_11231 0.0
V24946 n1_521_11264 n3_521_11264 0.0
V24947 n1_521_11447 n3_521_11447 0.0
V24948 n1_521_11480 n3_521_11480 0.0
V24949 n1_521_11663 n3_521_11663 0.0
V24950 n1_521_11696 n3_521_11696 0.0
V24951 n1_521_11879 n3_521_11879 0.0
V24952 n1_521_11912 n3_521_11912 0.0
V24953 n1_521_12095 n3_521_12095 0.0
V24954 n1_521_12128 n3_521_12128 0.0
V24955 n1_521_12311 n3_521_12311 0.0
V24956 n1_521_12344 n3_521_12344 0.0
V24957 n1_521_12527 n3_521_12527 0.0
V24958 n1_521_12560 n3_521_12560 0.0
V24959 n1_521_12743 n3_521_12743 0.0
V24960 n1_521_12776 n3_521_12776 0.0
V24961 n1_521_12959 n3_521_12959 0.0
V24962 n1_521_12992 n3_521_12992 0.0
V24963 n1_521_13175 n3_521_13175 0.0
V24964 n1_521_13208 n3_521_13208 0.0
V24965 n1_521_13391 n3_521_13391 0.0
V24966 n1_521_13424 n3_521_13424 0.0
V24967 n1_521_13607 n3_521_13607 0.0
V24968 n1_521_13640 n3_521_13640 0.0
V24969 n1_521_13774 n3_521_13774 0.0
V24970 n1_521_13823 n3_521_13823 0.0
V24971 n1_521_13856 n3_521_13856 0.0
V24972 n1_521_14039 n3_521_14039 0.0
V24973 n1_521_14072 n3_521_14072 0.0
V24974 n1_521_14255 n3_521_14255 0.0
V24975 n1_521_14288 n3_521_14288 0.0
V24976 n1_521_14471 n3_521_14471 0.0
V24977 n1_521_14504 n3_521_14504 0.0
V24978 n1_521_14687 n3_521_14687 0.0
V24979 n1_521_14720 n3_521_14720 0.0
V24980 n1_521_14903 n3_521_14903 0.0
V24981 n1_521_14936 n3_521_14936 0.0
V24982 n1_521_15119 n3_521_15119 0.0
V24983 n1_521_15152 n3_521_15152 0.0
V24984 n1_521_15335 n3_521_15335 0.0
V24985 n1_521_15368 n3_521_15368 0.0
V24986 n1_521_15551 n3_521_15551 0.0
V24987 n1_521_15584 n3_521_15584 0.0
V24988 n1_521_15767 n3_521_15767 0.0
V24989 n1_521_15800 n3_521_15800 0.0
V24990 n1_521_15983 n3_521_15983 0.0
V24991 n1_521_16016 n3_521_16016 0.0
V24992 n1_521_16199 n3_521_16199 0.0
V24993 n1_521_16415 n3_521_16415 0.0
V24994 n1_521_16448 n3_521_16448 0.0
V24995 n1_521_16631 n3_521_16631 0.0
V24996 n1_521_16664 n3_521_16664 0.0
V24997 n1_521_16847 n3_521_16847 0.0
V24998 n1_521_16880 n3_521_16880 0.0
V24999 n1_521_17063 n3_521_17063 0.0
V25000 n1_521_17096 n3_521_17096 0.0
V25001 n1_521_17279 n3_521_17279 0.0
V25002 n1_521_17312 n3_521_17312 0.0
V25003 n1_521_17495 n3_521_17495 0.0
V25004 n1_521_17528 n3_521_17528 0.0
V25005 n1_521_17711 n3_521_17711 0.0
V25006 n1_521_17744 n3_521_17744 0.0
V25007 n1_521_17927 n3_521_17927 0.0
V25008 n1_521_17960 n3_521_17960 0.0
V25009 n1_521_18116 n3_521_18116 0.0
V25010 n1_521_18143 n3_521_18143 0.0
V25011 n1_521_18176 n3_521_18176 0.0
V25012 n1_521_18359 n3_521_18359 0.0
V25013 n1_521_18392 n3_521_18392 0.0
V25014 n1_521_18527 n3_521_18527 0.0
V25015 n1_521_18575 n3_521_18575 0.0
V25016 n1_521_18608 n3_521_18608 0.0
V25017 n1_521_18791 n3_521_18791 0.0
V25018 n1_521_18824 n3_521_18824 0.0
V25019 n1_521_19007 n3_521_19007 0.0
V25020 n1_521_19040 n3_521_19040 0.0
V25021 n1_521_19196 n3_521_19196 0.0
V25022 n1_521_19223 n3_521_19223 0.0
V25023 n1_521_19256 n3_521_19256 0.0
V25024 n1_521_19412 n3_521_19412 0.0
V25025 n1_521_19439 n3_521_19439 0.0
V25026 n1_521_19472 n3_521_19472 0.0
V25027 n1_521_19655 n3_521_19655 0.0
V25028 n1_521_19688 n3_521_19688 0.0
V25029 n1_521_19871 n3_521_19871 0.0
V25030 n1_521_19904 n3_521_19904 0.0
V25031 n1_521_20087 n3_521_20087 0.0
V25032 n1_521_20120 n3_521_20120 0.0
V25033 n1_521_20303 n3_521_20303 0.0
V25034 n1_521_20336 n3_521_20336 0.0
V25035 n1_521_20519 n3_521_20519 0.0
V25036 n1_521_20552 n3_521_20552 0.0
V25037 n1_521_20687 n3_521_20687 0.0
V25038 n1_521_20768 n3_521_20768 0.0
V25039 n1_521_20951 n3_521_20951 0.0
V25040 n1_521_20984 n3_521_20984 0.0
V25041 n1_2400_215 n3_2400_215 0.0
V25042 n1_2400_248 n3_2400_248 0.0
V25043 n1_2400_383 n3_2400_383 0.0
V25044 n1_2400_431 n3_2400_431 0.0
V25045 n1_2400_464 n3_2400_464 0.0
V25046 n1_2400_647 n3_2400_647 0.0
V25047 n1_2400_680 n3_2400_680 0.0
V25048 n1_2400_863 n3_2400_863 0.0
V25049 n1_2400_896 n3_2400_896 0.0
V25050 n1_2400_1079 n3_2400_1079 0.0
V25051 n1_2400_1112 n3_2400_1112 0.0
V25052 n1_2400_1295 n3_2400_1295 0.0
V25053 n1_2400_1328 n3_2400_1328 0.0
V25054 n1_2400_1511 n3_2400_1511 0.0
V25055 n1_2400_1544 n3_2400_1544 0.0
V25056 n1_2400_1727 n3_2400_1727 0.0
V25057 n1_2400_1760 n3_2400_1760 0.0
V25058 n1_2400_1943 n3_2400_1943 0.0
V25059 n1_2400_1976 n3_2400_1976 0.0
V25060 n1_2400_2159 n3_2400_2159 0.0
V25061 n1_2400_2192 n3_2400_2192 0.0
V25062 n1_2400_2375 n3_2400_2375 0.0
V25063 n1_2400_2408 n3_2400_2408 0.0
V25064 n1_2400_2543 n3_2400_2543 0.0
V25065 n1_2400_2591 n3_2400_2591 0.0
V25066 n1_2400_2624 n3_2400_2624 0.0
V25067 n1_2400_18527 n3_2400_18527 0.0
V25068 n1_2400_18575 n3_2400_18575 0.0
V25069 n1_2400_18608 n3_2400_18608 0.0
V25070 n1_2400_18791 n3_2400_18791 0.0
V25071 n1_2400_18824 n3_2400_18824 0.0
V25072 n1_2400_19007 n3_2400_19007 0.0
V25073 n1_2400_19040 n3_2400_19040 0.0
V25074 n1_2400_19223 n3_2400_19223 0.0
V25075 n1_2400_19256 n3_2400_19256 0.0
V25076 n1_2400_19439 n3_2400_19439 0.0
V25077 n1_2400_19472 n3_2400_19472 0.0
V25078 n1_2400_19655 n3_2400_19655 0.0
V25079 n1_2400_19688 n3_2400_19688 0.0
V25080 n1_2400_19871 n3_2400_19871 0.0
V25081 n1_2400_19904 n3_2400_19904 0.0
V25082 n1_2400_20087 n3_2400_20087 0.0
V25083 n1_2400_20120 n3_2400_20120 0.0
V25084 n1_2400_20303 n3_2400_20303 0.0
V25085 n1_2400_20336 n3_2400_20336 0.0
V25086 n1_2400_20519 n3_2400_20519 0.0
V25087 n1_2400_20552 n3_2400_20552 0.0
V25088 n1_2400_20687 n3_2400_20687 0.0
V25089 n1_2400_20735 n3_2400_20735 0.0
V25090 n1_2400_20768 n3_2400_20768 0.0
V25091 n1_2400_20951 n3_2400_20951 0.0
V25092 n1_2400_20984 n3_2400_20984 0.0
V25093 n1_2583_215 n3_2583_215 0.0
V25094 n1_2583_248 n3_2583_248 0.0
V25095 n1_2583_383 n3_2583_383 0.0
V25096 n1_2583_431 n3_2583_431 0.0
V25097 n1_2583_464 n3_2583_464 0.0
V25098 n1_2583_647 n3_2583_647 0.0
V25099 n1_2583_680 n3_2583_680 0.0
V25100 n1_2583_863 n3_2583_863 0.0
V25101 n1_2583_896 n3_2583_896 0.0
V25102 n1_2583_1079 n3_2583_1079 0.0
V25103 n1_2583_1112 n3_2583_1112 0.0
V25104 n1_2583_1295 n3_2583_1295 0.0
V25105 n1_2583_1328 n3_2583_1328 0.0
V25106 n1_2583_1727 n3_2583_1727 0.0
V25107 n1_2583_1760 n3_2583_1760 0.0
V25108 n1_2583_1943 n3_2583_1943 0.0
V25109 n1_2583_1976 n3_2583_1976 0.0
V25110 n1_2583_2159 n3_2583_2159 0.0
V25111 n1_2583_2192 n3_2583_2192 0.0
V25112 n1_2583_2375 n3_2583_2375 0.0
V25113 n1_2583_2408 n3_2583_2408 0.0
V25114 n1_2583_2543 n3_2583_2543 0.0
V25115 n1_2583_2591 n3_2583_2591 0.0
V25116 n1_2583_2624 n3_2583_2624 0.0
V25117 n1_2583_2807 n3_2583_2807 0.0
V25118 n1_2583_2840 n3_2583_2840 0.0
V25119 n1_2583_3023 n3_2583_3023 0.0
V25120 n1_2583_3056 n3_2583_3056 0.0
V25121 n1_2583_3239 n3_2583_3239 0.0
V25122 n1_2583_3272 n3_2583_3272 0.0
V25123 n1_2583_3428 n3_2583_3428 0.0
V25124 n1_2583_3455 n3_2583_3455 0.0
V25125 n1_2583_3488 n3_2583_3488 0.0
V25126 n1_2583_3671 n3_2583_3671 0.0
V25127 n1_2583_3704 n3_2583_3704 0.0
V25128 n1_2583_4076 n3_2583_4076 0.0
V25129 n1_2583_4103 n3_2583_4103 0.0
V25130 n1_2583_4136 n3_2583_4136 0.0
V25131 n1_2583_4270 n3_2583_4270 0.0
V25132 n1_2583_4319 n3_2583_4319 0.0
V25133 n1_2583_4352 n3_2583_4352 0.0
V25134 n1_2583_4508 n3_2583_4508 0.0
V25135 n1_2583_4535 n3_2583_4535 0.0
V25136 n1_2583_4568 n3_2583_4568 0.0
V25137 n1_2583_4751 n3_2583_4751 0.0
V25138 n1_2583_4784 n3_2583_4784 0.0
V25139 n1_2583_4967 n3_2583_4967 0.0
V25140 n1_2583_5000 n3_2583_5000 0.0
V25141 n1_2583_5183 n3_2583_5183 0.0
V25142 n1_2583_5216 n3_2583_5216 0.0
V25143 n1_2583_5399 n3_2583_5399 0.0
V25144 n1_2583_5432 n3_2583_5432 0.0
V25145 n1_2583_5446 n3_2583_5446 0.0
V25146 n1_2583_5588 n3_2583_5588 0.0
V25147 n1_2583_5615 n3_2583_5615 0.0
V25148 n1_2583_5648 n3_2583_5648 0.0
V25149 n1_2583_5831 n3_2583_5831 0.0
V25150 n1_2583_5864 n3_2583_5864 0.0
V25151 n1_2583_6263 n3_2583_6263 0.0
V25152 n1_2583_6296 n3_2583_6296 0.0
V25153 n1_2583_6479 n3_2583_6479 0.0
V25154 n1_2583_6512 n3_2583_6512 0.0
V25155 n1_2583_6549 n3_2583_6549 0.0
V25156 n1_2583_6646 n3_2583_6646 0.0
V25157 n1_2583_6695 n3_2583_6695 0.0
V25158 n1_2583_6728 n3_2583_6728 0.0
V25159 n1_2583_6911 n3_2583_6911 0.0
V25160 n1_2583_6944 n3_2583_6944 0.0
V25161 n1_2583_7127 n3_2583_7127 0.0
V25162 n1_2583_7160 n3_2583_7160 0.0
V25163 n1_2583_7343 n3_2583_7343 0.0
V25164 n1_2583_7376 n3_2583_7376 0.0
V25165 n1_2583_7559 n3_2583_7559 0.0
V25166 n1_2583_7592 n3_2583_7592 0.0
V25167 n1_2583_7775 n3_2583_7775 0.0
V25168 n1_2583_7808 n3_2583_7808 0.0
V25169 n1_2583_7822 n3_2583_7822 0.0
V25170 n1_2583_7964 n3_2583_7964 0.0
V25171 n1_2583_7991 n3_2583_7991 0.0
V25172 n1_2583_8024 n3_2583_8024 0.0
V25173 n1_2583_8207 n3_2583_8207 0.0
V25174 n1_2583_8240 n3_2583_8240 0.0
V25175 n1_2583_8456 n3_2583_8456 0.0
V25176 n1_2583_8639 n3_2583_8639 0.0
V25177 n1_2583_8672 n3_2583_8672 0.0
V25178 n1_2583_8855 n3_2583_8855 0.0
V25179 n1_2583_8888 n3_2583_8888 0.0
V25180 n1_2583_8902 n3_2583_8902 0.0
V25181 n1_2583_9022 n3_2583_9022 0.0
V25182 n1_2583_9044 n3_2583_9044 0.0
V25183 n1_2583_9071 n3_2583_9071 0.0
V25184 n1_2583_9104 n3_2583_9104 0.0
V25185 n1_2583_9287 n3_2583_9287 0.0
V25186 n1_2583_9320 n3_2583_9320 0.0
V25187 n1_2583_9503 n3_2583_9503 0.0
V25188 n1_2583_9536 n3_2583_9536 0.0
V25189 n1_2583_9719 n3_2583_9719 0.0
V25190 n1_2583_9752 n3_2583_9752 0.0
V25191 n1_2583_9935 n3_2583_9935 0.0
V25192 n1_2583_9968 n3_2583_9968 0.0
V25193 n1_2583_9982 n3_2583_9982 0.0
V25194 n1_2583_10124 n3_2583_10124 0.0
V25195 n1_2583_10151 n3_2583_10151 0.0
V25196 n1_2583_10184 n3_2583_10184 0.0
V25197 n1_2583_10367 n3_2583_10367 0.0
V25198 n1_2583_10400 n3_2583_10400 0.0
V25199 n1_2583_10799 n3_2583_10799 0.0
V25200 n1_2583_10832 n3_2583_10832 0.0
V25201 n1_2583_11015 n3_2583_11015 0.0
V25202 n1_2583_11048 n3_2583_11048 0.0
V25203 n1_2583_11182 n3_2583_11182 0.0
V25204 n1_2583_11204 n3_2583_11204 0.0
V25205 n1_2583_11231 n3_2583_11231 0.0
V25206 n1_2583_11264 n3_2583_11264 0.0
V25207 n1_2583_11447 n3_2583_11447 0.0
V25208 n1_2583_11480 n3_2583_11480 0.0
V25209 n1_2583_11663 n3_2583_11663 0.0
V25210 n1_2583_11696 n3_2583_11696 0.0
V25211 n1_2583_11879 n3_2583_11879 0.0
V25212 n1_2583_11912 n3_2583_11912 0.0
V25213 n1_2583_12095 n3_2583_12095 0.0
V25214 n1_2583_12128 n3_2583_12128 0.0
V25215 n1_2583_12262 n3_2583_12262 0.0
V25216 n1_2583_12284 n3_2583_12284 0.0
V25217 n1_2583_12311 n3_2583_12311 0.0
V25218 n1_2583_12344 n3_2583_12344 0.0
V25219 n1_2583_12527 n3_2583_12527 0.0
V25220 n1_2583_12560 n3_2583_12560 0.0
V25221 n1_2583_12743 n3_2583_12743 0.0
V25222 n1_2583_12959 n3_2583_12959 0.0
V25223 n1_2583_12992 n3_2583_12992 0.0
V25224 n1_2583_13175 n3_2583_13175 0.0
V25225 n1_2583_13208 n3_2583_13208 0.0
V25226 n1_2583_13391 n3_2583_13391 0.0
V25227 n1_2583_13424 n3_2583_13424 0.0
V25228 n1_2583_13558 n3_2583_13558 0.0
V25229 n1_2583_13580 n3_2583_13580 0.0
V25230 n1_2583_13607 n3_2583_13607 0.0
V25231 n1_2583_13640 n3_2583_13640 0.0
V25232 n1_2583_13796 n3_2583_13796 0.0
V25233 n1_2583_13823 n3_2583_13823 0.0
V25234 n1_2583_13856 n3_2583_13856 0.0
V25235 n1_2583_13990 n3_2583_13990 0.0
V25236 n1_2583_14039 n3_2583_14039 0.0
V25237 n1_2583_14072 n3_2583_14072 0.0
V25238 n1_2583_14206 n3_2583_14206 0.0
V25239 n1_2583_14255 n3_2583_14255 0.0
V25240 n1_2583_14288 n3_2583_14288 0.0
V25241 n1_2583_14471 n3_2583_14471 0.0
V25242 n1_2583_14504 n3_2583_14504 0.0
V25243 n1_2583_14660 n3_2583_14660 0.0
V25244 n1_2583_14687 n3_2583_14687 0.0
V25245 n1_2583_14720 n3_2583_14720 0.0
V25246 n1_2583_14903 n3_2583_14903 0.0
V25247 n1_2583_14936 n3_2583_14936 0.0
V25248 n1_2583_15335 n3_2583_15335 0.0
V25249 n1_2583_15368 n3_2583_15368 0.0
V25250 n1_2583_15524 n3_2583_15524 0.0
V25251 n1_2583_15551 n3_2583_15551 0.0
V25252 n1_2583_15584 n3_2583_15584 0.0
V25253 n1_2583_15740 n3_2583_15740 0.0
V25254 n1_2583_15767 n3_2583_15767 0.0
V25255 n1_2583_15800 n3_2583_15800 0.0
V25256 n1_2583_15983 n3_2583_15983 0.0
V25257 n1_2583_16016 n3_2583_16016 0.0
V25258 n1_2583_16199 n3_2583_16199 0.0
V25259 n1_2583_16232 n3_2583_16232 0.0
V25260 n1_2583_16415 n3_2583_16415 0.0
V25261 n1_2583_16448 n3_2583_16448 0.0
V25262 n1_2583_16582 n3_2583_16582 0.0
V25263 n1_2583_16631 n3_2583_16631 0.0
V25264 n1_2583_16664 n3_2583_16664 0.0
V25265 n1_2583_16798 n3_2583_16798 0.0
V25266 n1_2583_16820 n3_2583_16820 0.0
V25267 n1_2583_16847 n3_2583_16847 0.0
V25268 n1_2583_16880 n3_2583_16880 0.0
V25269 n1_2583_17036 n3_2583_17036 0.0
V25270 n1_2583_17063 n3_2583_17063 0.0
V25271 n1_2583_17096 n3_2583_17096 0.0
V25272 n1_2583_17495 n3_2583_17495 0.0
V25273 n1_2583_17528 n3_2583_17528 0.0
V25274 n1_2583_17662 n3_2583_17662 0.0
V25275 n1_2583_17684 n3_2583_17684 0.0
V25276 n1_2583_17711 n3_2583_17711 0.0
V25277 n1_2583_17744 n3_2583_17744 0.0
V25278 n1_2583_17927 n3_2583_17927 0.0
V25279 n1_2583_17960 n3_2583_17960 0.0
V25280 n1_2583_18143 n3_2583_18143 0.0
V25281 n1_2583_18176 n3_2583_18176 0.0
V25282 n1_2583_18359 n3_2583_18359 0.0
V25283 n1_2583_18392 n3_2583_18392 0.0
V25284 n1_2583_18527 n3_2583_18527 0.0
V25285 n1_2583_18575 n3_2583_18575 0.0
V25286 n1_2583_18608 n3_2583_18608 0.0
V25287 n1_2583_18791 n3_2583_18791 0.0
V25288 n1_2583_18824 n3_2583_18824 0.0
V25289 n1_2583_19007 n3_2583_19007 0.0
V25290 n1_2583_19040 n3_2583_19040 0.0
V25291 n1_2583_19223 n3_2583_19223 0.0
V25292 n1_2583_19256 n3_2583_19256 0.0
V25293 n1_2583_19439 n3_2583_19439 0.0
V25294 n1_2583_19472 n3_2583_19472 0.0
V25295 n1_2583_19871 n3_2583_19871 0.0
V25296 n1_2583_19904 n3_2583_19904 0.0
V25297 n1_2583_20087 n3_2583_20087 0.0
V25298 n1_2583_20120 n3_2583_20120 0.0
V25299 n1_2583_20303 n3_2583_20303 0.0
V25300 n1_2583_20336 n3_2583_20336 0.0
V25301 n1_2583_20519 n3_2583_20519 0.0
V25302 n1_2583_20552 n3_2583_20552 0.0
V25303 n1_2583_20687 n3_2583_20687 0.0
V25304 n1_2583_20735 n3_2583_20735 0.0
V25305 n1_2583_20768 n3_2583_20768 0.0
V25306 n1_2583_20951 n3_2583_20951 0.0
V25307 n1_2583_20984 n3_2583_20984 0.0
V25308 n1_2630_431 n3_2630_431 0.0
V25309 n1_2630_464 n3_2630_464 0.0
V25310 n1_2630_4967 n3_2630_4967 0.0
V25311 n1_2630_5000 n3_2630_5000 0.0
V25312 n1_2630_7160 n3_2630_7160 0.0
V25313 n1_2630_9503 n3_2630_9503 0.0
V25314 n1_2630_9536 n3_2630_9536 0.0
V25315 n1_2630_11663 n3_2630_11663 0.0
V25316 n1_2630_11696 n3_2630_11696 0.0
V25317 n1_2630_13990 n3_2630_13990 0.0
V25318 n1_2630_14039 n3_2630_14039 0.0
V25319 n1_2630_16199 n3_2630_16199 0.0
V25320 n1_2630_16232 n3_2630_16232 0.0
V25321 n1_2630_18392 n3_2630_18392 0.0
V25322 n1_2630_18527 n3_2630_18527 0.0
V25323 n1_2630_20687 n3_2630_20687 0.0
V25324 n1_2630_20735 n3_2630_20735 0.0
V25325 n1_2630_20768 n3_2630_20768 0.0
V25326 n1_2771_215 n3_2771_215 0.0
V25327 n1_2771_248 n3_2771_248 0.0
V25328 n1_2771_383 n3_2771_383 0.0
V25329 n1_2771_431 n3_2771_431 0.0
V25330 n1_2771_647 n3_2771_647 0.0
V25331 n1_2771_680 n3_2771_680 0.0
V25332 n1_2771_863 n3_2771_863 0.0
V25333 n1_2771_896 n3_2771_896 0.0
V25334 n1_2771_1079 n3_2771_1079 0.0
V25335 n1_2771_1112 n3_2771_1112 0.0
V25336 n1_2771_1295 n3_2771_1295 0.0
V25337 n1_2771_1328 n3_2771_1328 0.0
V25338 n1_2771_1511 n3_2771_1511 0.0
V25339 n1_2771_1544 n3_2771_1544 0.0
V25340 n1_2771_1727 n3_2771_1727 0.0
V25341 n1_2771_1760 n3_2771_1760 0.0
V25342 n1_2771_1943 n3_2771_1943 0.0
V25343 n1_2771_1976 n3_2771_1976 0.0
V25344 n1_2771_2159 n3_2771_2159 0.0
V25345 n1_2771_2192 n3_2771_2192 0.0
V25346 n1_2771_2375 n3_2771_2375 0.0
V25347 n1_2771_2408 n3_2771_2408 0.0
V25348 n1_2771_2543 n3_2771_2543 0.0
V25349 n1_2771_2591 n3_2771_2591 0.0
V25350 n1_2771_2624 n3_2771_2624 0.0
V25351 n1_2771_2807 n3_2771_2807 0.0
V25352 n1_2771_2840 n3_2771_2840 0.0
V25353 n1_2771_3023 n3_2771_3023 0.0
V25354 n1_2771_3056 n3_2771_3056 0.0
V25355 n1_2771_3239 n3_2771_3239 0.0
V25356 n1_2771_3272 n3_2771_3272 0.0
V25357 n1_2771_3428 n3_2771_3428 0.0
V25358 n1_2771_3455 n3_2771_3455 0.0
V25359 n1_2771_3488 n3_2771_3488 0.0
V25360 n1_2771_3671 n3_2771_3671 0.0
V25361 n1_2771_3704 n3_2771_3704 0.0
V25362 n1_2771_3860 n3_2771_3860 0.0
V25363 n1_2771_3887 n3_2771_3887 0.0
V25364 n1_2771_3920 n3_2771_3920 0.0
V25365 n1_2771_4076 n3_2771_4076 0.0
V25366 n1_2771_4103 n3_2771_4103 0.0
V25367 n1_2771_4136 n3_2771_4136 0.0
V25368 n1_2771_4270 n3_2771_4270 0.0
V25369 n1_2771_4319 n3_2771_4319 0.0
V25370 n1_2771_4352 n3_2771_4352 0.0
V25371 n1_2771_4508 n3_2771_4508 0.0
V25372 n1_2771_4535 n3_2771_4535 0.0
V25373 n1_2771_4568 n3_2771_4568 0.0
V25374 n1_2771_4751 n3_2771_4751 0.0
V25375 n1_2771_4784 n3_2771_4784 0.0
V25376 n1_2771_5000 n3_2771_5000 0.0
V25377 n1_2771_5183 n3_2771_5183 0.0
V25378 n1_2771_5216 n3_2771_5216 0.0
V25379 n1_2771_5399 n3_2771_5399 0.0
V25380 n1_2771_5432 n3_2771_5432 0.0
V25381 n1_2771_5446 n3_2771_5446 0.0
V25382 n1_2771_5588 n3_2771_5588 0.0
V25383 n1_2771_5615 n3_2771_5615 0.0
V25384 n1_2771_5648 n3_2771_5648 0.0
V25385 n1_2771_5831 n3_2771_5831 0.0
V25386 n1_2771_5864 n3_2771_5864 0.0
V25387 n1_2771_6047 n3_2771_6047 0.0
V25388 n1_2771_6080 n3_2771_6080 0.0
V25389 n1_2771_6263 n3_2771_6263 0.0
V25390 n1_2771_6296 n3_2771_6296 0.0
V25391 n1_2771_6479 n3_2771_6479 0.0
V25392 n1_2771_6512 n3_2771_6512 0.0
V25393 n1_2771_6549 n3_2771_6549 0.0
V25394 n1_2771_6646 n3_2771_6646 0.0
V25395 n1_2771_6695 n3_2771_6695 0.0
V25396 n1_2771_6728 n3_2771_6728 0.0
V25397 n1_2771_6911 n3_2771_6911 0.0
V25398 n1_2771_6944 n3_2771_6944 0.0
V25399 n1_2771_7127 n3_2771_7127 0.0
V25400 n1_2771_7160 n3_2771_7160 0.0
V25401 n1_2771_7343 n3_2771_7343 0.0
V25402 n1_2771_7376 n3_2771_7376 0.0
V25403 n1_2771_7559 n3_2771_7559 0.0
V25404 n1_2771_7592 n3_2771_7592 0.0
V25405 n1_2771_7775 n3_2771_7775 0.0
V25406 n1_2771_7808 n3_2771_7808 0.0
V25407 n1_2771_7822 n3_2771_7822 0.0
V25408 n1_2771_7964 n3_2771_7964 0.0
V25409 n1_2771_7991 n3_2771_7991 0.0
V25410 n1_2771_8024 n3_2771_8024 0.0
V25411 n1_2771_8207 n3_2771_8207 0.0
V25412 n1_2771_8240 n3_2771_8240 0.0
V25413 n1_2771_8423 n3_2771_8423 0.0
V25414 n1_2771_8456 n3_2771_8456 0.0
V25415 n1_2771_8639 n3_2771_8639 0.0
V25416 n1_2771_8672 n3_2771_8672 0.0
V25417 n1_2771_8855 n3_2771_8855 0.0
V25418 n1_2771_8888 n3_2771_8888 0.0
V25419 n1_2771_8902 n3_2771_8902 0.0
V25420 n1_2771_9022 n3_2771_9022 0.0
V25421 n1_2771_9044 n3_2771_9044 0.0
V25422 n1_2771_9071 n3_2771_9071 0.0
V25423 n1_2771_9104 n3_2771_9104 0.0
V25424 n1_2771_9287 n3_2771_9287 0.0
V25425 n1_2771_9320 n3_2771_9320 0.0
V25426 n1_2771_9503 n3_2771_9503 0.0
V25427 n1_2771_9536 n3_2771_9536 0.0
V25428 n1_2771_9719 n3_2771_9719 0.0
V25429 n1_2771_9752 n3_2771_9752 0.0
V25430 n1_2771_9935 n3_2771_9935 0.0
V25431 n1_2771_9968 n3_2771_9968 0.0
V25432 n1_2771_9982 n3_2771_9982 0.0
V25433 n1_2771_10124 n3_2771_10124 0.0
V25434 n1_2771_10151 n3_2771_10151 0.0
V25435 n1_2771_10184 n3_2771_10184 0.0
V25436 n1_2771_10367 n3_2771_10367 0.0
V25437 n1_2771_10400 n3_2771_10400 0.0
V25438 n1_2771_10616 n3_2771_10616 0.0
V25439 n1_2771_10799 n3_2771_10799 0.0
V25440 n1_2771_10832 n3_2771_10832 0.0
V25441 n1_2771_11015 n3_2771_11015 0.0
V25442 n1_2771_11048 n3_2771_11048 0.0
V25443 n1_2771_11182 n3_2771_11182 0.0
V25444 n1_2771_11204 n3_2771_11204 0.0
V25445 n1_2771_11231 n3_2771_11231 0.0
V25446 n1_2771_11264 n3_2771_11264 0.0
V25447 n1_2771_11447 n3_2771_11447 0.0
V25448 n1_2771_11480 n3_2771_11480 0.0
V25449 n1_2771_11663 n3_2771_11663 0.0
V25450 n1_2771_11696 n3_2771_11696 0.0
V25451 n1_2771_11879 n3_2771_11879 0.0
V25452 n1_2771_11912 n3_2771_11912 0.0
V25453 n1_2771_12095 n3_2771_12095 0.0
V25454 n1_2771_12128 n3_2771_12128 0.0
V25455 n1_2771_12262 n3_2771_12262 0.0
V25456 n1_2771_12284 n3_2771_12284 0.0
V25457 n1_2771_12311 n3_2771_12311 0.0
V25458 n1_2771_12344 n3_2771_12344 0.0
V25459 n1_2771_12527 n3_2771_12527 0.0
V25460 n1_2771_12560 n3_2771_12560 0.0
V25461 n1_2771_12743 n3_2771_12743 0.0
V25462 n1_2771_12776 n3_2771_12776 0.0
V25463 n1_2771_12959 n3_2771_12959 0.0
V25464 n1_2771_12992 n3_2771_12992 0.0
V25465 n1_2771_13175 n3_2771_13175 0.0
V25466 n1_2771_13208 n3_2771_13208 0.0
V25467 n1_2771_13391 n3_2771_13391 0.0
V25468 n1_2771_13424 n3_2771_13424 0.0
V25469 n1_2771_13558 n3_2771_13558 0.0
V25470 n1_2771_13580 n3_2771_13580 0.0
V25471 n1_2771_13607 n3_2771_13607 0.0
V25472 n1_2771_13640 n3_2771_13640 0.0
V25473 n1_2771_13796 n3_2771_13796 0.0
V25474 n1_2771_13823 n3_2771_13823 0.0
V25475 n1_2771_13856 n3_2771_13856 0.0
V25476 n1_2771_13990 n3_2771_13990 0.0
V25477 n1_2771_14039 n3_2771_14039 0.0
V25478 n1_2771_14072 n3_2771_14072 0.0
V25479 n1_2771_14206 n3_2771_14206 0.0
V25480 n1_2771_14255 n3_2771_14255 0.0
V25481 n1_2771_14288 n3_2771_14288 0.0
V25482 n1_2771_14471 n3_2771_14471 0.0
V25483 n1_2771_14504 n3_2771_14504 0.0
V25484 n1_2771_14660 n3_2771_14660 0.0
V25485 n1_2771_14687 n3_2771_14687 0.0
V25486 n1_2771_14720 n3_2771_14720 0.0
V25487 n1_2771_14903 n3_2771_14903 0.0
V25488 n1_2771_14936 n3_2771_14936 0.0
V25489 n1_2771_15119 n3_2771_15119 0.0
V25490 n1_2771_15152 n3_2771_15152 0.0
V25491 n1_2771_15335 n3_2771_15335 0.0
V25492 n1_2771_15368 n3_2771_15368 0.0
V25493 n1_2771_15524 n3_2771_15524 0.0
V25494 n1_2771_15551 n3_2771_15551 0.0
V25495 n1_2771_15584 n3_2771_15584 0.0
V25496 n1_2771_15740 n3_2771_15740 0.0
V25497 n1_2771_15767 n3_2771_15767 0.0
V25498 n1_2771_15800 n3_2771_15800 0.0
V25499 n1_2771_15983 n3_2771_15983 0.0
V25500 n1_2771_16016 n3_2771_16016 0.0
V25501 n1_2771_16199 n3_2771_16199 0.0
V25502 n1_2771_16415 n3_2771_16415 0.0
V25503 n1_2771_16448 n3_2771_16448 0.0
V25504 n1_2771_16582 n3_2771_16582 0.0
V25505 n1_2771_16631 n3_2771_16631 0.0
V25506 n1_2771_16664 n3_2771_16664 0.0
V25507 n1_2771_16798 n3_2771_16798 0.0
V25508 n1_2771_16820 n3_2771_16820 0.0
V25509 n1_2771_16847 n3_2771_16847 0.0
V25510 n1_2771_16880 n3_2771_16880 0.0
V25511 n1_2771_17036 n3_2771_17036 0.0
V25512 n1_2771_17063 n3_2771_17063 0.0
V25513 n1_2771_17096 n3_2771_17096 0.0
V25514 n1_2771_17279 n3_2771_17279 0.0
V25515 n1_2771_17312 n3_2771_17312 0.0
V25516 n1_2771_17495 n3_2771_17495 0.0
V25517 n1_2771_17528 n3_2771_17528 0.0
V25518 n1_2771_17662 n3_2771_17662 0.0
V25519 n1_2771_17684 n3_2771_17684 0.0
V25520 n1_2771_17711 n3_2771_17711 0.0
V25521 n1_2771_17744 n3_2771_17744 0.0
V25522 n1_2771_17927 n3_2771_17927 0.0
V25523 n1_2771_17960 n3_2771_17960 0.0
V25524 n1_2771_18143 n3_2771_18143 0.0
V25525 n1_2771_18176 n3_2771_18176 0.0
V25526 n1_2771_18359 n3_2771_18359 0.0
V25527 n1_2771_18392 n3_2771_18392 0.0
V25528 n1_2771_18527 n3_2771_18527 0.0
V25529 n1_2771_18575 n3_2771_18575 0.0
V25530 n1_2771_18608 n3_2771_18608 0.0
V25531 n1_2771_18791 n3_2771_18791 0.0
V25532 n1_2771_18824 n3_2771_18824 0.0
V25533 n1_2771_19007 n3_2771_19007 0.0
V25534 n1_2771_19040 n3_2771_19040 0.0
V25535 n1_2771_19223 n3_2771_19223 0.0
V25536 n1_2771_19256 n3_2771_19256 0.0
V25537 n1_2771_19439 n3_2771_19439 0.0
V25538 n1_2771_19472 n3_2771_19472 0.0
V25539 n1_2771_19655 n3_2771_19655 0.0
V25540 n1_2771_19688 n3_2771_19688 0.0
V25541 n1_2771_19871 n3_2771_19871 0.0
V25542 n1_2771_19904 n3_2771_19904 0.0
V25543 n1_2771_20087 n3_2771_20087 0.0
V25544 n1_2771_20120 n3_2771_20120 0.0
V25545 n1_2771_20303 n3_2771_20303 0.0
V25546 n1_2771_20336 n3_2771_20336 0.0
V25547 n1_2771_20519 n3_2771_20519 0.0
V25548 n1_2771_20552 n3_2771_20552 0.0
V25549 n1_2771_20687 n3_2771_20687 0.0
V25550 n1_2771_20768 n3_2771_20768 0.0
V25551 n1_2771_20951 n3_2771_20951 0.0
V25552 n1_2771_20984 n3_2771_20984 0.0
V25553 n1_2864_215 n3_2864_215 0.0
V25554 n1_2864_248 n3_2864_248 0.0
V25555 n1_2864_383 n3_2864_383 0.0
V25556 n1_2864_431 n3_2864_431 0.0
V25557 n1_2864_464 n3_2864_464 0.0
V25558 n1_2864_647 n3_2864_647 0.0
V25559 n1_2864_680 n3_2864_680 0.0
V25560 n1_2864_863 n3_2864_863 0.0
V25561 n1_2864_896 n3_2864_896 0.0
V25562 n1_2864_1079 n3_2864_1079 0.0
V25563 n1_2864_1112 n3_2864_1112 0.0
V25564 n1_2864_1295 n3_2864_1295 0.0
V25565 n1_2864_1328 n3_2864_1328 0.0
V25566 n1_2864_1511 n3_2864_1511 0.0
V25567 n1_2864_1544 n3_2864_1544 0.0
V25568 n1_2864_1727 n3_2864_1727 0.0
V25569 n1_2864_1760 n3_2864_1760 0.0
V25570 n1_2864_1943 n3_2864_1943 0.0
V25571 n1_2864_1976 n3_2864_1976 0.0
V25572 n1_2864_2159 n3_2864_2159 0.0
V25573 n1_2864_2192 n3_2864_2192 0.0
V25574 n1_2864_2375 n3_2864_2375 0.0
V25575 n1_2864_2408 n3_2864_2408 0.0
V25576 n1_2864_2543 n3_2864_2543 0.0
V25577 n1_2864_2591 n3_2864_2591 0.0
V25578 n1_2864_2624 n3_2864_2624 0.0
V25579 n1_2864_18527 n3_2864_18527 0.0
V25580 n1_2864_18575 n3_2864_18575 0.0
V25581 n1_2864_18608 n3_2864_18608 0.0
V25582 n1_2864_18791 n3_2864_18791 0.0
V25583 n1_2864_18824 n3_2864_18824 0.0
V25584 n1_2864_19007 n3_2864_19007 0.0
V25585 n1_2864_19040 n3_2864_19040 0.0
V25586 n1_2864_19223 n3_2864_19223 0.0
V25587 n1_2864_19256 n3_2864_19256 0.0
V25588 n1_2864_19439 n3_2864_19439 0.0
V25589 n1_2864_19472 n3_2864_19472 0.0
V25590 n1_2864_19655 n3_2864_19655 0.0
V25591 n1_2864_19688 n3_2864_19688 0.0
V25592 n1_2864_19871 n3_2864_19871 0.0
V25593 n1_2864_19904 n3_2864_19904 0.0
V25594 n1_2864_20087 n3_2864_20087 0.0
V25595 n1_2864_20120 n3_2864_20120 0.0
V25596 n1_2864_20303 n3_2864_20303 0.0
V25597 n1_2864_20336 n3_2864_20336 0.0
V25598 n1_2864_20519 n3_2864_20519 0.0
V25599 n1_2864_20552 n3_2864_20552 0.0
V25600 n1_2864_20687 n3_2864_20687 0.0
V25601 n1_2864_20735 n3_2864_20735 0.0
V25602 n1_2864_20768 n3_2864_20768 0.0
V25603 n1_2864_20951 n3_2864_20951 0.0
V25604 n1_2864_20984 n3_2864_20984 0.0
V25605 n1_4650_215 n3_4650_215 0.0
V25606 n1_4650_248 n3_4650_248 0.0
V25607 n1_4650_431 n3_4650_431 0.0
V25608 n1_4650_464 n3_4650_464 0.0
V25609 n1_4650_513 n3_4650_513 0.0
V25610 n1_4650_647 n3_4650_647 0.0
V25611 n1_4650_680 n3_4650_680 0.0
V25612 n1_4650_863 n3_4650_863 0.0
V25613 n1_4650_896 n3_4650_896 0.0
V25614 n1_4650_945 n3_4650_945 0.0
V25615 n1_4650_1079 n3_4650_1079 0.0
V25616 n1_4650_1112 n3_4650_1112 0.0
V25617 n1_4650_1295 n3_4650_1295 0.0
V25618 n1_4650_1328 n3_4650_1328 0.0
V25619 n1_4650_1511 n3_4650_1511 0.0
V25620 n1_4650_1544 n3_4650_1544 0.0
V25621 n1_4650_1727 n3_4650_1727 0.0
V25622 n1_4650_1760 n3_4650_1760 0.0
V25623 n1_4650_1943 n3_4650_1943 0.0
V25624 n1_4650_1976 n3_4650_1976 0.0
V25625 n1_4650_2132 n3_4650_2132 0.0
V25626 n1_4650_2159 n3_4650_2159 0.0
V25627 n1_4650_2192 n3_4650_2192 0.0
V25628 n1_4650_2375 n3_4650_2375 0.0
V25629 n1_4650_2408 n3_4650_2408 0.0
V25630 n1_4650_2543 n3_4650_2543 0.0
V25631 n1_4650_2591 n3_4650_2591 0.0
V25632 n1_4650_2624 n3_4650_2624 0.0
V25633 n1_4650_18527 n3_4650_18527 0.0
V25634 n1_4650_18575 n3_4650_18575 0.0
V25635 n1_4650_18608 n3_4650_18608 0.0
V25636 n1_4650_18791 n3_4650_18791 0.0
V25637 n1_4650_18824 n3_4650_18824 0.0
V25638 n1_4650_19007 n3_4650_19007 0.0
V25639 n1_4650_19040 n3_4650_19040 0.0
V25640 n1_4650_19223 n3_4650_19223 0.0
V25641 n1_4650_19256 n3_4650_19256 0.0
V25642 n1_4650_19439 n3_4650_19439 0.0
V25643 n1_4650_19472 n3_4650_19472 0.0
V25644 n1_4650_19655 n3_4650_19655 0.0
V25645 n1_4650_19688 n3_4650_19688 0.0
V25646 n1_4650_19871 n3_4650_19871 0.0
V25647 n1_4650_19904 n3_4650_19904 0.0
V25648 n1_4650_20087 n3_4650_20087 0.0
V25649 n1_4650_20120 n3_4650_20120 0.0
V25650 n1_4650_20303 n3_4650_20303 0.0
V25651 n1_4650_20336 n3_4650_20336 0.0
V25652 n1_4650_20519 n3_4650_20519 0.0
V25653 n1_4650_20552 n3_4650_20552 0.0
V25654 n1_4650_20687 n3_4650_20687 0.0
V25655 n1_4650_20735 n3_4650_20735 0.0
V25656 n1_4650_20768 n3_4650_20768 0.0
V25657 n1_4650_20951 n3_4650_20951 0.0
V25658 n1_4650_20984 n3_4650_20984 0.0
V25659 n1_4833_215 n3_4833_215 0.0
V25660 n1_4833_248 n3_4833_248 0.0
V25661 n1_4833_431 n3_4833_431 0.0
V25662 n1_4833_464 n3_4833_464 0.0
V25663 n1_4833_513 n3_4833_513 0.0
V25664 n1_4833_647 n3_4833_647 0.0
V25665 n1_4833_680 n3_4833_680 0.0
V25666 n1_4833_863 n3_4833_863 0.0
V25667 n1_4833_896 n3_4833_896 0.0
V25668 n1_4833_945 n3_4833_945 0.0
V25669 n1_4833_1079 n3_4833_1079 0.0
V25670 n1_4833_1112 n3_4833_1112 0.0
V25671 n1_4833_1295 n3_4833_1295 0.0
V25672 n1_4833_1328 n3_4833_1328 0.0
V25673 n1_4833_1727 n3_4833_1727 0.0
V25674 n1_4833_1760 n3_4833_1760 0.0
V25675 n1_4833_1916 n3_4833_1916 0.0
V25676 n1_4833_1943 n3_4833_1943 0.0
V25677 n1_4833_1976 n3_4833_1976 0.0
V25678 n1_4833_2132 n3_4833_2132 0.0
V25679 n1_4833_2159 n3_4833_2159 0.0
V25680 n1_4833_2192 n3_4833_2192 0.0
V25681 n1_4833_2375 n3_4833_2375 0.0
V25682 n1_4833_2408 n3_4833_2408 0.0
V25683 n1_4833_2543 n3_4833_2543 0.0
V25684 n1_4833_2564 n3_4833_2564 0.0
V25685 n1_4833_2591 n3_4833_2591 0.0
V25686 n1_4833_2624 n3_4833_2624 0.0
V25687 n1_4833_2807 n3_4833_2807 0.0
V25688 n1_4833_2840 n3_4833_2840 0.0
V25689 n1_4833_2996 n3_4833_2996 0.0
V25690 n1_4833_3023 n3_4833_3023 0.0
V25691 n1_4833_3056 n3_4833_3056 0.0
V25692 n1_4833_3212 n3_4833_3212 0.0
V25693 n1_4833_3239 n3_4833_3239 0.0
V25694 n1_4833_3272 n3_4833_3272 0.0
V25695 n1_4833_3455 n3_4833_3455 0.0
V25696 n1_4833_3488 n3_4833_3488 0.0
V25697 n1_4833_3644 n3_4833_3644 0.0
V25698 n1_4833_3671 n3_4833_3671 0.0
V25699 n1_4833_3704 n3_4833_3704 0.0
V25700 n1_4833_4103 n3_4833_4103 0.0
V25701 n1_4833_4136 n3_4833_4136 0.0
V25702 n1_4833_4292 n3_4833_4292 0.0
V25703 n1_4833_4319 n3_4833_4319 0.0
V25704 n1_4833_4352 n3_4833_4352 0.0
V25705 n1_4833_4486 n3_4833_4486 0.0
V25706 n1_4833_4508 n3_4833_4508 0.0
V25707 n1_4833_4535 n3_4833_4535 0.0
V25708 n1_4833_4568 n3_4833_4568 0.0
V25709 n1_4833_4751 n3_4833_4751 0.0
V25710 n1_4833_4784 n3_4833_4784 0.0
V25711 n1_4833_4967 n3_4833_4967 0.0
V25712 n1_4833_5000 n3_4833_5000 0.0
V25713 n1_4833_5183 n3_4833_5183 0.0
V25714 n1_4833_5216 n3_4833_5216 0.0
V25715 n1_4833_5399 n3_4833_5399 0.0
V25716 n1_4833_5432 n3_4833_5432 0.0
V25717 n1_4833_5446 n3_4833_5446 0.0
V25718 n1_4833_5588 n3_4833_5588 0.0
V25719 n1_4833_5615 n3_4833_5615 0.0
V25720 n1_4833_5648 n3_4833_5648 0.0
V25721 n1_4833_5831 n3_4833_5831 0.0
V25722 n1_4833_5864 n3_4833_5864 0.0
V25723 n1_4833_6263 n3_4833_6263 0.0
V25724 n1_4833_6296 n3_4833_6296 0.0
V25725 n1_4833_6479 n3_4833_6479 0.0
V25726 n1_4833_6512 n3_4833_6512 0.0
V25727 n1_4833_6549 n3_4833_6549 0.0
V25728 n1_4833_6646 n3_4833_6646 0.0
V25729 n1_4833_6695 n3_4833_6695 0.0
V25730 n1_4833_6728 n3_4833_6728 0.0
V25731 n1_4833_6911 n3_4833_6911 0.0
V25732 n1_4833_6944 n3_4833_6944 0.0
V25733 n1_4833_7127 n3_4833_7127 0.0
V25734 n1_4833_7160 n3_4833_7160 0.0
V25735 n1_4833_7343 n3_4833_7343 0.0
V25736 n1_4833_7376 n3_4833_7376 0.0
V25737 n1_4833_7559 n3_4833_7559 0.0
V25738 n1_4833_7592 n3_4833_7592 0.0
V25739 n1_4833_7775 n3_4833_7775 0.0
V25740 n1_4833_7808 n3_4833_7808 0.0
V25741 n1_4833_7822 n3_4833_7822 0.0
V25742 n1_4833_7964 n3_4833_7964 0.0
V25743 n1_4833_7991 n3_4833_7991 0.0
V25744 n1_4833_8024 n3_4833_8024 0.0
V25745 n1_4833_8207 n3_4833_8207 0.0
V25746 n1_4833_8240 n3_4833_8240 0.0
V25747 n1_4833_8456 n3_4833_8456 0.0
V25748 n1_4833_8639 n3_4833_8639 0.0
V25749 n1_4833_8672 n3_4833_8672 0.0
V25750 n1_4833_8855 n3_4833_8855 0.0
V25751 n1_4833_8888 n3_4833_8888 0.0
V25752 n1_4833_8902 n3_4833_8902 0.0
V25753 n1_4833_9022 n3_4833_9022 0.0
V25754 n1_4833_9044 n3_4833_9044 0.0
V25755 n1_4833_9071 n3_4833_9071 0.0
V25756 n1_4833_9104 n3_4833_9104 0.0
V25757 n1_4833_9287 n3_4833_9287 0.0
V25758 n1_4833_9320 n3_4833_9320 0.0
V25759 n1_4833_9503 n3_4833_9503 0.0
V25760 n1_4833_9536 n3_4833_9536 0.0
V25761 n1_4833_9719 n3_4833_9719 0.0
V25762 n1_4833_9752 n3_4833_9752 0.0
V25763 n1_4833_9935 n3_4833_9935 0.0
V25764 n1_4833_9968 n3_4833_9968 0.0
V25765 n1_4833_9982 n3_4833_9982 0.0
V25766 n1_4833_10124 n3_4833_10124 0.0
V25767 n1_4833_10151 n3_4833_10151 0.0
V25768 n1_4833_10184 n3_4833_10184 0.0
V25769 n1_4833_10367 n3_4833_10367 0.0
V25770 n1_4833_10400 n3_4833_10400 0.0
V25771 n1_4833_10799 n3_4833_10799 0.0
V25772 n1_4833_10832 n3_4833_10832 0.0
V25773 n1_4833_11015 n3_4833_11015 0.0
V25774 n1_4833_11048 n3_4833_11048 0.0
V25775 n1_4833_11182 n3_4833_11182 0.0
V25776 n1_4833_11204 n3_4833_11204 0.0
V25777 n1_4833_11231 n3_4833_11231 0.0
V25778 n1_4833_11264 n3_4833_11264 0.0
V25779 n1_4833_11447 n3_4833_11447 0.0
V25780 n1_4833_11480 n3_4833_11480 0.0
V25781 n1_4833_11663 n3_4833_11663 0.0
V25782 n1_4833_11696 n3_4833_11696 0.0
V25783 n1_4833_11879 n3_4833_11879 0.0
V25784 n1_4833_11912 n3_4833_11912 0.0
V25785 n1_4833_12095 n3_4833_12095 0.0
V25786 n1_4833_12128 n3_4833_12128 0.0
V25787 n1_4833_12284 n3_4833_12284 0.0
V25788 n1_4833_12311 n3_4833_12311 0.0
V25789 n1_4833_12344 n3_4833_12344 0.0
V25790 n1_4833_12527 n3_4833_12527 0.0
V25791 n1_4833_12560 n3_4833_12560 0.0
V25792 n1_4833_12743 n3_4833_12743 0.0
V25793 n1_4833_12959 n3_4833_12959 0.0
V25794 n1_4833_12992 n3_4833_12992 0.0
V25795 n1_4833_13175 n3_4833_13175 0.0
V25796 n1_4833_13208 n3_4833_13208 0.0
V25797 n1_4833_13391 n3_4833_13391 0.0
V25798 n1_4833_13424 n3_4833_13424 0.0
V25799 n1_4833_13580 n3_4833_13580 0.0
V25800 n1_4833_13607 n3_4833_13607 0.0
V25801 n1_4833_13640 n3_4833_13640 0.0
V25802 n1_4833_13823 n3_4833_13823 0.0
V25803 n1_4833_13856 n3_4833_13856 0.0
V25804 n1_4833_13990 n3_4833_13990 0.0
V25805 n1_4833_14039 n3_4833_14039 0.0
V25806 n1_4833_14072 n3_4833_14072 0.0
V25807 n1_4833_14206 n3_4833_14206 0.0
V25808 n1_4833_14255 n3_4833_14255 0.0
V25809 n1_4833_14288 n3_4833_14288 0.0
V25810 n1_4833_14471 n3_4833_14471 0.0
V25811 n1_4833_14504 n3_4833_14504 0.0
V25812 n1_4833_14687 n3_4833_14687 0.0
V25813 n1_4833_14720 n3_4833_14720 0.0
V25814 n1_4833_14903 n3_4833_14903 0.0
V25815 n1_4833_14936 n3_4833_14936 0.0
V25816 n1_4833_15335 n3_4833_15335 0.0
V25817 n1_4833_15368 n3_4833_15368 0.0
V25818 n1_4833_15524 n3_4833_15524 0.0
V25819 n1_4833_15551 n3_4833_15551 0.0
V25820 n1_4833_15584 n3_4833_15584 0.0
V25821 n1_4833_15740 n3_4833_15740 0.0
V25822 n1_4833_15767 n3_4833_15767 0.0
V25823 n1_4833_15800 n3_4833_15800 0.0
V25824 n1_4833_15983 n3_4833_15983 0.0
V25825 n1_4833_16016 n3_4833_16016 0.0
V25826 n1_4833_16172 n3_4833_16172 0.0
V25827 n1_4833_16199 n3_4833_16199 0.0
V25828 n1_4833_16232 n3_4833_16232 0.0
V25829 n1_4833_16415 n3_4833_16415 0.0
V25830 n1_4833_16448 n3_4833_16448 0.0
V25831 n1_4833_16631 n3_4833_16631 0.0
V25832 n1_4833_16664 n3_4833_16664 0.0
V25833 n1_4833_16847 n3_4833_16847 0.0
V25834 n1_4833_16880 n3_4833_16880 0.0
V25835 n1_4833_17036 n3_4833_17036 0.0
V25836 n1_4833_17063 n3_4833_17063 0.0
V25837 n1_4833_17096 n3_4833_17096 0.0
V25838 n1_4833_17468 n3_4833_17468 0.0
V25839 n1_4833_17495 n3_4833_17495 0.0
V25840 n1_4833_17528 n3_4833_17528 0.0
V25841 n1_4833_17684 n3_4833_17684 0.0
V25842 n1_4833_17711 n3_4833_17711 0.0
V25843 n1_4833_17744 n3_4833_17744 0.0
V25844 n1_4833_17927 n3_4833_17927 0.0
V25845 n1_4833_17960 n3_4833_17960 0.0
V25846 n1_4833_18143 n3_4833_18143 0.0
V25847 n1_4833_18176 n3_4833_18176 0.0
V25848 n1_4833_18359 n3_4833_18359 0.0
V25849 n1_4833_18392 n3_4833_18392 0.0
V25850 n1_4833_18527 n3_4833_18527 0.0
V25851 n1_4833_18548 n3_4833_18548 0.0
V25852 n1_4833_18575 n3_4833_18575 0.0
V25853 n1_4833_18608 n3_4833_18608 0.0
V25854 n1_4833_18764 n3_4833_18764 0.0
V25855 n1_4833_18791 n3_4833_18791 0.0
V25856 n1_4833_18824 n3_4833_18824 0.0
V25857 n1_4833_18980 n3_4833_18980 0.0
V25858 n1_4833_19007 n3_4833_19007 0.0
V25859 n1_4833_19040 n3_4833_19040 0.0
V25860 n1_4833_19196 n3_4833_19196 0.0
V25861 n1_4833_19223 n3_4833_19223 0.0
V25862 n1_4833_19256 n3_4833_19256 0.0
V25863 n1_4833_19439 n3_4833_19439 0.0
V25864 n1_4833_19472 n3_4833_19472 0.0
V25865 n1_4833_19871 n3_4833_19871 0.0
V25866 n1_4833_19904 n3_4833_19904 0.0
V25867 n1_4833_20087 n3_4833_20087 0.0
V25868 n1_4833_20120 n3_4833_20120 0.0
V25869 n1_4833_20303 n3_4833_20303 0.0
V25870 n1_4833_20336 n3_4833_20336 0.0
V25871 n1_4833_20519 n3_4833_20519 0.0
V25872 n1_4833_20552 n3_4833_20552 0.0
V25873 n1_4833_20687 n3_4833_20687 0.0
V25874 n1_4833_20735 n3_4833_20735 0.0
V25875 n1_4833_20768 n3_4833_20768 0.0
V25876 n1_4833_20951 n3_4833_20951 0.0
V25877 n1_4833_20984 n3_4833_20984 0.0
V25878 n1_4880_431 n3_4880_431 0.0
V25879 n1_4880_464 n3_4880_464 0.0
V25880 n1_4880_513 n3_4880_513 0.0
V25881 n1_4880_4967 n3_4880_4967 0.0
V25882 n1_4880_5000 n3_4880_5000 0.0
V25883 n1_4880_7160 n3_4880_7160 0.0
V25884 n1_4880_9503 n3_4880_9503 0.0
V25885 n1_4880_9536 n3_4880_9536 0.0
V25886 n1_4880_11663 n3_4880_11663 0.0
V25887 n1_4880_11696 n3_4880_11696 0.0
V25888 n1_4880_13990 n3_4880_13990 0.0
V25889 n1_4880_14039 n3_4880_14039 0.0
V25890 n1_4880_16172 n3_4880_16172 0.0
V25891 n1_4880_16199 n3_4880_16199 0.0
V25892 n1_4880_16232 n3_4880_16232 0.0
V25893 n1_4880_18392 n3_4880_18392 0.0
V25894 n1_4880_18527 n3_4880_18527 0.0
V25895 n1_4880_18548 n3_4880_18548 0.0
V25896 n1_4880_20687 n3_4880_20687 0.0
V25897 n1_4880_20735 n3_4880_20735 0.0
V25898 n1_4880_20768 n3_4880_20768 0.0
V25899 n1_5021_215 n3_5021_215 0.0
V25900 n1_5021_248 n3_5021_248 0.0
V25901 n1_5021_431 n3_5021_431 0.0
V25902 n1_5021_513 n3_5021_513 0.0
V25903 n1_5021_647 n3_5021_647 0.0
V25904 n1_5021_680 n3_5021_680 0.0
V25905 n1_5021_863 n3_5021_863 0.0
V25906 n1_5021_896 n3_5021_896 0.0
V25907 n1_5021_945 n3_5021_945 0.0
V25908 n1_5021_1079 n3_5021_1079 0.0
V25909 n1_5021_1112 n3_5021_1112 0.0
V25910 n1_5021_1295 n3_5021_1295 0.0
V25911 n1_5021_1328 n3_5021_1328 0.0
V25912 n1_5021_1511 n3_5021_1511 0.0
V25913 n1_5021_1544 n3_5021_1544 0.0
V25914 n1_5021_1727 n3_5021_1727 0.0
V25915 n1_5021_1760 n3_5021_1760 0.0
V25916 n1_5021_1916 n3_5021_1916 0.0
V25917 n1_5021_1943 n3_5021_1943 0.0
V25918 n1_5021_1976 n3_5021_1976 0.0
V25919 n1_5021_2132 n3_5021_2132 0.0
V25920 n1_5021_2159 n3_5021_2159 0.0
V25921 n1_5021_2192 n3_5021_2192 0.0
V25922 n1_5021_2375 n3_5021_2375 0.0
V25923 n1_5021_2408 n3_5021_2408 0.0
V25924 n1_5021_2543 n3_5021_2543 0.0
V25925 n1_5021_2564 n3_5021_2564 0.0
V25926 n1_5021_2591 n3_5021_2591 0.0
V25927 n1_5021_2624 n3_5021_2624 0.0
V25928 n1_5021_2807 n3_5021_2807 0.0
V25929 n1_5021_2840 n3_5021_2840 0.0
V25930 n1_5021_2996 n3_5021_2996 0.0
V25931 n1_5021_3023 n3_5021_3023 0.0
V25932 n1_5021_3056 n3_5021_3056 0.0
V25933 n1_5021_3212 n3_5021_3212 0.0
V25934 n1_5021_3239 n3_5021_3239 0.0
V25935 n1_5021_3272 n3_5021_3272 0.0
V25936 n1_5021_3455 n3_5021_3455 0.0
V25937 n1_5021_3488 n3_5021_3488 0.0
V25938 n1_5021_3644 n3_5021_3644 0.0
V25939 n1_5021_3671 n3_5021_3671 0.0
V25940 n1_5021_3704 n3_5021_3704 0.0
V25941 n1_5021_3887 n3_5021_3887 0.0
V25942 n1_5021_3920 n3_5021_3920 0.0
V25943 n1_5021_4103 n3_5021_4103 0.0
V25944 n1_5021_4136 n3_5021_4136 0.0
V25945 n1_5021_4292 n3_5021_4292 0.0
V25946 n1_5021_4319 n3_5021_4319 0.0
V25947 n1_5021_4352 n3_5021_4352 0.0
V25948 n1_5021_4486 n3_5021_4486 0.0
V25949 n1_5021_4508 n3_5021_4508 0.0
V25950 n1_5021_4535 n3_5021_4535 0.0
V25951 n1_5021_4568 n3_5021_4568 0.0
V25952 n1_5021_4751 n3_5021_4751 0.0
V25953 n1_5021_4784 n3_5021_4784 0.0
V25954 n1_5021_5000 n3_5021_5000 0.0
V25955 n1_5021_5183 n3_5021_5183 0.0
V25956 n1_5021_5216 n3_5021_5216 0.0
V25957 n1_5021_5399 n3_5021_5399 0.0
V25958 n1_5021_5432 n3_5021_5432 0.0
V25959 n1_5021_5446 n3_5021_5446 0.0
V25960 n1_5021_5588 n3_5021_5588 0.0
V25961 n1_5021_5615 n3_5021_5615 0.0
V25962 n1_5021_5648 n3_5021_5648 0.0
V25963 n1_5021_5831 n3_5021_5831 0.0
V25964 n1_5021_5864 n3_5021_5864 0.0
V25965 n1_5021_6047 n3_5021_6047 0.0
V25966 n1_5021_6080 n3_5021_6080 0.0
V25967 n1_5021_6263 n3_5021_6263 0.0
V25968 n1_5021_6296 n3_5021_6296 0.0
V25969 n1_5021_6479 n3_5021_6479 0.0
V25970 n1_5021_6512 n3_5021_6512 0.0
V25971 n1_5021_6549 n3_5021_6549 0.0
V25972 n1_5021_6646 n3_5021_6646 0.0
V25973 n1_5021_6695 n3_5021_6695 0.0
V25974 n1_5021_6728 n3_5021_6728 0.0
V25975 n1_5021_6911 n3_5021_6911 0.0
V25976 n1_5021_6944 n3_5021_6944 0.0
V25977 n1_5021_7127 n3_5021_7127 0.0
V25978 n1_5021_7160 n3_5021_7160 0.0
V25979 n1_5021_7343 n3_5021_7343 0.0
V25980 n1_5021_7376 n3_5021_7376 0.0
V25981 n1_5021_7559 n3_5021_7559 0.0
V25982 n1_5021_7592 n3_5021_7592 0.0
V25983 n1_5021_7775 n3_5021_7775 0.0
V25984 n1_5021_7808 n3_5021_7808 0.0
V25985 n1_5021_7822 n3_5021_7822 0.0
V25986 n1_5021_7964 n3_5021_7964 0.0
V25987 n1_5021_7991 n3_5021_7991 0.0
V25988 n1_5021_8024 n3_5021_8024 0.0
V25989 n1_5021_8207 n3_5021_8207 0.0
V25990 n1_5021_8240 n3_5021_8240 0.0
V25991 n1_5021_8423 n3_5021_8423 0.0
V25992 n1_5021_8456 n3_5021_8456 0.0
V25993 n1_5021_8639 n3_5021_8639 0.0
V25994 n1_5021_8672 n3_5021_8672 0.0
V25995 n1_5021_8855 n3_5021_8855 0.0
V25996 n1_5021_8888 n3_5021_8888 0.0
V25997 n1_5021_8902 n3_5021_8902 0.0
V25998 n1_5021_9022 n3_5021_9022 0.0
V25999 n1_5021_9044 n3_5021_9044 0.0
V26000 n1_5021_9071 n3_5021_9071 0.0
V26001 n1_5021_9104 n3_5021_9104 0.0
V26002 n1_5021_9287 n3_5021_9287 0.0
V26003 n1_5021_9320 n3_5021_9320 0.0
V26004 n1_5021_9503 n3_5021_9503 0.0
V26005 n1_5021_9536 n3_5021_9536 0.0
V26006 n1_5021_9719 n3_5021_9719 0.0
V26007 n1_5021_9752 n3_5021_9752 0.0
V26008 n1_5021_9935 n3_5021_9935 0.0
V26009 n1_5021_9968 n3_5021_9968 0.0
V26010 n1_5021_9982 n3_5021_9982 0.0
V26011 n1_5021_10124 n3_5021_10124 0.0
V26012 n1_5021_10151 n3_5021_10151 0.0
V26013 n1_5021_10184 n3_5021_10184 0.0
V26014 n1_5021_10367 n3_5021_10367 0.0
V26015 n1_5021_10400 n3_5021_10400 0.0
V26016 n1_5021_10616 n3_5021_10616 0.0
V26017 n1_5021_10799 n3_5021_10799 0.0
V26018 n1_5021_10832 n3_5021_10832 0.0
V26019 n1_5021_11015 n3_5021_11015 0.0
V26020 n1_5021_11048 n3_5021_11048 0.0
V26021 n1_5021_11182 n3_5021_11182 0.0
V26022 n1_5021_11204 n3_5021_11204 0.0
V26023 n1_5021_11231 n3_5021_11231 0.0
V26024 n1_5021_11264 n3_5021_11264 0.0
V26025 n1_5021_11447 n3_5021_11447 0.0
V26026 n1_5021_11480 n3_5021_11480 0.0
V26027 n1_5021_11663 n3_5021_11663 0.0
V26028 n1_5021_11696 n3_5021_11696 0.0
V26029 n1_5021_11879 n3_5021_11879 0.0
V26030 n1_5021_11912 n3_5021_11912 0.0
V26031 n1_5021_12095 n3_5021_12095 0.0
V26032 n1_5021_12128 n3_5021_12128 0.0
V26033 n1_5021_12284 n3_5021_12284 0.0
V26034 n1_5021_12311 n3_5021_12311 0.0
V26035 n1_5021_12344 n3_5021_12344 0.0
V26036 n1_5021_12527 n3_5021_12527 0.0
V26037 n1_5021_12560 n3_5021_12560 0.0
V26038 n1_5021_12743 n3_5021_12743 0.0
V26039 n1_5021_12776 n3_5021_12776 0.0
V26040 n1_5021_12959 n3_5021_12959 0.0
V26041 n1_5021_12992 n3_5021_12992 0.0
V26042 n1_5021_13175 n3_5021_13175 0.0
V26043 n1_5021_13208 n3_5021_13208 0.0
V26044 n1_5021_13391 n3_5021_13391 0.0
V26045 n1_5021_13424 n3_5021_13424 0.0
V26046 n1_5021_13580 n3_5021_13580 0.0
V26047 n1_5021_13607 n3_5021_13607 0.0
V26048 n1_5021_13640 n3_5021_13640 0.0
V26049 n1_5021_13823 n3_5021_13823 0.0
V26050 n1_5021_13856 n3_5021_13856 0.0
V26051 n1_5021_14039 n3_5021_14039 0.0
V26052 n1_5021_14072 n3_5021_14072 0.0
V26053 n1_5021_14206 n3_5021_14206 0.0
V26054 n1_5021_14255 n3_5021_14255 0.0
V26055 n1_5021_14288 n3_5021_14288 0.0
V26056 n1_5021_14471 n3_5021_14471 0.0
V26057 n1_5021_14504 n3_5021_14504 0.0
V26058 n1_5021_14687 n3_5021_14687 0.0
V26059 n1_5021_14720 n3_5021_14720 0.0
V26060 n1_5021_14903 n3_5021_14903 0.0
V26061 n1_5021_14936 n3_5021_14936 0.0
V26062 n1_5021_15119 n3_5021_15119 0.0
V26063 n1_5021_15152 n3_5021_15152 0.0
V26064 n1_5021_15335 n3_5021_15335 0.0
V26065 n1_5021_15368 n3_5021_15368 0.0
V26066 n1_5021_15524 n3_5021_15524 0.0
V26067 n1_5021_15551 n3_5021_15551 0.0
V26068 n1_5021_15584 n3_5021_15584 0.0
V26069 n1_5021_15740 n3_5021_15740 0.0
V26070 n1_5021_15767 n3_5021_15767 0.0
V26071 n1_5021_15800 n3_5021_15800 0.0
V26072 n1_5021_15983 n3_5021_15983 0.0
V26073 n1_5021_16016 n3_5021_16016 0.0
V26074 n1_5021_16172 n3_5021_16172 0.0
V26075 n1_5021_16199 n3_5021_16199 0.0
V26076 n1_5021_16415 n3_5021_16415 0.0
V26077 n1_5021_16448 n3_5021_16448 0.0
V26078 n1_5021_16631 n3_5021_16631 0.0
V26079 n1_5021_16664 n3_5021_16664 0.0
V26080 n1_5021_16847 n3_5021_16847 0.0
V26081 n1_5021_16880 n3_5021_16880 0.0
V26082 n1_5021_17036 n3_5021_17036 0.0
V26083 n1_5021_17063 n3_5021_17063 0.0
V26084 n1_5021_17096 n3_5021_17096 0.0
V26085 n1_5021_17252 n3_5021_17252 0.0
V26086 n1_5021_17279 n3_5021_17279 0.0
V26087 n1_5021_17312 n3_5021_17312 0.0
V26088 n1_5021_17446 n3_5021_17446 0.0
V26089 n1_5021_17468 n3_5021_17468 0.0
V26090 n1_5021_17495 n3_5021_17495 0.0
V26091 n1_5021_17528 n3_5021_17528 0.0
V26092 n1_5021_17684 n3_5021_17684 0.0
V26093 n1_5021_17711 n3_5021_17711 0.0
V26094 n1_5021_17744 n3_5021_17744 0.0
V26095 n1_5021_17927 n3_5021_17927 0.0
V26096 n1_5021_17960 n3_5021_17960 0.0
V26097 n1_5021_18143 n3_5021_18143 0.0
V26098 n1_5021_18176 n3_5021_18176 0.0
V26099 n1_5021_18359 n3_5021_18359 0.0
V26100 n1_5021_18392 n3_5021_18392 0.0
V26101 n1_5021_18527 n3_5021_18527 0.0
V26102 n1_5021_18548 n3_5021_18548 0.0
V26103 n1_5021_18575 n3_5021_18575 0.0
V26104 n1_5021_18608 n3_5021_18608 0.0
V26105 n1_5021_18764 n3_5021_18764 0.0
V26106 n1_5021_18791 n3_5021_18791 0.0
V26107 n1_5021_18824 n3_5021_18824 0.0
V26108 n1_5021_18980 n3_5021_18980 0.0
V26109 n1_5021_19007 n3_5021_19007 0.0
V26110 n1_5021_19040 n3_5021_19040 0.0
V26111 n1_5021_19196 n3_5021_19196 0.0
V26112 n1_5021_19223 n3_5021_19223 0.0
V26113 n1_5021_19256 n3_5021_19256 0.0
V26114 n1_5021_19439 n3_5021_19439 0.0
V26115 n1_5021_19472 n3_5021_19472 0.0
V26116 n1_5021_19628 n3_5021_19628 0.0
V26117 n1_5021_19655 n3_5021_19655 0.0
V26118 n1_5021_19688 n3_5021_19688 0.0
V26119 n1_5021_19871 n3_5021_19871 0.0
V26120 n1_5021_19904 n3_5021_19904 0.0
V26121 n1_5021_20087 n3_5021_20087 0.0
V26122 n1_5021_20120 n3_5021_20120 0.0
V26123 n1_5021_20303 n3_5021_20303 0.0
V26124 n1_5021_20336 n3_5021_20336 0.0
V26125 n1_5021_20519 n3_5021_20519 0.0
V26126 n1_5021_20552 n3_5021_20552 0.0
V26127 n1_5021_20687 n3_5021_20687 0.0
V26128 n1_5021_20768 n3_5021_20768 0.0
V26129 n1_5021_20951 n3_5021_20951 0.0
V26130 n1_5021_20984 n3_5021_20984 0.0
V26131 n1_5114_215 n3_5114_215 0.0
V26132 n1_5114_248 n3_5114_248 0.0
V26133 n1_5114_431 n3_5114_431 0.0
V26134 n1_5114_464 n3_5114_464 0.0
V26135 n1_5114_513 n3_5114_513 0.0
V26136 n1_5114_647 n3_5114_647 0.0
V26137 n1_5114_680 n3_5114_680 0.0
V26138 n1_5114_863 n3_5114_863 0.0
V26139 n1_5114_896 n3_5114_896 0.0
V26140 n1_5114_945 n3_5114_945 0.0
V26141 n1_5114_1079 n3_5114_1079 0.0
V26142 n1_5114_1112 n3_5114_1112 0.0
V26143 n1_5114_1295 n3_5114_1295 0.0
V26144 n1_5114_1328 n3_5114_1328 0.0
V26145 n1_5114_1511 n3_5114_1511 0.0
V26146 n1_5114_1544 n3_5114_1544 0.0
V26147 n1_5114_1727 n3_5114_1727 0.0
V26148 n1_5114_1760 n3_5114_1760 0.0
V26149 n1_5114_1916 n3_5114_1916 0.0
V26150 n1_5114_1943 n3_5114_1943 0.0
V26151 n1_5114_1976 n3_5114_1976 0.0
V26152 n1_5114_2159 n3_5114_2159 0.0
V26153 n1_5114_2192 n3_5114_2192 0.0
V26154 n1_5114_2375 n3_5114_2375 0.0
V26155 n1_5114_2408 n3_5114_2408 0.0
V26156 n1_5114_2543 n3_5114_2543 0.0
V26157 n1_5114_2564 n3_5114_2564 0.0
V26158 n1_5114_2591 n3_5114_2591 0.0
V26159 n1_5114_2624 n3_5114_2624 0.0
V26160 n1_5114_18527 n3_5114_18527 0.0
V26161 n1_5114_18548 n3_5114_18548 0.0
V26162 n1_5114_18575 n3_5114_18575 0.0
V26163 n1_5114_18608 n3_5114_18608 0.0
V26164 n1_5114_18764 n3_5114_18764 0.0
V26165 n1_5114_18791 n3_5114_18791 0.0
V26166 n1_5114_18824 n3_5114_18824 0.0
V26167 n1_5114_18980 n3_5114_18980 0.0
V26168 n1_5114_19007 n3_5114_19007 0.0
V26169 n1_5114_19040 n3_5114_19040 0.0
V26170 n1_5114_19196 n3_5114_19196 0.0
V26171 n1_5114_19223 n3_5114_19223 0.0
V26172 n1_5114_19256 n3_5114_19256 0.0
V26173 n1_5114_19439 n3_5114_19439 0.0
V26174 n1_5114_19472 n3_5114_19472 0.0
V26175 n1_5114_19628 n3_5114_19628 0.0
V26176 n1_5114_19655 n3_5114_19655 0.0
V26177 n1_5114_19688 n3_5114_19688 0.0
V26178 n1_5114_19871 n3_5114_19871 0.0
V26179 n1_5114_19904 n3_5114_19904 0.0
V26180 n1_5114_20087 n3_5114_20087 0.0
V26181 n1_5114_20120 n3_5114_20120 0.0
V26182 n1_5114_20303 n3_5114_20303 0.0
V26183 n1_5114_20336 n3_5114_20336 0.0
V26184 n1_5114_20519 n3_5114_20519 0.0
V26185 n1_5114_20552 n3_5114_20552 0.0
V26186 n1_5114_20687 n3_5114_20687 0.0
V26187 n1_5114_20735 n3_5114_20735 0.0
V26188 n1_5114_20768 n3_5114_20768 0.0
V26189 n1_5114_20951 n3_5114_20951 0.0
V26190 n1_5114_20984 n3_5114_20984 0.0
V26191 n1_6900_215 n3_6900_215 0.0
V26192 n1_6900_248 n3_6900_248 0.0
V26193 n1_6900_383 n3_6900_383 0.0
V26194 n1_6900_431 n3_6900_431 0.0
V26195 n1_6900_464 n3_6900_464 0.0
V26196 n1_6900_647 n3_6900_647 0.0
V26197 n1_6900_680 n3_6900_680 0.0
V26198 n1_6900_863 n3_6900_863 0.0
V26199 n1_6900_896 n3_6900_896 0.0
V26200 n1_6900_1079 n3_6900_1079 0.0
V26201 n1_6900_1112 n3_6900_1112 0.0
V26202 n1_6900_1295 n3_6900_1295 0.0
V26203 n1_6900_1328 n3_6900_1328 0.0
V26204 n1_6900_1511 n3_6900_1511 0.0
V26205 n1_6900_1544 n3_6900_1544 0.0
V26206 n1_6900_1727 n3_6900_1727 0.0
V26207 n1_6900_1760 n3_6900_1760 0.0
V26208 n1_6900_1916 n3_6900_1916 0.0
V26209 n1_6900_1943 n3_6900_1943 0.0
V26210 n1_6900_1976 n3_6900_1976 0.0
V26211 n1_6900_2159 n3_6900_2159 0.0
V26212 n1_6900_2192 n3_6900_2192 0.0
V26213 n1_6900_2375 n3_6900_2375 0.0
V26214 n1_6900_2408 n3_6900_2408 0.0
V26215 n1_6900_2543 n3_6900_2543 0.0
V26216 n1_6900_2564 n3_6900_2564 0.0
V26217 n1_6900_2591 n3_6900_2591 0.0
V26218 n1_6900_2624 n3_6900_2624 0.0
V26219 n1_6900_18527 n3_6900_18527 0.0
V26220 n1_6900_18548 n3_6900_18548 0.0
V26221 n1_6900_18575 n3_6900_18575 0.0
V26222 n1_6900_18608 n3_6900_18608 0.0
V26223 n1_6900_18764 n3_6900_18764 0.0
V26224 n1_6900_18791 n3_6900_18791 0.0
V26225 n1_6900_18824 n3_6900_18824 0.0
V26226 n1_6900_19007 n3_6900_19007 0.0
V26227 n1_6900_19040 n3_6900_19040 0.0
V26228 n1_6900_19196 n3_6900_19196 0.0
V26229 n1_6900_19223 n3_6900_19223 0.0
V26230 n1_6900_19256 n3_6900_19256 0.0
V26231 n1_6900_19439 n3_6900_19439 0.0
V26232 n1_6900_19472 n3_6900_19472 0.0
V26233 n1_6900_19655 n3_6900_19655 0.0
V26234 n1_6900_19688 n3_6900_19688 0.0
V26235 n1_6900_19871 n3_6900_19871 0.0
V26236 n1_6900_19904 n3_6900_19904 0.0
V26237 n1_6900_20087 n3_6900_20087 0.0
V26238 n1_6900_20120 n3_6900_20120 0.0
V26239 n1_6900_20303 n3_6900_20303 0.0
V26240 n1_6900_20336 n3_6900_20336 0.0
V26241 n1_6900_20519 n3_6900_20519 0.0
V26242 n1_6900_20552 n3_6900_20552 0.0
V26243 n1_6900_20687 n3_6900_20687 0.0
V26244 n1_6900_20735 n3_6900_20735 0.0
V26245 n1_6900_20768 n3_6900_20768 0.0
V26246 n1_6900_20951 n3_6900_20951 0.0
V26247 n1_6900_20984 n3_6900_20984 0.0
V26248 n1_7083_215 n3_7083_215 0.0
V26249 n1_7083_248 n3_7083_248 0.0
V26250 n1_7083_383 n3_7083_383 0.0
V26251 n1_7083_431 n3_7083_431 0.0
V26252 n1_7083_464 n3_7083_464 0.0
V26253 n1_7083_647 n3_7083_647 0.0
V26254 n1_7083_680 n3_7083_680 0.0
V26255 n1_7083_863 n3_7083_863 0.0
V26256 n1_7083_896 n3_7083_896 0.0
V26257 n1_7083_1079 n3_7083_1079 0.0
V26258 n1_7083_1112 n3_7083_1112 0.0
V26259 n1_7083_1295 n3_7083_1295 0.0
V26260 n1_7083_1328 n3_7083_1328 0.0
V26261 n1_7083_1727 n3_7083_1727 0.0
V26262 n1_7083_1760 n3_7083_1760 0.0
V26263 n1_7083_1916 n3_7083_1916 0.0
V26264 n1_7083_1943 n3_7083_1943 0.0
V26265 n1_7083_1976 n3_7083_1976 0.0
V26266 n1_7083_2159 n3_7083_2159 0.0
V26267 n1_7083_2192 n3_7083_2192 0.0
V26268 n1_7083_2375 n3_7083_2375 0.0
V26269 n1_7083_2408 n3_7083_2408 0.0
V26270 n1_7083_2543 n3_7083_2543 0.0
V26271 n1_7083_2564 n3_7083_2564 0.0
V26272 n1_7083_2591 n3_7083_2591 0.0
V26273 n1_7083_2624 n3_7083_2624 0.0
V26274 n1_7083_2807 n3_7083_2807 0.0
V26275 n1_7083_2840 n3_7083_2840 0.0
V26276 n1_7083_2974 n3_7083_2974 0.0
V26277 n1_7083_2996 n3_7083_2996 0.0
V26278 n1_7083_3023 n3_7083_3023 0.0
V26279 n1_7083_3056 n3_7083_3056 0.0
V26280 n1_7083_3239 n3_7083_3239 0.0
V26281 n1_7083_3272 n3_7083_3272 0.0
V26282 n1_7083_3455 n3_7083_3455 0.0
V26283 n1_7083_3488 n3_7083_3488 0.0
V26284 n1_7083_3644 n3_7083_3644 0.0
V26285 n1_7083_3671 n3_7083_3671 0.0
V26286 n1_7083_3704 n3_7083_3704 0.0
V26287 n1_7083_4103 n3_7083_4103 0.0
V26288 n1_7083_4136 n3_7083_4136 0.0
V26289 n1_7083_4292 n3_7083_4292 0.0
V26290 n1_7083_4319 n3_7083_4319 0.0
V26291 n1_7083_4352 n3_7083_4352 0.0
V26292 n1_7083_4535 n3_7083_4535 0.0
V26293 n1_7083_4568 n3_7083_4568 0.0
V26294 n1_7083_4724 n3_7083_4724 0.0
V26295 n1_7083_4751 n3_7083_4751 0.0
V26296 n1_7083_4784 n3_7083_4784 0.0
V26297 n1_7083_4967 n3_7083_4967 0.0
V26298 n1_7083_5000 n3_7083_5000 0.0
V26299 n1_7083_5183 n3_7083_5183 0.0
V26300 n1_7083_5216 n3_7083_5216 0.0
V26301 n1_7083_5372 n3_7083_5372 0.0
V26302 n1_7083_5399 n3_7083_5399 0.0
V26303 n1_7083_5432 n3_7083_5432 0.0
V26304 n1_7083_5566 n3_7083_5566 0.0
V26305 n1_7083_5588 n3_7083_5588 0.0
V26306 n1_7083_5615 n3_7083_5615 0.0
V26307 n1_7083_5648 n3_7083_5648 0.0
V26308 n1_7083_5831 n3_7083_5831 0.0
V26309 n1_7083_5864 n3_7083_5864 0.0
V26310 n1_7083_6263 n3_7083_6263 0.0
V26311 n1_7083_6296 n3_7083_6296 0.0
V26312 n1_7083_6479 n3_7083_6479 0.0
V26313 n1_7083_6512 n3_7083_6512 0.0
V26314 n1_7083_6646 n3_7083_6646 0.0
V26315 n1_7083_6695 n3_7083_6695 0.0
V26316 n1_7083_6728 n3_7083_6728 0.0
V26317 n1_7083_6911 n3_7083_6911 0.0
V26318 n1_7083_6944 n3_7083_6944 0.0
V26319 n1_7083_7127 n3_7083_7127 0.0
V26320 n1_7083_7160 n3_7083_7160 0.0
V26321 n1_7083_7343 n3_7083_7343 0.0
V26322 n1_7083_7376 n3_7083_7376 0.0
V26323 n1_7083_7559 n3_7083_7559 0.0
V26324 n1_7083_7592 n3_7083_7592 0.0
V26325 n1_7083_7775 n3_7083_7775 0.0
V26326 n1_7083_7808 n3_7083_7808 0.0
V26327 n1_7083_7822 n3_7083_7822 0.0
V26328 n1_7083_7964 n3_7083_7964 0.0
V26329 n1_7083_7991 n3_7083_7991 0.0
V26330 n1_7083_8024 n3_7083_8024 0.0
V26331 n1_7083_8207 n3_7083_8207 0.0
V26332 n1_7083_8240 n3_7083_8240 0.0
V26333 n1_7083_8456 n3_7083_8456 0.0
V26334 n1_7083_8639 n3_7083_8639 0.0
V26335 n1_7083_8672 n3_7083_8672 0.0
V26336 n1_7083_8855 n3_7083_8855 0.0
V26337 n1_7083_8888 n3_7083_8888 0.0
V26338 n1_7083_8902 n3_7083_8902 0.0
V26339 n1_7083_9044 n3_7083_9044 0.0
V26340 n1_7083_9071 n3_7083_9071 0.0
V26341 n1_7083_9104 n3_7083_9104 0.0
V26342 n1_7083_9287 n3_7083_9287 0.0
V26343 n1_7083_9320 n3_7083_9320 0.0
V26344 n1_7083_9503 n3_7083_9503 0.0
V26345 n1_7083_9536 n3_7083_9536 0.0
V26346 n1_7083_9719 n3_7083_9719 0.0
V26347 n1_7083_9752 n3_7083_9752 0.0
V26348 n1_7083_9935 n3_7083_9935 0.0
V26349 n1_7083_9968 n3_7083_9968 0.0
V26350 n1_7083_9982 n3_7083_9982 0.0
V26351 n1_7083_10124 n3_7083_10124 0.0
V26352 n1_7083_10151 n3_7083_10151 0.0
V26353 n1_7083_10184 n3_7083_10184 0.0
V26354 n1_7083_10367 n3_7083_10367 0.0
V26355 n1_7083_10400 n3_7083_10400 0.0
V26356 n1_7083_10799 n3_7083_10799 0.0
V26357 n1_7083_10832 n3_7083_10832 0.0
V26358 n1_7083_11015 n3_7083_11015 0.0
V26359 n1_7083_11048 n3_7083_11048 0.0
V26360 n1_7083_11204 n3_7083_11204 0.0
V26361 n1_7083_11231 n3_7083_11231 0.0
V26362 n1_7083_11264 n3_7083_11264 0.0
V26363 n1_7083_11447 n3_7083_11447 0.0
V26364 n1_7083_11480 n3_7083_11480 0.0
V26365 n1_7083_11663 n3_7083_11663 0.0
V26366 n1_7083_11696 n3_7083_11696 0.0
V26367 n1_7083_11879 n3_7083_11879 0.0
V26368 n1_7083_11912 n3_7083_11912 0.0
V26369 n1_7083_12095 n3_7083_12095 0.0
V26370 n1_7083_12128 n3_7083_12128 0.0
V26371 n1_7083_12284 n3_7083_12284 0.0
V26372 n1_7083_12311 n3_7083_12311 0.0
V26373 n1_7083_12344 n3_7083_12344 0.0
V26374 n1_7083_12527 n3_7083_12527 0.0
V26375 n1_7083_12560 n3_7083_12560 0.0
V26376 n1_7083_12743 n3_7083_12743 0.0
V26377 n1_7083_12959 n3_7083_12959 0.0
V26378 n1_7083_12992 n3_7083_12992 0.0
V26379 n1_7083_13175 n3_7083_13175 0.0
V26380 n1_7083_13208 n3_7083_13208 0.0
V26381 n1_7083_13391 n3_7083_13391 0.0
V26382 n1_7083_13424 n3_7083_13424 0.0
V26383 n1_7083_13580 n3_7083_13580 0.0
V26384 n1_7083_13607 n3_7083_13607 0.0
V26385 n1_7083_13640 n3_7083_13640 0.0
V26386 n1_7083_13823 n3_7083_13823 0.0
V26387 n1_7083_13856 n3_7083_13856 0.0
V26388 n1_7083_14039 n3_7083_14039 0.0
V26389 n1_7083_14072 n3_7083_14072 0.0
V26390 n1_7083_14255 n3_7083_14255 0.0
V26391 n1_7083_14288 n3_7083_14288 0.0
V26392 n1_7083_14471 n3_7083_14471 0.0
V26393 n1_7083_14504 n3_7083_14504 0.0
V26394 n1_7083_14553 n3_7083_14553 0.0
V26395 n1_7083_14687 n3_7083_14687 0.0
V26396 n1_7083_14720 n3_7083_14720 0.0
V26397 n1_7083_14903 n3_7083_14903 0.0
V26398 n1_7083_14936 n3_7083_14936 0.0
V26399 n1_7083_15335 n3_7083_15335 0.0
V26400 n1_7083_15368 n3_7083_15368 0.0
V26401 n1_7083_15551 n3_7083_15551 0.0
V26402 n1_7083_15584 n3_7083_15584 0.0
V26403 n1_7083_15740 n3_7083_15740 0.0
V26404 n1_7083_15767 n3_7083_15767 0.0
V26405 n1_7083_15800 n3_7083_15800 0.0
V26406 n1_7083_15956 n3_7083_15956 0.0
V26407 n1_7083_15983 n3_7083_15983 0.0
V26408 n1_7083_16016 n3_7083_16016 0.0
V26409 n1_7083_16172 n3_7083_16172 0.0
V26410 n1_7083_16199 n3_7083_16199 0.0
V26411 n1_7083_16232 n3_7083_16232 0.0
V26412 n1_7083_16415 n3_7083_16415 0.0
V26413 n1_7083_16448 n3_7083_16448 0.0
V26414 n1_7083_16631 n3_7083_16631 0.0
V26415 n1_7083_16664 n3_7083_16664 0.0
V26416 n1_7083_16847 n3_7083_16847 0.0
V26417 n1_7083_16880 n3_7083_16880 0.0
V26418 n1_7083_17063 n3_7083_17063 0.0
V26419 n1_7083_17096 n3_7083_17096 0.0
V26420 n1_7083_17230 n3_7083_17230 0.0
V26421 n1_7083_17468 n3_7083_17468 0.0
V26422 n1_7083_17495 n3_7083_17495 0.0
V26423 n1_7083_17528 n3_7083_17528 0.0
V26424 n1_7083_17711 n3_7083_17711 0.0
V26425 n1_7083_17744 n3_7083_17744 0.0
V26426 n1_7083_17927 n3_7083_17927 0.0
V26427 n1_7083_17960 n3_7083_17960 0.0
V26428 n1_7083_18143 n3_7083_18143 0.0
V26429 n1_7083_18176 n3_7083_18176 0.0
V26430 n1_7083_18359 n3_7083_18359 0.0
V26431 n1_7083_18392 n3_7083_18392 0.0
V26432 n1_7083_18526 n3_7083_18526 0.0
V26433 n1_7083_18527 n3_7083_18527 0.0
V26434 n1_7083_18548 n3_7083_18548 0.0
V26435 n1_7083_18575 n3_7083_18575 0.0
V26436 n1_7083_18608 n3_7083_18608 0.0
V26437 n1_7083_18764 n3_7083_18764 0.0
V26438 n1_7083_18791 n3_7083_18791 0.0
V26439 n1_7083_18824 n3_7083_18824 0.0
V26440 n1_7083_19007 n3_7083_19007 0.0
V26441 n1_7083_19040 n3_7083_19040 0.0
V26442 n1_7083_19196 n3_7083_19196 0.0
V26443 n1_7083_19223 n3_7083_19223 0.0
V26444 n1_7083_19256 n3_7083_19256 0.0
V26445 n1_7083_19390 n3_7083_19390 0.0
V26446 n1_7083_19439 n3_7083_19439 0.0
V26447 n1_7083_19472 n3_7083_19472 0.0
V26448 n1_7083_19871 n3_7083_19871 0.0
V26449 n1_7083_19904 n3_7083_19904 0.0
V26450 n1_7083_20087 n3_7083_20087 0.0
V26451 n1_7083_20120 n3_7083_20120 0.0
V26452 n1_7083_20303 n3_7083_20303 0.0
V26453 n1_7083_20336 n3_7083_20336 0.0
V26454 n1_7083_20519 n3_7083_20519 0.0
V26455 n1_7083_20552 n3_7083_20552 0.0
V26456 n1_7083_20687 n3_7083_20687 0.0
V26457 n1_7083_20735 n3_7083_20735 0.0
V26458 n1_7083_20768 n3_7083_20768 0.0
V26459 n1_7083_20951 n3_7083_20951 0.0
V26460 n1_7083_20984 n3_7083_20984 0.0
V26461 n1_7130_431 n3_7130_431 0.0
V26462 n1_7130_464 n3_7130_464 0.0
V26463 n1_7130_4967 n3_7130_4967 0.0
V26464 n1_7130_5000 n3_7130_5000 0.0
V26465 n1_7130_7160 n3_7130_7160 0.0
V26466 n1_7130_9503 n3_7130_9503 0.0
V26467 n1_7130_9536 n3_7130_9536 0.0
V26468 n1_7130_11663 n3_7130_11663 0.0
V26469 n1_7130_11696 n3_7130_11696 0.0
V26470 n1_7130_14039 n3_7130_14039 0.0
V26471 n1_7130_16172 n3_7130_16172 0.0
V26472 n1_7130_16199 n3_7130_16199 0.0
V26473 n1_7130_16232 n3_7130_16232 0.0
V26474 n1_7130_18392 n3_7130_18392 0.0
V26475 n1_7130_18526 n3_7130_18526 0.0
V26476 n1_7130_18527 n3_7130_18527 0.0
V26477 n1_7130_18548 n3_7130_18548 0.0
V26478 n1_7130_20687 n3_7130_20687 0.0
V26479 n1_7130_20735 n3_7130_20735 0.0
V26480 n1_7130_20768 n3_7130_20768 0.0
V26481 n1_7271_215 n3_7271_215 0.0
V26482 n1_7271_248 n3_7271_248 0.0
V26483 n1_7271_383 n3_7271_383 0.0
V26484 n1_7271_431 n3_7271_431 0.0
V26485 n1_7271_647 n3_7271_647 0.0
V26486 n1_7271_680 n3_7271_680 0.0
V26487 n1_7271_863 n3_7271_863 0.0
V26488 n1_7271_896 n3_7271_896 0.0
V26489 n1_7271_1079 n3_7271_1079 0.0
V26490 n1_7271_1112 n3_7271_1112 0.0
V26491 n1_7271_1295 n3_7271_1295 0.0
V26492 n1_7271_1328 n3_7271_1328 0.0
V26493 n1_7271_1511 n3_7271_1511 0.0
V26494 n1_7271_1544 n3_7271_1544 0.0
V26495 n1_7271_1727 n3_7271_1727 0.0
V26496 n1_7271_1760 n3_7271_1760 0.0
V26497 n1_7271_1916 n3_7271_1916 0.0
V26498 n1_7271_1943 n3_7271_1943 0.0
V26499 n1_7271_1976 n3_7271_1976 0.0
V26500 n1_7271_2159 n3_7271_2159 0.0
V26501 n1_7271_2192 n3_7271_2192 0.0
V26502 n1_7271_2375 n3_7271_2375 0.0
V26503 n1_7271_2408 n3_7271_2408 0.0
V26504 n1_7271_2543 n3_7271_2543 0.0
V26505 n1_7271_2564 n3_7271_2564 0.0
V26506 n1_7271_2591 n3_7271_2591 0.0
V26507 n1_7271_2624 n3_7271_2624 0.0
V26508 n1_7271_2807 n3_7271_2807 0.0
V26509 n1_7271_2840 n3_7271_2840 0.0
V26510 n1_7271_2974 n3_7271_2974 0.0
V26511 n1_7271_2996 n3_7271_2996 0.0
V26512 n1_7271_3023 n3_7271_3023 0.0
V26513 n1_7271_3056 n3_7271_3056 0.0
V26514 n1_7271_3239 n3_7271_3239 0.0
V26515 n1_7271_3272 n3_7271_3272 0.0
V26516 n1_7271_3455 n3_7271_3455 0.0
V26517 n1_7271_3488 n3_7271_3488 0.0
V26518 n1_7271_3644 n3_7271_3644 0.0
V26519 n1_7271_3671 n3_7271_3671 0.0
V26520 n1_7271_3704 n3_7271_3704 0.0
V26521 n1_7271_3887 n3_7271_3887 0.0
V26522 n1_7271_3920 n3_7271_3920 0.0
V26523 n1_7271_4103 n3_7271_4103 0.0
V26524 n1_7271_4136 n3_7271_4136 0.0
V26525 n1_7271_4292 n3_7271_4292 0.0
V26526 n1_7271_4319 n3_7271_4319 0.0
V26527 n1_7271_4352 n3_7271_4352 0.0
V26528 n1_7271_4535 n3_7271_4535 0.0
V26529 n1_7271_4568 n3_7271_4568 0.0
V26530 n1_7271_4724 n3_7271_4724 0.0
V26531 n1_7271_4751 n3_7271_4751 0.0
V26532 n1_7271_4784 n3_7271_4784 0.0
V26533 n1_7271_5000 n3_7271_5000 0.0
V26534 n1_7271_5183 n3_7271_5183 0.0
V26535 n1_7271_5216 n3_7271_5216 0.0
V26536 n1_7271_5372 n3_7271_5372 0.0
V26537 n1_7271_5399 n3_7271_5399 0.0
V26538 n1_7271_5432 n3_7271_5432 0.0
V26539 n1_7271_5566 n3_7271_5566 0.0
V26540 n1_7271_5588 n3_7271_5588 0.0
V26541 n1_7271_5615 n3_7271_5615 0.0
V26542 n1_7271_5648 n3_7271_5648 0.0
V26543 n1_7271_5831 n3_7271_5831 0.0
V26544 n1_7271_5864 n3_7271_5864 0.0
V26545 n1_7271_6047 n3_7271_6047 0.0
V26546 n1_7271_6080 n3_7271_6080 0.0
V26547 n1_7271_6263 n3_7271_6263 0.0
V26548 n1_7271_6296 n3_7271_6296 0.0
V26549 n1_7271_6479 n3_7271_6479 0.0
V26550 n1_7271_6512 n3_7271_6512 0.0
V26551 n1_7271_6646 n3_7271_6646 0.0
V26552 n1_7271_6695 n3_7271_6695 0.0
V26553 n1_7271_6728 n3_7271_6728 0.0
V26554 n1_7271_6911 n3_7271_6911 0.0
V26555 n1_7271_6944 n3_7271_6944 0.0
V26556 n1_7271_7127 n3_7271_7127 0.0
V26557 n1_7271_7160 n3_7271_7160 0.0
V26558 n1_7271_7343 n3_7271_7343 0.0
V26559 n1_7271_7376 n3_7271_7376 0.0
V26560 n1_7271_7559 n3_7271_7559 0.0
V26561 n1_7271_7592 n3_7271_7592 0.0
V26562 n1_7271_7775 n3_7271_7775 0.0
V26563 n1_7271_7808 n3_7271_7808 0.0
V26564 n1_7271_7822 n3_7271_7822 0.0
V26565 n1_7271_7964 n3_7271_7964 0.0
V26566 n1_7271_7991 n3_7271_7991 0.0
V26567 n1_7271_8024 n3_7271_8024 0.0
V26568 n1_7271_8207 n3_7271_8207 0.0
V26569 n1_7271_8240 n3_7271_8240 0.0
V26570 n1_7271_8423 n3_7271_8423 0.0
V26571 n1_7271_8456 n3_7271_8456 0.0
V26572 n1_7271_8639 n3_7271_8639 0.0
V26573 n1_7271_8672 n3_7271_8672 0.0
V26574 n1_7271_8855 n3_7271_8855 0.0
V26575 n1_7271_8888 n3_7271_8888 0.0
V26576 n1_7271_8902 n3_7271_8902 0.0
V26577 n1_7271_9044 n3_7271_9044 0.0
V26578 n1_7271_9071 n3_7271_9071 0.0
V26579 n1_7271_9104 n3_7271_9104 0.0
V26580 n1_7271_9287 n3_7271_9287 0.0
V26581 n1_7271_9320 n3_7271_9320 0.0
V26582 n1_7271_9503 n3_7271_9503 0.0
V26583 n1_7271_9536 n3_7271_9536 0.0
V26584 n1_7271_9719 n3_7271_9719 0.0
V26585 n1_7271_9752 n3_7271_9752 0.0
V26586 n1_7271_9935 n3_7271_9935 0.0
V26587 n1_7271_9968 n3_7271_9968 0.0
V26588 n1_7271_9982 n3_7271_9982 0.0
V26589 n1_7271_10124 n3_7271_10124 0.0
V26590 n1_7271_10151 n3_7271_10151 0.0
V26591 n1_7271_10184 n3_7271_10184 0.0
V26592 n1_7271_10367 n3_7271_10367 0.0
V26593 n1_7271_10400 n3_7271_10400 0.0
V26594 n1_7271_10616 n3_7271_10616 0.0
V26595 n1_7271_10799 n3_7271_10799 0.0
V26596 n1_7271_10832 n3_7271_10832 0.0
V26597 n1_7271_11015 n3_7271_11015 0.0
V26598 n1_7271_11048 n3_7271_11048 0.0
V26599 n1_7271_11204 n3_7271_11204 0.0
V26600 n1_7271_11231 n3_7271_11231 0.0
V26601 n1_7271_11264 n3_7271_11264 0.0
V26602 n1_7271_11447 n3_7271_11447 0.0
V26603 n1_7271_11480 n3_7271_11480 0.0
V26604 n1_7271_11663 n3_7271_11663 0.0
V26605 n1_7271_11696 n3_7271_11696 0.0
V26606 n1_7271_11879 n3_7271_11879 0.0
V26607 n1_7271_11912 n3_7271_11912 0.0
V26608 n1_7271_12095 n3_7271_12095 0.0
V26609 n1_7271_12128 n3_7271_12128 0.0
V26610 n1_7271_12284 n3_7271_12284 0.0
V26611 n1_7271_12311 n3_7271_12311 0.0
V26612 n1_7271_12344 n3_7271_12344 0.0
V26613 n1_7271_12527 n3_7271_12527 0.0
V26614 n1_7271_12560 n3_7271_12560 0.0
V26615 n1_7271_12743 n3_7271_12743 0.0
V26616 n1_7271_12776 n3_7271_12776 0.0
V26617 n1_7271_12959 n3_7271_12959 0.0
V26618 n1_7271_12992 n3_7271_12992 0.0
V26619 n1_7271_13175 n3_7271_13175 0.0
V26620 n1_7271_13208 n3_7271_13208 0.0
V26621 n1_7271_13391 n3_7271_13391 0.0
V26622 n1_7271_13424 n3_7271_13424 0.0
V26623 n1_7271_13580 n3_7271_13580 0.0
V26624 n1_7271_13607 n3_7271_13607 0.0
V26625 n1_7271_13640 n3_7271_13640 0.0
V26626 n1_7271_13823 n3_7271_13823 0.0
V26627 n1_7271_13856 n3_7271_13856 0.0
V26628 n1_7271_14039 n3_7271_14039 0.0
V26629 n1_7271_14072 n3_7271_14072 0.0
V26630 n1_7271_14255 n3_7271_14255 0.0
V26631 n1_7271_14288 n3_7271_14288 0.0
V26632 n1_7271_14471 n3_7271_14471 0.0
V26633 n1_7271_14504 n3_7271_14504 0.0
V26634 n1_7271_14553 n3_7271_14553 0.0
V26635 n1_7271_14687 n3_7271_14687 0.0
V26636 n1_7271_14720 n3_7271_14720 0.0
V26637 n1_7271_14903 n3_7271_14903 0.0
V26638 n1_7271_14936 n3_7271_14936 0.0
V26639 n1_7271_15119 n3_7271_15119 0.0
V26640 n1_7271_15152 n3_7271_15152 0.0
V26641 n1_7271_15335 n3_7271_15335 0.0
V26642 n1_7271_15368 n3_7271_15368 0.0
V26643 n1_7271_15551 n3_7271_15551 0.0
V26644 n1_7271_15584 n3_7271_15584 0.0
V26645 n1_7271_15740 n3_7271_15740 0.0
V26646 n1_7271_15767 n3_7271_15767 0.0
V26647 n1_7271_15800 n3_7271_15800 0.0
V26648 n1_7271_15956 n3_7271_15956 0.0
V26649 n1_7271_15983 n3_7271_15983 0.0
V26650 n1_7271_16016 n3_7271_16016 0.0
V26651 n1_7271_16172 n3_7271_16172 0.0
V26652 n1_7271_16199 n3_7271_16199 0.0
V26653 n1_7271_16415 n3_7271_16415 0.0
V26654 n1_7271_16448 n3_7271_16448 0.0
V26655 n1_7271_16631 n3_7271_16631 0.0
V26656 n1_7271_16664 n3_7271_16664 0.0
V26657 n1_7271_16847 n3_7271_16847 0.0
V26658 n1_7271_16880 n3_7271_16880 0.0
V26659 n1_7271_17063 n3_7271_17063 0.0
V26660 n1_7271_17096 n3_7271_17096 0.0
V26661 n1_7271_17230 n3_7271_17230 0.0
V26662 n1_7271_17252 n3_7271_17252 0.0
V26663 n1_7271_17279 n3_7271_17279 0.0
V26664 n1_7271_17312 n3_7271_17312 0.0
V26665 n1_7271_17468 n3_7271_17468 0.0
V26666 n1_7271_17495 n3_7271_17495 0.0
V26667 n1_7271_17528 n3_7271_17528 0.0
V26668 n1_7271_17711 n3_7271_17711 0.0
V26669 n1_7271_17744 n3_7271_17744 0.0
V26670 n1_7271_17927 n3_7271_17927 0.0
V26671 n1_7271_17960 n3_7271_17960 0.0
V26672 n1_7271_18143 n3_7271_18143 0.0
V26673 n1_7271_18176 n3_7271_18176 0.0
V26674 n1_7271_18359 n3_7271_18359 0.0
V26675 n1_7271_18392 n3_7271_18392 0.0
V26676 n1_7271_18526 n3_7271_18526 0.0
V26677 n1_7271_18527 n3_7271_18527 0.0
V26678 n1_7271_18548 n3_7271_18548 0.0
V26679 n1_7271_18575 n3_7271_18575 0.0
V26680 n1_7271_18608 n3_7271_18608 0.0
V26681 n1_7271_18764 n3_7271_18764 0.0
V26682 n1_7271_18791 n3_7271_18791 0.0
V26683 n1_7271_18824 n3_7271_18824 0.0
V26684 n1_7271_19007 n3_7271_19007 0.0
V26685 n1_7271_19040 n3_7271_19040 0.0
V26686 n1_7271_19196 n3_7271_19196 0.0
V26687 n1_7271_19223 n3_7271_19223 0.0
V26688 n1_7271_19256 n3_7271_19256 0.0
V26689 n1_7271_19390 n3_7271_19390 0.0
V26690 n1_7271_19439 n3_7271_19439 0.0
V26691 n1_7271_19472 n3_7271_19472 0.0
V26692 n1_7271_19655 n3_7271_19655 0.0
V26693 n1_7271_19688 n3_7271_19688 0.0
V26694 n1_7271_19871 n3_7271_19871 0.0
V26695 n1_7271_19904 n3_7271_19904 0.0
V26696 n1_7271_20087 n3_7271_20087 0.0
V26697 n1_7271_20120 n3_7271_20120 0.0
V26698 n1_7271_20303 n3_7271_20303 0.0
V26699 n1_7271_20336 n3_7271_20336 0.0
V26700 n1_7271_20519 n3_7271_20519 0.0
V26701 n1_7271_20552 n3_7271_20552 0.0
V26702 n1_7271_20687 n3_7271_20687 0.0
V26703 n1_7271_20768 n3_7271_20768 0.0
V26704 n1_7271_20951 n3_7271_20951 0.0
V26705 n1_7271_20984 n3_7271_20984 0.0
V26706 n1_7364_215 n3_7364_215 0.0
V26707 n1_7364_248 n3_7364_248 0.0
V26708 n1_7364_383 n3_7364_383 0.0
V26709 n1_7364_431 n3_7364_431 0.0
V26710 n1_7364_464 n3_7364_464 0.0
V26711 n1_7364_647 n3_7364_647 0.0
V26712 n1_7364_680 n3_7364_680 0.0
V26713 n1_7364_863 n3_7364_863 0.0
V26714 n1_7364_896 n3_7364_896 0.0
V26715 n1_7364_1079 n3_7364_1079 0.0
V26716 n1_7364_1112 n3_7364_1112 0.0
V26717 n1_7364_1295 n3_7364_1295 0.0
V26718 n1_7364_1328 n3_7364_1328 0.0
V26719 n1_7364_1511 n3_7364_1511 0.0
V26720 n1_7364_1544 n3_7364_1544 0.0
V26721 n1_7364_1727 n3_7364_1727 0.0
V26722 n1_7364_1760 n3_7364_1760 0.0
V26723 n1_7364_1916 n3_7364_1916 0.0
V26724 n1_7364_1943 n3_7364_1943 0.0
V26725 n1_7364_1976 n3_7364_1976 0.0
V26726 n1_7364_2159 n3_7364_2159 0.0
V26727 n1_7364_2192 n3_7364_2192 0.0
V26728 n1_7364_2375 n3_7364_2375 0.0
V26729 n1_7364_2408 n3_7364_2408 0.0
V26730 n1_7364_2543 n3_7364_2543 0.0
V26731 n1_7364_2564 n3_7364_2564 0.0
V26732 n1_7364_2591 n3_7364_2591 0.0
V26733 n1_7364_2624 n3_7364_2624 0.0
V26734 n1_7364_18526 n3_7364_18526 0.0
V26735 n1_7364_18527 n3_7364_18527 0.0
V26736 n1_7364_18575 n3_7364_18575 0.0
V26737 n1_7364_18608 n3_7364_18608 0.0
V26738 n1_7364_18764 n3_7364_18764 0.0
V26739 n1_7364_18791 n3_7364_18791 0.0
V26740 n1_7364_18824 n3_7364_18824 0.0
V26741 n1_7364_19007 n3_7364_19007 0.0
V26742 n1_7364_19040 n3_7364_19040 0.0
V26743 n1_7364_19223 n3_7364_19223 0.0
V26744 n1_7364_19256 n3_7364_19256 0.0
V26745 n1_7364_19390 n3_7364_19390 0.0
V26746 n1_7364_19439 n3_7364_19439 0.0
V26747 n1_7364_19472 n3_7364_19472 0.0
V26748 n1_7364_19655 n3_7364_19655 0.0
V26749 n1_7364_19688 n3_7364_19688 0.0
V26750 n1_7364_19871 n3_7364_19871 0.0
V26751 n1_7364_19904 n3_7364_19904 0.0
V26752 n1_7364_20087 n3_7364_20087 0.0
V26753 n1_7364_20120 n3_7364_20120 0.0
V26754 n1_7364_20303 n3_7364_20303 0.0
V26755 n1_7364_20336 n3_7364_20336 0.0
V26756 n1_7364_20519 n3_7364_20519 0.0
V26757 n1_7364_20552 n3_7364_20552 0.0
V26758 n1_7364_20687 n3_7364_20687 0.0
V26759 n1_7364_20735 n3_7364_20735 0.0
V26760 n1_7364_20768 n3_7364_20768 0.0
V26761 n1_7364_20951 n3_7364_20951 0.0
V26762 n1_7364_20984 n3_7364_20984 0.0
V26763 n1_9150_215 n3_9150_215 0.0
V26764 n1_9150_248 n3_9150_248 0.0
V26765 n1_9150_383 n3_9150_383 0.0
V26766 n1_9150_431 n3_9150_431 0.0
V26767 n1_9150_464 n3_9150_464 0.0
V26768 n1_9150_647 n3_9150_647 0.0
V26769 n1_9150_680 n3_9150_680 0.0
V26770 n1_9150_863 n3_9150_863 0.0
V26771 n1_9150_896 n3_9150_896 0.0
V26772 n1_9150_1079 n3_9150_1079 0.0
V26773 n1_9150_1112 n3_9150_1112 0.0
V26774 n1_9150_1295 n3_9150_1295 0.0
V26775 n1_9150_1328 n3_9150_1328 0.0
V26776 n1_9150_1511 n3_9150_1511 0.0
V26777 n1_9150_1544 n3_9150_1544 0.0
V26778 n1_9150_1727 n3_9150_1727 0.0
V26779 n1_9150_1760 n3_9150_1760 0.0
V26780 n1_9150_1894 n3_9150_1894 0.0
V26781 n1_9150_1943 n3_9150_1943 0.0
V26782 n1_9150_1976 n3_9150_1976 0.0
V26783 n1_9150_2159 n3_9150_2159 0.0
V26784 n1_9150_2192 n3_9150_2192 0.0
V26785 n1_9150_2375 n3_9150_2375 0.0
V26786 n1_9150_2408 n3_9150_2408 0.0
V26787 n1_9150_2543 n3_9150_2543 0.0
V26788 n1_9150_2564 n3_9150_2564 0.0
V26789 n1_9150_2591 n3_9150_2591 0.0
V26790 n1_9150_2624 n3_9150_2624 0.0
V26791 n1_9150_18527 n3_9150_18527 0.0
V26792 n1_9150_18548 n3_9150_18548 0.0
V26793 n1_9150_18575 n3_9150_18575 0.0
V26794 n1_9150_18608 n3_9150_18608 0.0
V26795 n1_9150_18764 n3_9150_18764 0.0
V26796 n1_9150_18791 n3_9150_18791 0.0
V26797 n1_9150_18824 n3_9150_18824 0.0
V26798 n1_9150_19007 n3_9150_19007 0.0
V26799 n1_9150_19040 n3_9150_19040 0.0
V26800 n1_9150_19223 n3_9150_19223 0.0
V26801 n1_9150_19256 n3_9150_19256 0.0
V26802 n1_9150_19412 n3_9150_19412 0.0
V26803 n1_9150_19439 n3_9150_19439 0.0
V26804 n1_9150_19472 n3_9150_19472 0.0
V26805 n1_9150_19655 n3_9150_19655 0.0
V26806 n1_9150_19688 n3_9150_19688 0.0
V26807 n1_9150_19871 n3_9150_19871 0.0
V26808 n1_9150_19904 n3_9150_19904 0.0
V26809 n1_9150_20087 n3_9150_20087 0.0
V26810 n1_9150_20120 n3_9150_20120 0.0
V26811 n1_9150_20303 n3_9150_20303 0.0
V26812 n1_9150_20336 n3_9150_20336 0.0
V26813 n1_9150_20519 n3_9150_20519 0.0
V26814 n1_9150_20552 n3_9150_20552 0.0
V26815 n1_9150_20687 n3_9150_20687 0.0
V26816 n1_9150_20735 n3_9150_20735 0.0
V26817 n1_9150_20768 n3_9150_20768 0.0
V26818 n1_9150_20951 n3_9150_20951 0.0
V26819 n1_9150_20984 n3_9150_20984 0.0
V26820 n1_9333_215 n3_9333_215 0.0
V26821 n1_9333_248 n3_9333_248 0.0
V26822 n1_9333_383 n3_9333_383 0.0
V26823 n1_9333_431 n3_9333_431 0.0
V26824 n1_9333_464 n3_9333_464 0.0
V26825 n1_9333_647 n3_9333_647 0.0
V26826 n1_9333_680 n3_9333_680 0.0
V26827 n1_9333_863 n3_9333_863 0.0
V26828 n1_9333_896 n3_9333_896 0.0
V26829 n1_9333_1079 n3_9333_1079 0.0
V26830 n1_9333_1112 n3_9333_1112 0.0
V26831 n1_9333_1295 n3_9333_1295 0.0
V26832 n1_9333_1328 n3_9333_1328 0.0
V26833 n1_9333_1727 n3_9333_1727 0.0
V26834 n1_9333_1760 n3_9333_1760 0.0
V26835 n1_9333_1894 n3_9333_1894 0.0
V26836 n1_9333_1916 n3_9333_1916 0.0
V26837 n1_9333_1943 n3_9333_1943 0.0
V26838 n1_9333_1976 n3_9333_1976 0.0
V26839 n1_9333_2159 n3_9333_2159 0.0
V26840 n1_9333_2192 n3_9333_2192 0.0
V26841 n1_9333_2375 n3_9333_2375 0.0
V26842 n1_9333_2408 n3_9333_2408 0.0
V26843 n1_9333_2543 n3_9333_2543 0.0
V26844 n1_9333_2564 n3_9333_2564 0.0
V26845 n1_9333_2591 n3_9333_2591 0.0
V26846 n1_9333_2624 n3_9333_2624 0.0
V26847 n1_9333_2807 n3_9333_2807 0.0
V26848 n1_9333_2840 n3_9333_2840 0.0
V26849 n1_9333_2996 n3_9333_2996 0.0
V26850 n1_9333_3023 n3_9333_3023 0.0
V26851 n1_9333_3056 n3_9333_3056 0.0
V26852 n1_9333_3239 n3_9333_3239 0.0
V26853 n1_9333_3272 n3_9333_3272 0.0
V26854 n1_9333_3455 n3_9333_3455 0.0
V26855 n1_9333_3488 n3_9333_3488 0.0
V26856 n1_9333_3644 n3_9333_3644 0.0
V26857 n1_9333_3671 n3_9333_3671 0.0
V26858 n1_9333_3704 n3_9333_3704 0.0
V26859 n1_9333_4103 n3_9333_4103 0.0
V26860 n1_9333_4136 n3_9333_4136 0.0
V26861 n1_9333_4292 n3_9333_4292 0.0
V26862 n1_9333_4319 n3_9333_4319 0.0
V26863 n1_9333_4352 n3_9333_4352 0.0
V26864 n1_9333_4535 n3_9333_4535 0.0
V26865 n1_9333_4568 n3_9333_4568 0.0
V26866 n1_9333_4724 n3_9333_4724 0.0
V26867 n1_9333_4751 n3_9333_4751 0.0
V26868 n1_9333_4784 n3_9333_4784 0.0
V26869 n1_9333_4967 n3_9333_4967 0.0
V26870 n1_9333_5000 n3_9333_5000 0.0
V26871 n1_9333_5183 n3_9333_5183 0.0
V26872 n1_9333_5216 n3_9333_5216 0.0
V26873 n1_9333_5350 n3_9333_5350 0.0
V26874 n1_9333_5372 n3_9333_5372 0.0
V26875 n1_9333_5399 n3_9333_5399 0.0
V26876 n1_9333_5432 n3_9333_5432 0.0
V26877 n1_9333_5588 n3_9333_5588 0.0
V26878 n1_9333_5615 n3_9333_5615 0.0
V26879 n1_9333_5648 n3_9333_5648 0.0
V26880 n1_9333_5831 n3_9333_5831 0.0
V26881 n1_9333_5864 n3_9333_5864 0.0
V26882 n1_9333_6263 n3_9333_6263 0.0
V26883 n1_9333_6296 n3_9333_6296 0.0
V26884 n1_9333_6479 n3_9333_6479 0.0
V26885 n1_9333_6512 n3_9333_6512 0.0
V26886 n1_9333_6668 n3_9333_6668 0.0
V26887 n1_9333_6695 n3_9333_6695 0.0
V26888 n1_9333_6728 n3_9333_6728 0.0
V26889 n1_9333_6911 n3_9333_6911 0.0
V26890 n1_9333_6944 n3_9333_6944 0.0
V26891 n1_9333_7100 n3_9333_7100 0.0
V26892 n1_9333_7127 n3_9333_7127 0.0
V26893 n1_9333_7160 n3_9333_7160 0.0
V26894 n1_9333_7316 n3_9333_7316 0.0
V26895 n1_9333_7343 n3_9333_7343 0.0
V26896 n1_9333_7376 n3_9333_7376 0.0
V26897 n1_9333_7532 n3_9333_7532 0.0
V26898 n1_9333_7559 n3_9333_7559 0.0
V26899 n1_9333_7592 n3_9333_7592 0.0
V26900 n1_9333_7775 n3_9333_7775 0.0
V26901 n1_9333_7808 n3_9333_7808 0.0
V26902 n1_9333_7991 n3_9333_7991 0.0
V26903 n1_9333_8024 n3_9333_8024 0.0
V26904 n1_9333_8207 n3_9333_8207 0.0
V26905 n1_9333_8240 n3_9333_8240 0.0
V26906 n1_9333_8456 n3_9333_8456 0.0
V26907 n1_9333_8639 n3_9333_8639 0.0
V26908 n1_9333_8672 n3_9333_8672 0.0
V26909 n1_9333_8855 n3_9333_8855 0.0
V26910 n1_9333_8888 n3_9333_8888 0.0
V26911 n1_9333_9071 n3_9333_9071 0.0
V26912 n1_9333_9104 n3_9333_9104 0.0
V26913 n1_9333_9287 n3_9333_9287 0.0
V26914 n1_9333_9320 n3_9333_9320 0.0
V26915 n1_9333_9503 n3_9333_9503 0.0
V26916 n1_9333_9536 n3_9333_9536 0.0
V26917 n1_9333_9719 n3_9333_9719 0.0
V26918 n1_9333_9752 n3_9333_9752 0.0
V26919 n1_9333_9935 n3_9333_9935 0.0
V26920 n1_9333_9968 n3_9333_9968 0.0
V26921 n1_9333_10151 n3_9333_10151 0.0
V26922 n1_9333_10184 n3_9333_10184 0.0
V26923 n1_9333_10367 n3_9333_10367 0.0
V26924 n1_9333_10400 n3_9333_10400 0.0
V26925 n1_9333_10799 n3_9333_10799 0.0
V26926 n1_9333_10832 n3_9333_10832 0.0
V26927 n1_9333_11015 n3_9333_11015 0.0
V26928 n1_9333_11048 n3_9333_11048 0.0
V26929 n1_9333_11231 n3_9333_11231 0.0
V26930 n1_9333_11264 n3_9333_11264 0.0
V26931 n1_9333_11447 n3_9333_11447 0.0
V26932 n1_9333_11480 n3_9333_11480 0.0
V26933 n1_9333_11663 n3_9333_11663 0.0
V26934 n1_9333_11696 n3_9333_11696 0.0
V26935 n1_9333_11879 n3_9333_11879 0.0
V26936 n1_9333_11912 n3_9333_11912 0.0
V26937 n1_9333_12095 n3_9333_12095 0.0
V26938 n1_9333_12128 n3_9333_12128 0.0
V26939 n1_9333_12311 n3_9333_12311 0.0
V26940 n1_9333_12344 n3_9333_12344 0.0
V26941 n1_9333_12527 n3_9333_12527 0.0
V26942 n1_9333_12560 n3_9333_12560 0.0
V26943 n1_9333_12743 n3_9333_12743 0.0
V26944 n1_9333_12959 n3_9333_12959 0.0
V26945 n1_9333_12992 n3_9333_12992 0.0
V26946 n1_9333_13175 n3_9333_13175 0.0
V26947 n1_9333_13208 n3_9333_13208 0.0
V26948 n1_9333_13391 n3_9333_13391 0.0
V26949 n1_9333_13424 n3_9333_13424 0.0
V26950 n1_9333_13607 n3_9333_13607 0.0
V26951 n1_9333_13640 n3_9333_13640 0.0
V26952 n1_9333_13796 n3_9333_13796 0.0
V26953 n1_9333_13823 n3_9333_13823 0.0
V26954 n1_9333_13856 n3_9333_13856 0.0
V26955 n1_9333_13990 n3_9333_13990 0.0
V26956 n1_9333_14012 n3_9333_14012 0.0
V26957 n1_9333_14039 n3_9333_14039 0.0
V26958 n1_9333_14072 n3_9333_14072 0.0
V26959 n1_9333_14228 n3_9333_14228 0.0
V26960 n1_9333_14255 n3_9333_14255 0.0
V26961 n1_9333_14288 n3_9333_14288 0.0
V26962 n1_9333_14471 n3_9333_14471 0.0
V26963 n1_9333_14504 n3_9333_14504 0.0
V26964 n1_9333_14660 n3_9333_14660 0.0
V26965 n1_9333_14687 n3_9333_14687 0.0
V26966 n1_9333_14720 n3_9333_14720 0.0
V26967 n1_9333_14903 n3_9333_14903 0.0
V26968 n1_9333_14936 n3_9333_14936 0.0
V26969 n1_9333_15335 n3_9333_15335 0.0
V26970 n1_9333_15368 n3_9333_15368 0.0
V26971 n1_9333_15551 n3_9333_15551 0.0
V26972 n1_9333_15584 n3_9333_15584 0.0
V26973 n1_9333_15740 n3_9333_15740 0.0
V26974 n1_9333_15767 n3_9333_15767 0.0
V26975 n1_9333_15800 n3_9333_15800 0.0
V26976 n1_9333_15934 n3_9333_15934 0.0
V26977 n1_9333_15956 n3_9333_15956 0.0
V26978 n1_9333_15983 n3_9333_15983 0.0
V26979 n1_9333_16016 n3_9333_16016 0.0
V26980 n1_9333_16172 n3_9333_16172 0.0
V26981 n1_9333_16199 n3_9333_16199 0.0
V26982 n1_9333_16232 n3_9333_16232 0.0
V26983 n1_9333_16415 n3_9333_16415 0.0
V26984 n1_9333_16448 n3_9333_16448 0.0
V26985 n1_9333_16631 n3_9333_16631 0.0
V26986 n1_9333_16664 n3_9333_16664 0.0
V26987 n1_9333_16847 n3_9333_16847 0.0
V26988 n1_9333_16880 n3_9333_16880 0.0
V26989 n1_9333_17063 n3_9333_17063 0.0
V26990 n1_9333_17096 n3_9333_17096 0.0
V26991 n1_9333_17230 n3_9333_17230 0.0
V26992 n1_9333_17468 n3_9333_17468 0.0
V26993 n1_9333_17495 n3_9333_17495 0.0
V26994 n1_9333_17528 n3_9333_17528 0.0
V26995 n1_9333_17711 n3_9333_17711 0.0
V26996 n1_9333_17744 n3_9333_17744 0.0
V26997 n1_9333_17927 n3_9333_17927 0.0
V26998 n1_9333_17960 n3_9333_17960 0.0
V26999 n1_9333_18143 n3_9333_18143 0.0
V27000 n1_9333_18176 n3_9333_18176 0.0
V27001 n1_9333_18359 n3_9333_18359 0.0
V27002 n1_9333_18392 n3_9333_18392 0.0
V27003 n1_9333_18527 n3_9333_18527 0.0
V27004 n1_9333_18548 n3_9333_18548 0.0
V27005 n1_9333_18575 n3_9333_18575 0.0
V27006 n1_9333_18608 n3_9333_18608 0.0
V27007 n1_9333_18764 n3_9333_18764 0.0
V27008 n1_9333_18791 n3_9333_18791 0.0
V27009 n1_9333_18824 n3_9333_18824 0.0
V27010 n1_9333_19007 n3_9333_19007 0.0
V27011 n1_9333_19040 n3_9333_19040 0.0
V27012 n1_9333_19223 n3_9333_19223 0.0
V27013 n1_9333_19256 n3_9333_19256 0.0
V27014 n1_9333_19412 n3_9333_19412 0.0
V27015 n1_9333_19439 n3_9333_19439 0.0
V27016 n1_9333_19472 n3_9333_19472 0.0
V27017 n1_9333_19871 n3_9333_19871 0.0
V27018 n1_9333_19904 n3_9333_19904 0.0
V27019 n1_9333_20087 n3_9333_20087 0.0
V27020 n1_9333_20120 n3_9333_20120 0.0
V27021 n1_9333_20303 n3_9333_20303 0.0
V27022 n1_9333_20336 n3_9333_20336 0.0
V27023 n1_9333_20519 n3_9333_20519 0.0
V27024 n1_9333_20552 n3_9333_20552 0.0
V27025 n1_9333_20687 n3_9333_20687 0.0
V27026 n1_9333_20735 n3_9333_20735 0.0
V27027 n1_9333_20768 n3_9333_20768 0.0
V27028 n1_9333_20951 n3_9333_20951 0.0
V27029 n1_9333_20984 n3_9333_20984 0.0
V27030 n1_9380_431 n3_9380_431 0.0
V27031 n1_9380_464 n3_9380_464 0.0
V27032 n1_9380_4967 n3_9380_4967 0.0
V27033 n1_9380_5000 n3_9380_5000 0.0
V27034 n1_9380_7160 n3_9380_7160 0.0
V27035 n1_9380_9503 n3_9380_9503 0.0
V27036 n1_9380_9536 n3_9380_9536 0.0
V27037 n1_9380_11663 n3_9380_11663 0.0
V27038 n1_9380_11696 n3_9380_11696 0.0
V27039 n1_9380_13990 n3_9380_13990 0.0
V27040 n1_9380_14012 n3_9380_14012 0.0
V27041 n1_9380_14039 n3_9380_14039 0.0
V27042 n1_9380_16172 n3_9380_16172 0.0
V27043 n1_9380_16199 n3_9380_16199 0.0
V27044 n1_9380_16232 n3_9380_16232 0.0
V27045 n1_9380_18392 n3_9380_18392 0.0
V27046 n1_9380_18527 n3_9380_18527 0.0
V27047 n1_9380_18548 n3_9380_18548 0.0
V27048 n1_9380_20687 n3_9380_20687 0.0
V27049 n1_9380_20735 n3_9380_20735 0.0
V27050 n1_9380_20768 n3_9380_20768 0.0
V27051 n1_9521_215 n3_9521_215 0.0
V27052 n1_9521_248 n3_9521_248 0.0
V27053 n1_9521_383 n3_9521_383 0.0
V27054 n1_9521_431 n3_9521_431 0.0
V27055 n1_9521_647 n3_9521_647 0.0
V27056 n1_9521_680 n3_9521_680 0.0
V27057 n1_9521_863 n3_9521_863 0.0
V27058 n1_9521_896 n3_9521_896 0.0
V27059 n1_9521_1079 n3_9521_1079 0.0
V27060 n1_9521_1112 n3_9521_1112 0.0
V27061 n1_9521_1295 n3_9521_1295 0.0
V27062 n1_9521_1328 n3_9521_1328 0.0
V27063 n1_9521_1511 n3_9521_1511 0.0
V27064 n1_9521_1544 n3_9521_1544 0.0
V27065 n1_9521_1727 n3_9521_1727 0.0
V27066 n1_9521_1760 n3_9521_1760 0.0
V27067 n1_9521_1894 n3_9521_1894 0.0
V27068 n1_9521_1916 n3_9521_1916 0.0
V27069 n1_9521_1943 n3_9521_1943 0.0
V27070 n1_9521_1976 n3_9521_1976 0.0
V27071 n1_9521_2159 n3_9521_2159 0.0
V27072 n1_9521_2192 n3_9521_2192 0.0
V27073 n1_9521_2375 n3_9521_2375 0.0
V27074 n1_9521_2408 n3_9521_2408 0.0
V27075 n1_9521_2543 n3_9521_2543 0.0
V27076 n1_9521_2564 n3_9521_2564 0.0
V27077 n1_9521_2591 n3_9521_2591 0.0
V27078 n1_9521_2624 n3_9521_2624 0.0
V27079 n1_9521_2807 n3_9521_2807 0.0
V27080 n1_9521_2840 n3_9521_2840 0.0
V27081 n1_9521_2996 n3_9521_2996 0.0
V27082 n1_9521_3023 n3_9521_3023 0.0
V27083 n1_9521_3056 n3_9521_3056 0.0
V27084 n1_9521_3239 n3_9521_3239 0.0
V27085 n1_9521_3272 n3_9521_3272 0.0
V27086 n1_9521_3455 n3_9521_3455 0.0
V27087 n1_9521_3488 n3_9521_3488 0.0
V27088 n1_9521_3644 n3_9521_3644 0.0
V27089 n1_9521_3671 n3_9521_3671 0.0
V27090 n1_9521_3704 n3_9521_3704 0.0
V27091 n1_9521_3887 n3_9521_3887 0.0
V27092 n1_9521_3920 n3_9521_3920 0.0
V27093 n1_9521_4103 n3_9521_4103 0.0
V27094 n1_9521_4136 n3_9521_4136 0.0
V27095 n1_9521_4292 n3_9521_4292 0.0
V27096 n1_9521_4319 n3_9521_4319 0.0
V27097 n1_9521_4352 n3_9521_4352 0.0
V27098 n1_9521_4535 n3_9521_4535 0.0
V27099 n1_9521_4568 n3_9521_4568 0.0
V27100 n1_9521_4724 n3_9521_4724 0.0
V27101 n1_9521_4751 n3_9521_4751 0.0
V27102 n1_9521_4784 n3_9521_4784 0.0
V27103 n1_9521_5000 n3_9521_5000 0.0
V27104 n1_9521_5183 n3_9521_5183 0.0
V27105 n1_9521_5216 n3_9521_5216 0.0
V27106 n1_9521_5350 n3_9521_5350 0.0
V27107 n1_9521_5372 n3_9521_5372 0.0
V27108 n1_9521_5399 n3_9521_5399 0.0
V27109 n1_9521_5432 n3_9521_5432 0.0
V27110 n1_9521_5588 n3_9521_5588 0.0
V27111 n1_9521_5615 n3_9521_5615 0.0
V27112 n1_9521_5648 n3_9521_5648 0.0
V27113 n1_9521_5831 n3_9521_5831 0.0
V27114 n1_9521_5864 n3_9521_5864 0.0
V27115 n1_9521_6047 n3_9521_6047 0.0
V27116 n1_9521_6080 n3_9521_6080 0.0
V27117 n1_9521_6263 n3_9521_6263 0.0
V27118 n1_9521_6296 n3_9521_6296 0.0
V27119 n1_9521_6479 n3_9521_6479 0.0
V27120 n1_9521_6512 n3_9521_6512 0.0
V27121 n1_9521_6668 n3_9521_6668 0.0
V27122 n1_9521_6695 n3_9521_6695 0.0
V27123 n1_9521_6728 n3_9521_6728 0.0
V27124 n1_9521_6911 n3_9521_6911 0.0
V27125 n1_9521_6944 n3_9521_6944 0.0
V27126 n1_9521_7100 n3_9521_7100 0.0
V27127 n1_9521_7127 n3_9521_7127 0.0
V27128 n1_9521_7160 n3_9521_7160 0.0
V27129 n1_9521_7316 n3_9521_7316 0.0
V27130 n1_9521_7343 n3_9521_7343 0.0
V27131 n1_9521_7376 n3_9521_7376 0.0
V27132 n1_9521_7532 n3_9521_7532 0.0
V27133 n1_9521_7559 n3_9521_7559 0.0
V27134 n1_9521_7592 n3_9521_7592 0.0
V27135 n1_9521_7775 n3_9521_7775 0.0
V27136 n1_9521_7808 n3_9521_7808 0.0
V27137 n1_9521_7991 n3_9521_7991 0.0
V27138 n1_9521_8024 n3_9521_8024 0.0
V27139 n1_9521_8207 n3_9521_8207 0.0
V27140 n1_9521_8240 n3_9521_8240 0.0
V27141 n1_9521_8423 n3_9521_8423 0.0
V27142 n1_9521_8456 n3_9521_8456 0.0
V27143 n1_9521_8639 n3_9521_8639 0.0
V27144 n1_9521_8672 n3_9521_8672 0.0
V27145 n1_9521_8855 n3_9521_8855 0.0
V27146 n1_9521_8888 n3_9521_8888 0.0
V27147 n1_9521_9071 n3_9521_9071 0.0
V27148 n1_9521_9104 n3_9521_9104 0.0
V27149 n1_9521_9287 n3_9521_9287 0.0
V27150 n1_9521_9320 n3_9521_9320 0.0
V27151 n1_9521_9503 n3_9521_9503 0.0
V27152 n1_9521_9536 n3_9521_9536 0.0
V27153 n1_9521_9719 n3_9521_9719 0.0
V27154 n1_9521_9752 n3_9521_9752 0.0
V27155 n1_9521_9935 n3_9521_9935 0.0
V27156 n1_9521_9968 n3_9521_9968 0.0
V27157 n1_9521_10151 n3_9521_10151 0.0
V27158 n1_9521_10184 n3_9521_10184 0.0
V27159 n1_9521_10367 n3_9521_10367 0.0
V27160 n1_9521_10400 n3_9521_10400 0.0
V27161 n1_9521_10616 n3_9521_10616 0.0
V27162 n1_9521_10799 n3_9521_10799 0.0
V27163 n1_9521_10832 n3_9521_10832 0.0
V27164 n1_9521_11015 n3_9521_11015 0.0
V27165 n1_9521_11048 n3_9521_11048 0.0
V27166 n1_9521_11231 n3_9521_11231 0.0
V27167 n1_9521_11264 n3_9521_11264 0.0
V27168 n1_9521_11447 n3_9521_11447 0.0
V27169 n1_9521_11480 n3_9521_11480 0.0
V27170 n1_9521_11663 n3_9521_11663 0.0
V27171 n1_9521_11696 n3_9521_11696 0.0
V27172 n1_9521_11879 n3_9521_11879 0.0
V27173 n1_9521_11912 n3_9521_11912 0.0
V27174 n1_9521_12095 n3_9521_12095 0.0
V27175 n1_9521_12128 n3_9521_12128 0.0
V27176 n1_9521_12311 n3_9521_12311 0.0
V27177 n1_9521_12344 n3_9521_12344 0.0
V27178 n1_9521_12527 n3_9521_12527 0.0
V27179 n1_9521_12560 n3_9521_12560 0.0
V27180 n1_9521_12743 n3_9521_12743 0.0
V27181 n1_9521_12776 n3_9521_12776 0.0
V27182 n1_9521_12959 n3_9521_12959 0.0
V27183 n1_9521_12992 n3_9521_12992 0.0
V27184 n1_9521_13175 n3_9521_13175 0.0
V27185 n1_9521_13208 n3_9521_13208 0.0
V27186 n1_9521_13391 n3_9521_13391 0.0
V27187 n1_9521_13424 n3_9521_13424 0.0
V27188 n1_9521_13607 n3_9521_13607 0.0
V27189 n1_9521_13640 n3_9521_13640 0.0
V27190 n1_9521_13796 n3_9521_13796 0.0
V27191 n1_9521_13823 n3_9521_13823 0.0
V27192 n1_9521_13856 n3_9521_13856 0.0
V27193 n1_9521_13990 n3_9521_13990 0.0
V27194 n1_9521_14012 n3_9521_14012 0.0
V27195 n1_9521_14039 n3_9521_14039 0.0
V27196 n1_9521_14072 n3_9521_14072 0.0
V27197 n1_9521_14228 n3_9521_14228 0.0
V27198 n1_9521_14255 n3_9521_14255 0.0
V27199 n1_9521_14288 n3_9521_14288 0.0
V27200 n1_9521_14471 n3_9521_14471 0.0
V27201 n1_9521_14504 n3_9521_14504 0.0
V27202 n1_9521_14660 n3_9521_14660 0.0
V27203 n1_9521_14687 n3_9521_14687 0.0
V27204 n1_9521_14720 n3_9521_14720 0.0
V27205 n1_9521_14903 n3_9521_14903 0.0
V27206 n1_9521_14936 n3_9521_14936 0.0
V27207 n1_9521_15119 n3_9521_15119 0.0
V27208 n1_9521_15152 n3_9521_15152 0.0
V27209 n1_9521_15335 n3_9521_15335 0.0
V27210 n1_9521_15368 n3_9521_15368 0.0
V27211 n1_9521_15551 n3_9521_15551 0.0
V27212 n1_9521_15584 n3_9521_15584 0.0
V27213 n1_9521_15740 n3_9521_15740 0.0
V27214 n1_9521_15767 n3_9521_15767 0.0
V27215 n1_9521_15800 n3_9521_15800 0.0
V27216 n1_9521_15934 n3_9521_15934 0.0
V27217 n1_9521_15956 n3_9521_15956 0.0
V27218 n1_9521_15983 n3_9521_15983 0.0
V27219 n1_9521_16016 n3_9521_16016 0.0
V27220 n1_9521_16172 n3_9521_16172 0.0
V27221 n1_9521_16199 n3_9521_16199 0.0
V27222 n1_9521_16415 n3_9521_16415 0.0
V27223 n1_9521_16448 n3_9521_16448 0.0
V27224 n1_9521_16631 n3_9521_16631 0.0
V27225 n1_9521_16664 n3_9521_16664 0.0
V27226 n1_9521_16847 n3_9521_16847 0.0
V27227 n1_9521_16880 n3_9521_16880 0.0
V27228 n1_9521_17063 n3_9521_17063 0.0
V27229 n1_9521_17096 n3_9521_17096 0.0
V27230 n1_9521_17230 n3_9521_17230 0.0
V27231 n1_9521_17252 n3_9521_17252 0.0
V27232 n1_9521_17279 n3_9521_17279 0.0
V27233 n1_9521_17312 n3_9521_17312 0.0
V27234 n1_9521_17468 n3_9521_17468 0.0
V27235 n1_9521_17495 n3_9521_17495 0.0
V27236 n1_9521_17528 n3_9521_17528 0.0
V27237 n1_9521_17711 n3_9521_17711 0.0
V27238 n1_9521_17744 n3_9521_17744 0.0
V27239 n1_9521_17927 n3_9521_17927 0.0
V27240 n1_9521_17960 n3_9521_17960 0.0
V27241 n1_9521_18143 n3_9521_18143 0.0
V27242 n1_9521_18176 n3_9521_18176 0.0
V27243 n1_9521_18359 n3_9521_18359 0.0
V27244 n1_9521_18392 n3_9521_18392 0.0
V27245 n1_9521_18527 n3_9521_18527 0.0
V27246 n1_9521_18548 n3_9521_18548 0.0
V27247 n1_9521_18575 n3_9521_18575 0.0
V27248 n1_9521_18608 n3_9521_18608 0.0
V27249 n1_9521_18764 n3_9521_18764 0.0
V27250 n1_9521_18791 n3_9521_18791 0.0
V27251 n1_9521_18824 n3_9521_18824 0.0
V27252 n1_9521_19007 n3_9521_19007 0.0
V27253 n1_9521_19040 n3_9521_19040 0.0
V27254 n1_9521_19223 n3_9521_19223 0.0
V27255 n1_9521_19256 n3_9521_19256 0.0
V27256 n1_9521_19412 n3_9521_19412 0.0
V27257 n1_9521_19439 n3_9521_19439 0.0
V27258 n1_9521_19472 n3_9521_19472 0.0
V27259 n1_9521_19655 n3_9521_19655 0.0
V27260 n1_9521_19688 n3_9521_19688 0.0
V27261 n1_9521_19871 n3_9521_19871 0.0
V27262 n1_9521_19904 n3_9521_19904 0.0
V27263 n1_9521_20087 n3_9521_20087 0.0
V27264 n1_9521_20120 n3_9521_20120 0.0
V27265 n1_9521_20303 n3_9521_20303 0.0
V27266 n1_9521_20336 n3_9521_20336 0.0
V27267 n1_9521_20519 n3_9521_20519 0.0
V27268 n1_9521_20552 n3_9521_20552 0.0
V27269 n1_9521_20687 n3_9521_20687 0.0
V27270 n1_9521_20768 n3_9521_20768 0.0
V27271 n1_9521_20951 n3_9521_20951 0.0
V27272 n1_9521_20984 n3_9521_20984 0.0
V27273 n1_9614_215 n3_9614_215 0.0
V27274 n1_9614_248 n3_9614_248 0.0
V27275 n1_9614_383 n3_9614_383 0.0
V27276 n1_9614_431 n3_9614_431 0.0
V27277 n1_9614_464 n3_9614_464 0.0
V27278 n1_9614_647 n3_9614_647 0.0
V27279 n1_9614_680 n3_9614_680 0.0
V27280 n1_9614_863 n3_9614_863 0.0
V27281 n1_9614_896 n3_9614_896 0.0
V27282 n1_9614_1079 n3_9614_1079 0.0
V27283 n1_9614_1112 n3_9614_1112 0.0
V27284 n1_9614_1295 n3_9614_1295 0.0
V27285 n1_9614_1328 n3_9614_1328 0.0
V27286 n1_9614_1511 n3_9614_1511 0.0
V27287 n1_9614_1544 n3_9614_1544 0.0
V27288 n1_9614_1727 n3_9614_1727 0.0
V27289 n1_9614_1760 n3_9614_1760 0.0
V27290 n1_9614_1916 n3_9614_1916 0.0
V27291 n1_9614_1943 n3_9614_1943 0.0
V27292 n1_9614_1976 n3_9614_1976 0.0
V27293 n1_9614_2159 n3_9614_2159 0.0
V27294 n1_9614_2192 n3_9614_2192 0.0
V27295 n1_9614_2375 n3_9614_2375 0.0
V27296 n1_9614_2408 n3_9614_2408 0.0
V27297 n1_9614_2543 n3_9614_2543 0.0
V27298 n1_9614_2564 n3_9614_2564 0.0
V27299 n1_9614_2591 n3_9614_2591 0.0
V27300 n1_9614_2624 n3_9614_2624 0.0
V27301 n1_9614_18527 n3_9614_18527 0.0
V27302 n1_9614_18548 n3_9614_18548 0.0
V27303 n1_9614_18575 n3_9614_18575 0.0
V27304 n1_9614_18608 n3_9614_18608 0.0
V27305 n1_9614_18764 n3_9614_18764 0.0
V27306 n1_9614_18791 n3_9614_18791 0.0
V27307 n1_9614_18824 n3_9614_18824 0.0
V27308 n1_9614_19007 n3_9614_19007 0.0
V27309 n1_9614_19040 n3_9614_19040 0.0
V27310 n1_9614_19223 n3_9614_19223 0.0
V27311 n1_9614_19256 n3_9614_19256 0.0
V27312 n1_9614_19412 n3_9614_19412 0.0
V27313 n1_9614_19439 n3_9614_19439 0.0
V27314 n1_9614_19472 n3_9614_19472 0.0
V27315 n1_9614_19655 n3_9614_19655 0.0
V27316 n1_9614_19688 n3_9614_19688 0.0
V27317 n1_9614_19871 n3_9614_19871 0.0
V27318 n1_9614_19904 n3_9614_19904 0.0
V27319 n1_9614_20087 n3_9614_20087 0.0
V27320 n1_9614_20120 n3_9614_20120 0.0
V27321 n1_9614_20303 n3_9614_20303 0.0
V27322 n1_9614_20336 n3_9614_20336 0.0
V27323 n1_9614_20519 n3_9614_20519 0.0
V27324 n1_9614_20552 n3_9614_20552 0.0
V27325 n1_9614_20687 n3_9614_20687 0.0
V27326 n1_9614_20735 n3_9614_20735 0.0
V27327 n1_9614_20768 n3_9614_20768 0.0
V27328 n1_9614_20951 n3_9614_20951 0.0
V27329 n1_9614_20984 n3_9614_20984 0.0
V27330 n1_11400_215 n3_11400_215 0.0
V27331 n1_11400_248 n3_11400_248 0.0
V27332 n1_11400_383 n3_11400_383 0.0
V27333 n1_11400_431 n3_11400_431 0.0
V27334 n1_11400_464 n3_11400_464 0.0
V27335 n1_11400_647 n3_11400_647 0.0
V27336 n1_11400_680 n3_11400_680 0.0
V27337 n1_11400_863 n3_11400_863 0.0
V27338 n1_11400_896 n3_11400_896 0.0
V27339 n1_11400_1079 n3_11400_1079 0.0
V27340 n1_11400_1112 n3_11400_1112 0.0
V27341 n1_11400_1295 n3_11400_1295 0.0
V27342 n1_11400_1328 n3_11400_1328 0.0
V27343 n1_11400_1511 n3_11400_1511 0.0
V27344 n1_11400_1544 n3_11400_1544 0.0
V27345 n1_11400_1727 n3_11400_1727 0.0
V27346 n1_11400_1760 n3_11400_1760 0.0
V27347 n1_11400_1894 n3_11400_1894 0.0
V27348 n1_11400_1943 n3_11400_1943 0.0
V27349 n1_11400_1976 n3_11400_1976 0.0
V27350 n1_11400_2159 n3_11400_2159 0.0
V27351 n1_11400_2192 n3_11400_2192 0.0
V27352 n1_11400_2375 n3_11400_2375 0.0
V27353 n1_11400_2408 n3_11400_2408 0.0
V27354 n1_11400_2543 n3_11400_2543 0.0
V27355 n1_11400_2591 n3_11400_2591 0.0
V27356 n1_11400_2624 n3_11400_2624 0.0
V27357 n1_11400_18527 n3_11400_18527 0.0
V27358 n1_11400_18548 n3_11400_18548 0.0
V27359 n1_11400_18575 n3_11400_18575 0.0
V27360 n1_11400_18608 n3_11400_18608 0.0
V27361 n1_11400_18764 n3_11400_18764 0.0
V27362 n1_11400_18791 n3_11400_18791 0.0
V27363 n1_11400_18824 n3_11400_18824 0.0
V27364 n1_11400_19007 n3_11400_19007 0.0
V27365 n1_11400_19040 n3_11400_19040 0.0
V27366 n1_11400_19223 n3_11400_19223 0.0
V27367 n1_11400_19256 n3_11400_19256 0.0
V27368 n1_11400_19412 n3_11400_19412 0.0
V27369 n1_11400_19439 n3_11400_19439 0.0
V27370 n1_11400_19472 n3_11400_19472 0.0
V27371 n1_11400_19655 n3_11400_19655 0.0
V27372 n1_11400_19688 n3_11400_19688 0.0
V27373 n1_11400_19871 n3_11400_19871 0.0
V27374 n1_11400_19904 n3_11400_19904 0.0
V27375 n1_11400_20087 n3_11400_20087 0.0
V27376 n1_11400_20120 n3_11400_20120 0.0
V27377 n1_11400_20303 n3_11400_20303 0.0
V27378 n1_11400_20336 n3_11400_20336 0.0
V27379 n1_11400_20519 n3_11400_20519 0.0
V27380 n1_11400_20552 n3_11400_20552 0.0
V27381 n1_11400_20687 n3_11400_20687 0.0
V27382 n1_11400_20735 n3_11400_20735 0.0
V27383 n1_11400_20768 n3_11400_20768 0.0
V27384 n1_11400_20951 n3_11400_20951 0.0
V27385 n1_11400_20984 n3_11400_20984 0.0
V27386 n1_11583_215 n3_11583_215 0.0
V27387 n1_11583_248 n3_11583_248 0.0
V27388 n1_11583_383 n3_11583_383 0.0
V27389 n1_11583_431 n3_11583_431 0.0
V27390 n1_11583_464 n3_11583_464 0.0
V27391 n1_11583_647 n3_11583_647 0.0
V27392 n1_11583_680 n3_11583_680 0.0
V27393 n1_11583_863 n3_11583_863 0.0
V27394 n1_11583_896 n3_11583_896 0.0
V27395 n1_11583_1079 n3_11583_1079 0.0
V27396 n1_11583_1112 n3_11583_1112 0.0
V27397 n1_11583_1295 n3_11583_1295 0.0
V27398 n1_11583_1328 n3_11583_1328 0.0
V27399 n1_11583_1727 n3_11583_1727 0.0
V27400 n1_11583_1760 n3_11583_1760 0.0
V27401 n1_11583_1894 n3_11583_1894 0.0
V27402 n1_11583_1943 n3_11583_1943 0.0
V27403 n1_11583_1976 n3_11583_1976 0.0
V27404 n1_11583_2159 n3_11583_2159 0.0
V27405 n1_11583_2192 n3_11583_2192 0.0
V27406 n1_11583_2375 n3_11583_2375 0.0
V27407 n1_11583_2408 n3_11583_2408 0.0
V27408 n1_11583_2542 n3_11583_2542 0.0
V27409 n1_11583_2543 n3_11583_2543 0.0
V27410 n1_11583_2591 n3_11583_2591 0.0
V27411 n1_11583_2624 n3_11583_2624 0.0
V27412 n1_11583_2760 n3_11583_2760 0.0
V27413 n1_11583_2807 n3_11583_2807 0.0
V27414 n1_11583_2840 n3_11583_2840 0.0
V27415 n1_11583_2974 n3_11583_2974 0.0
V27416 n1_11583_3023 n3_11583_3023 0.0
V27417 n1_11583_3056 n3_11583_3056 0.0
V27418 n1_11583_3239 n3_11583_3239 0.0
V27419 n1_11583_3272 n3_11583_3272 0.0
V27420 n1_11583_3455 n3_11583_3455 0.0
V27421 n1_11583_3488 n3_11583_3488 0.0
V27422 n1_11583_3622 n3_11583_3622 0.0
V27423 n1_11583_3671 n3_11583_3671 0.0
V27424 n1_11583_3704 n3_11583_3704 0.0
V27425 n1_11583_4103 n3_11583_4103 0.0
V27426 n1_11583_4136 n3_11583_4136 0.0
V27427 n1_11583_4270 n3_11583_4270 0.0
V27428 n1_11583_4319 n3_11583_4319 0.0
V27429 n1_11583_4352 n3_11583_4352 0.0
V27430 n1_11583_4535 n3_11583_4535 0.0
V27431 n1_11583_4568 n3_11583_4568 0.0
V27432 n1_11583_4702 n3_11583_4702 0.0
V27433 n1_11583_4751 n3_11583_4751 0.0
V27434 n1_11583_4784 n3_11583_4784 0.0
V27435 n1_11583_4967 n3_11583_4967 0.0
V27436 n1_11583_5000 n3_11583_5000 0.0
V27437 n1_11583_5183 n3_11583_5183 0.0
V27438 n1_11583_5216 n3_11583_5216 0.0
V27439 n1_11583_5350 n3_11583_5350 0.0
V27440 n1_11583_5399 n3_11583_5399 0.0
V27441 n1_11583_5432 n3_11583_5432 0.0
V27442 n1_11583_5566 n3_11583_5566 0.0
V27443 n1_11583_5615 n3_11583_5615 0.0
V27444 n1_11583_5648 n3_11583_5648 0.0
V27445 n1_11583_5782 n3_11583_5782 0.0
V27446 n1_11583_5831 n3_11583_5831 0.0
V27447 n1_11583_5864 n3_11583_5864 0.0
V27448 n1_11583_6263 n3_11583_6263 0.0
V27449 n1_11583_6296 n3_11583_6296 0.0
V27450 n1_11583_6430 n3_11583_6430 0.0
V27451 n1_11583_6479 n3_11583_6479 0.0
V27452 n1_11583_6512 n3_11583_6512 0.0
V27453 n1_11583_6646 n3_11583_6646 0.0
V27454 n1_11583_6695 n3_11583_6695 0.0
V27455 n1_11583_6728 n3_11583_6728 0.0
V27456 n1_11583_6862 n3_11583_6862 0.0
V27457 n1_11583_6911 n3_11583_6911 0.0
V27458 n1_11583_6944 n3_11583_6944 0.0
V27459 n1_11583_7078 n3_11583_7078 0.0
V27460 n1_11583_7127 n3_11583_7127 0.0
V27461 n1_11583_7160 n3_11583_7160 0.0
V27462 n1_11583_7294 n3_11583_7294 0.0
V27463 n1_11583_7343 n3_11583_7343 0.0
V27464 n1_11583_7376 n3_11583_7376 0.0
V27465 n1_11583_7510 n3_11583_7510 0.0
V27466 n1_11583_7559 n3_11583_7559 0.0
V27467 n1_11583_7592 n3_11583_7592 0.0
V27468 n1_11583_7775 n3_11583_7775 0.0
V27469 n1_11583_7808 n3_11583_7808 0.0
V27470 n1_11583_7991 n3_11583_7991 0.0
V27471 n1_11583_8024 n3_11583_8024 0.0
V27472 n1_11583_8207 n3_11583_8207 0.0
V27473 n1_11583_8240 n3_11583_8240 0.0
V27474 n1_11583_8456 n3_11583_8456 0.0
V27475 n1_11583_8639 n3_11583_8639 0.0
V27476 n1_11583_8672 n3_11583_8672 0.0
V27477 n1_11583_8855 n3_11583_8855 0.0
V27478 n1_11583_8888 n3_11583_8888 0.0
V27479 n1_11583_9071 n3_11583_9071 0.0
V27480 n1_11583_9104 n3_11583_9104 0.0
V27481 n1_11583_9287 n3_11583_9287 0.0
V27482 n1_11583_9320 n3_11583_9320 0.0
V27483 n1_11583_9503 n3_11583_9503 0.0
V27484 n1_11583_9536 n3_11583_9536 0.0
V27485 n1_11583_9719 n3_11583_9719 0.0
V27486 n1_11583_9752 n3_11583_9752 0.0
V27487 n1_11583_9935 n3_11583_9935 0.0
V27488 n1_11583_9968 n3_11583_9968 0.0
V27489 n1_11583_10151 n3_11583_10151 0.0
V27490 n1_11583_10184 n3_11583_10184 0.0
V27491 n1_11583_10367 n3_11583_10367 0.0
V27492 n1_11583_10400 n3_11583_10400 0.0
V27493 n1_11583_10799 n3_11583_10799 0.0
V27494 n1_11583_10832 n3_11583_10832 0.0
V27495 n1_11583_11015 n3_11583_11015 0.0
V27496 n1_11583_11048 n3_11583_11048 0.0
V27497 n1_11583_11231 n3_11583_11231 0.0
V27498 n1_11583_11264 n3_11583_11264 0.0
V27499 n1_11583_11447 n3_11583_11447 0.0
V27500 n1_11583_11480 n3_11583_11480 0.0
V27501 n1_11583_11663 n3_11583_11663 0.0
V27502 n1_11583_11696 n3_11583_11696 0.0
V27503 n1_11583_11879 n3_11583_11879 0.0
V27504 n1_11583_11912 n3_11583_11912 0.0
V27505 n1_11583_12095 n3_11583_12095 0.0
V27506 n1_11583_12128 n3_11583_12128 0.0
V27507 n1_11583_12311 n3_11583_12311 0.0
V27508 n1_11583_12344 n3_11583_12344 0.0
V27509 n1_11583_12527 n3_11583_12527 0.0
V27510 n1_11583_12560 n3_11583_12560 0.0
V27511 n1_11583_12743 n3_11583_12743 0.0
V27512 n1_11583_12959 n3_11583_12959 0.0
V27513 n1_11583_12992 n3_11583_12992 0.0
V27514 n1_11583_13175 n3_11583_13175 0.0
V27515 n1_11583_13208 n3_11583_13208 0.0
V27516 n1_11583_13391 n3_11583_13391 0.0
V27517 n1_11583_13424 n3_11583_13424 0.0
V27518 n1_11583_13607 n3_11583_13607 0.0
V27519 n1_11583_13640 n3_11583_13640 0.0
V27520 n1_11583_13774 n3_11583_13774 0.0
V27521 n1_11583_13823 n3_11583_13823 0.0
V27522 n1_11583_13856 n3_11583_13856 0.0
V27523 n1_11583_14012 n3_11583_14012 0.0
V27524 n1_11583_14039 n3_11583_14039 0.0
V27525 n1_11583_14072 n3_11583_14072 0.0
V27526 n1_11583_14220 n3_11583_14220 0.0
V27527 n1_11583_14255 n3_11583_14255 0.0
V27528 n1_11583_14288 n3_11583_14288 0.0
V27529 n1_11583_14471 n3_11583_14471 0.0
V27530 n1_11583_14504 n3_11583_14504 0.0
V27531 n1_11583_14660 n3_11583_14660 0.0
V27532 n1_11583_14687 n3_11583_14687 0.0
V27533 n1_11583_14720 n3_11583_14720 0.0
V27534 n1_11583_14903 n3_11583_14903 0.0
V27535 n1_11583_14936 n3_11583_14936 0.0
V27536 n1_11583_15335 n3_11583_15335 0.0
V27537 n1_11583_15368 n3_11583_15368 0.0
V27538 n1_11583_15551 n3_11583_15551 0.0
V27539 n1_11583_15584 n3_11583_15584 0.0
V27540 n1_11583_15740 n3_11583_15740 0.0
V27541 n1_11583_15767 n3_11583_15767 0.0
V27542 n1_11583_15800 n3_11583_15800 0.0
V27543 n1_11583_15948 n3_11583_15948 0.0
V27544 n1_11583_15956 n3_11583_15956 0.0
V27545 n1_11583_15983 n3_11583_15983 0.0
V27546 n1_11583_16016 n3_11583_16016 0.0
V27547 n1_11583_16172 n3_11583_16172 0.0
V27548 n1_11583_16199 n3_11583_16199 0.0
V27549 n1_11583_16232 n3_11583_16232 0.0
V27550 n1_11583_16415 n3_11583_16415 0.0
V27551 n1_11583_16448 n3_11583_16448 0.0
V27552 n1_11583_16604 n3_11583_16604 0.0
V27553 n1_11583_16631 n3_11583_16631 0.0
V27554 n1_11583_16664 n3_11583_16664 0.0
V27555 n1_11583_16847 n3_11583_16847 0.0
V27556 n1_11583_16880 n3_11583_16880 0.0
V27557 n1_11583_17063 n3_11583_17063 0.0
V27558 n1_11583_17096 n3_11583_17096 0.0
V27559 n1_11583_17244 n3_11583_17244 0.0
V27560 n1_11583_17468 n3_11583_17468 0.0
V27561 n1_11583_17495 n3_11583_17495 0.0
V27562 n1_11583_17528 n3_11583_17528 0.0
V27563 n1_11583_17684 n3_11583_17684 0.0
V27564 n1_11583_17711 n3_11583_17711 0.0
V27565 n1_11583_17744 n3_11583_17744 0.0
V27566 n1_11583_17927 n3_11583_17927 0.0
V27567 n1_11583_17960 n3_11583_17960 0.0
V27568 n1_11583_18143 n3_11583_18143 0.0
V27569 n1_11583_18176 n3_11583_18176 0.0
V27570 n1_11583_18332 n3_11583_18332 0.0
V27571 n1_11583_18359 n3_11583_18359 0.0
V27572 n1_11583_18392 n3_11583_18392 0.0
V27573 n1_11583_18527 n3_11583_18527 0.0
V27574 n1_11583_18548 n3_11583_18548 0.0
V27575 n1_11583_18575 n3_11583_18575 0.0
V27576 n1_11583_18608 n3_11583_18608 0.0
V27577 n1_11583_18764 n3_11583_18764 0.0
V27578 n1_11583_18791 n3_11583_18791 0.0
V27579 n1_11583_18824 n3_11583_18824 0.0
V27580 n1_11583_19007 n3_11583_19007 0.0
V27581 n1_11583_19040 n3_11583_19040 0.0
V27582 n1_11583_19223 n3_11583_19223 0.0
V27583 n1_11583_19256 n3_11583_19256 0.0
V27584 n1_11583_19404 n3_11583_19404 0.0
V27585 n1_11583_19412 n3_11583_19412 0.0
V27586 n1_11583_19439 n3_11583_19439 0.0
V27587 n1_11583_19472 n3_11583_19472 0.0
V27588 n1_11583_19871 n3_11583_19871 0.0
V27589 n1_11583_19904 n3_11583_19904 0.0
V27590 n1_11583_20087 n3_11583_20087 0.0
V27591 n1_11583_20120 n3_11583_20120 0.0
V27592 n1_11583_20303 n3_11583_20303 0.0
V27593 n1_11583_20336 n3_11583_20336 0.0
V27594 n1_11583_20519 n3_11583_20519 0.0
V27595 n1_11583_20552 n3_11583_20552 0.0
V27596 n1_11583_20687 n3_11583_20687 0.0
V27597 n1_11583_20735 n3_11583_20735 0.0
V27598 n1_11583_20768 n3_11583_20768 0.0
V27599 n1_11583_20951 n3_11583_20951 0.0
V27600 n1_11583_20984 n3_11583_20984 0.0
V27601 n1_11630_431 n3_11630_431 0.0
V27602 n1_11630_464 n3_11630_464 0.0
V27603 n1_11630_2760 n3_11630_2760 0.0
V27604 n1_11630_4967 n3_11630_4967 0.0
V27605 n1_11630_5000 n3_11630_5000 0.0
V27606 n1_11630_7160 n3_11630_7160 0.0
V27607 n1_11630_7294 n3_11630_7294 0.0
V27608 n1_11630_9503 n3_11630_9503 0.0
V27609 n1_11630_9536 n3_11630_9536 0.0
V27610 n1_11630_11663 n3_11630_11663 0.0
V27611 n1_11630_11696 n3_11630_11696 0.0
V27612 n1_11630_14012 n3_11630_14012 0.0
V27613 n1_11630_14039 n3_11630_14039 0.0
V27614 n1_11630_16172 n3_11630_16172 0.0
V27615 n1_11630_16199 n3_11630_16199 0.0
V27616 n1_11630_16232 n3_11630_16232 0.0
V27617 n1_11630_18392 n3_11630_18392 0.0
V27618 n1_11630_18527 n3_11630_18527 0.0
V27619 n1_11630_18548 n3_11630_18548 0.0
V27620 n1_11630_20687 n3_11630_20687 0.0
V27621 n1_11630_20735 n3_11630_20735 0.0
V27622 n1_11630_20768 n3_11630_20768 0.0
V27623 n1_11771_215 n3_11771_215 0.0
V27624 n1_11771_248 n3_11771_248 0.0
V27625 n1_11771_383 n3_11771_383 0.0
V27626 n1_11771_431 n3_11771_431 0.0
V27627 n1_11771_647 n3_11771_647 0.0
V27628 n1_11771_680 n3_11771_680 0.0
V27629 n1_11771_863 n3_11771_863 0.0
V27630 n1_11771_896 n3_11771_896 0.0
V27631 n1_11771_1079 n3_11771_1079 0.0
V27632 n1_11771_1112 n3_11771_1112 0.0
V27633 n1_11771_1295 n3_11771_1295 0.0
V27634 n1_11771_1328 n3_11771_1328 0.0
V27635 n1_11771_1511 n3_11771_1511 0.0
V27636 n1_11771_1544 n3_11771_1544 0.0
V27637 n1_11771_1727 n3_11771_1727 0.0
V27638 n1_11771_1760 n3_11771_1760 0.0
V27639 n1_11771_1894 n3_11771_1894 0.0
V27640 n1_11771_1943 n3_11771_1943 0.0
V27641 n1_11771_1976 n3_11771_1976 0.0
V27642 n1_11771_2159 n3_11771_2159 0.0
V27643 n1_11771_2192 n3_11771_2192 0.0
V27644 n1_11771_2375 n3_11771_2375 0.0
V27645 n1_11771_2408 n3_11771_2408 0.0
V27646 n1_11771_2542 n3_11771_2542 0.0
V27647 n1_11771_2543 n3_11771_2543 0.0
V27648 n1_11771_2591 n3_11771_2591 0.0
V27649 n1_11771_2624 n3_11771_2624 0.0
V27650 n1_11771_2760 n3_11771_2760 0.0
V27651 n1_11771_2807 n3_11771_2807 0.0
V27652 n1_11771_2840 n3_11771_2840 0.0
V27653 n1_11771_2974 n3_11771_2974 0.0
V27654 n1_11771_3023 n3_11771_3023 0.0
V27655 n1_11771_3056 n3_11771_3056 0.0
V27656 n1_11771_3239 n3_11771_3239 0.0
V27657 n1_11771_3272 n3_11771_3272 0.0
V27658 n1_11771_3455 n3_11771_3455 0.0
V27659 n1_11771_3488 n3_11771_3488 0.0
V27660 n1_11771_3622 n3_11771_3622 0.0
V27661 n1_11771_3671 n3_11771_3671 0.0
V27662 n1_11771_3704 n3_11771_3704 0.0
V27663 n1_11771_3887 n3_11771_3887 0.0
V27664 n1_11771_3920 n3_11771_3920 0.0
V27665 n1_11771_4103 n3_11771_4103 0.0
V27666 n1_11771_4136 n3_11771_4136 0.0
V27667 n1_11771_4270 n3_11771_4270 0.0
V27668 n1_11771_4319 n3_11771_4319 0.0
V27669 n1_11771_4352 n3_11771_4352 0.0
V27670 n1_11771_4535 n3_11771_4535 0.0
V27671 n1_11771_4568 n3_11771_4568 0.0
V27672 n1_11771_4702 n3_11771_4702 0.0
V27673 n1_11771_4751 n3_11771_4751 0.0
V27674 n1_11771_4784 n3_11771_4784 0.0
V27675 n1_11771_5000 n3_11771_5000 0.0
V27676 n1_11771_5183 n3_11771_5183 0.0
V27677 n1_11771_5216 n3_11771_5216 0.0
V27678 n1_11771_5350 n3_11771_5350 0.0
V27679 n1_11771_5399 n3_11771_5399 0.0
V27680 n1_11771_5432 n3_11771_5432 0.0
V27681 n1_11771_5566 n3_11771_5566 0.0
V27682 n1_11771_5615 n3_11771_5615 0.0
V27683 n1_11771_5648 n3_11771_5648 0.0
V27684 n1_11771_5782 n3_11771_5782 0.0
V27685 n1_11771_5831 n3_11771_5831 0.0
V27686 n1_11771_5864 n3_11771_5864 0.0
V27687 n1_11771_6047 n3_11771_6047 0.0
V27688 n1_11771_6080 n3_11771_6080 0.0
V27689 n1_11771_6263 n3_11771_6263 0.0
V27690 n1_11771_6296 n3_11771_6296 0.0
V27691 n1_11771_6430 n3_11771_6430 0.0
V27692 n1_11771_6479 n3_11771_6479 0.0
V27693 n1_11771_6512 n3_11771_6512 0.0
V27694 n1_11771_6646 n3_11771_6646 0.0
V27695 n1_11771_6695 n3_11771_6695 0.0
V27696 n1_11771_6728 n3_11771_6728 0.0
V27697 n1_11771_6862 n3_11771_6862 0.0
V27698 n1_11771_6911 n3_11771_6911 0.0
V27699 n1_11771_6944 n3_11771_6944 0.0
V27700 n1_11771_7078 n3_11771_7078 0.0
V27701 n1_11771_7127 n3_11771_7127 0.0
V27702 n1_11771_7160 n3_11771_7160 0.0
V27703 n1_11771_7294 n3_11771_7294 0.0
V27704 n1_11771_7343 n3_11771_7343 0.0
V27705 n1_11771_7376 n3_11771_7376 0.0
V27706 n1_11771_7510 n3_11771_7510 0.0
V27707 n1_11771_7559 n3_11771_7559 0.0
V27708 n1_11771_7592 n3_11771_7592 0.0
V27709 n1_11771_7775 n3_11771_7775 0.0
V27710 n1_11771_7808 n3_11771_7808 0.0
V27711 n1_11771_7991 n3_11771_7991 0.0
V27712 n1_11771_8024 n3_11771_8024 0.0
V27713 n1_11771_8207 n3_11771_8207 0.0
V27714 n1_11771_8240 n3_11771_8240 0.0
V27715 n1_11771_8423 n3_11771_8423 0.0
V27716 n1_11771_8456 n3_11771_8456 0.0
V27717 n1_11771_8639 n3_11771_8639 0.0
V27718 n1_11771_8672 n3_11771_8672 0.0
V27719 n1_11771_8855 n3_11771_8855 0.0
V27720 n1_11771_8888 n3_11771_8888 0.0
V27721 n1_11771_9071 n3_11771_9071 0.0
V27722 n1_11771_9104 n3_11771_9104 0.0
V27723 n1_11771_9287 n3_11771_9287 0.0
V27724 n1_11771_9320 n3_11771_9320 0.0
V27725 n1_11771_9503 n3_11771_9503 0.0
V27726 n1_11771_9536 n3_11771_9536 0.0
V27727 n1_11771_9719 n3_11771_9719 0.0
V27728 n1_11771_9752 n3_11771_9752 0.0
V27729 n1_11771_9935 n3_11771_9935 0.0
V27730 n1_11771_9968 n3_11771_9968 0.0
V27731 n1_11771_10151 n3_11771_10151 0.0
V27732 n1_11771_10184 n3_11771_10184 0.0
V27733 n1_11771_10367 n3_11771_10367 0.0
V27734 n1_11771_10400 n3_11771_10400 0.0
V27735 n1_11771_10616 n3_11771_10616 0.0
V27736 n1_11771_10799 n3_11771_10799 0.0
V27737 n1_11771_10832 n3_11771_10832 0.0
V27738 n1_11771_11015 n3_11771_11015 0.0
V27739 n1_11771_11048 n3_11771_11048 0.0
V27740 n1_11771_11231 n3_11771_11231 0.0
V27741 n1_11771_11264 n3_11771_11264 0.0
V27742 n1_11771_11447 n3_11771_11447 0.0
V27743 n1_11771_11480 n3_11771_11480 0.0
V27744 n1_11771_11663 n3_11771_11663 0.0
V27745 n1_11771_11696 n3_11771_11696 0.0
V27746 n1_11771_11879 n3_11771_11879 0.0
V27747 n1_11771_11912 n3_11771_11912 0.0
V27748 n1_11771_12095 n3_11771_12095 0.0
V27749 n1_11771_12128 n3_11771_12128 0.0
V27750 n1_11771_12311 n3_11771_12311 0.0
V27751 n1_11771_12344 n3_11771_12344 0.0
V27752 n1_11771_12527 n3_11771_12527 0.0
V27753 n1_11771_12560 n3_11771_12560 0.0
V27754 n1_11771_12743 n3_11771_12743 0.0
V27755 n1_11771_12776 n3_11771_12776 0.0
V27756 n1_11771_12959 n3_11771_12959 0.0
V27757 n1_11771_12992 n3_11771_12992 0.0
V27758 n1_11771_13175 n3_11771_13175 0.0
V27759 n1_11771_13208 n3_11771_13208 0.0
V27760 n1_11771_13391 n3_11771_13391 0.0
V27761 n1_11771_13424 n3_11771_13424 0.0
V27762 n1_11771_13607 n3_11771_13607 0.0
V27763 n1_11771_13640 n3_11771_13640 0.0
V27764 n1_11771_13774 n3_11771_13774 0.0
V27765 n1_11771_13823 n3_11771_13823 0.0
V27766 n1_11771_13856 n3_11771_13856 0.0
V27767 n1_11771_14012 n3_11771_14012 0.0
V27768 n1_11771_14039 n3_11771_14039 0.0
V27769 n1_11771_14072 n3_11771_14072 0.0
V27770 n1_11771_14220 n3_11771_14220 0.0
V27771 n1_11771_14255 n3_11771_14255 0.0
V27772 n1_11771_14288 n3_11771_14288 0.0
V27773 n1_11771_14471 n3_11771_14471 0.0
V27774 n1_11771_14504 n3_11771_14504 0.0
V27775 n1_11771_14660 n3_11771_14660 0.0
V27776 n1_11771_14687 n3_11771_14687 0.0
V27777 n1_11771_14720 n3_11771_14720 0.0
V27778 n1_11771_14903 n3_11771_14903 0.0
V27779 n1_11771_14936 n3_11771_14936 0.0
V27780 n1_11771_15119 n3_11771_15119 0.0
V27781 n1_11771_15152 n3_11771_15152 0.0
V27782 n1_11771_15335 n3_11771_15335 0.0
V27783 n1_11771_15368 n3_11771_15368 0.0
V27784 n1_11771_15551 n3_11771_15551 0.0
V27785 n1_11771_15584 n3_11771_15584 0.0
V27786 n1_11771_15740 n3_11771_15740 0.0
V27787 n1_11771_15767 n3_11771_15767 0.0
V27788 n1_11771_15800 n3_11771_15800 0.0
V27789 n1_11771_15948 n3_11771_15948 0.0
V27790 n1_11771_15956 n3_11771_15956 0.0
V27791 n1_11771_15983 n3_11771_15983 0.0
V27792 n1_11771_16016 n3_11771_16016 0.0
V27793 n1_11771_16172 n3_11771_16172 0.0
V27794 n1_11771_16199 n3_11771_16199 0.0
V27795 n1_11771_16415 n3_11771_16415 0.0
V27796 n1_11771_16448 n3_11771_16448 0.0
V27797 n1_11771_16604 n3_11771_16604 0.0
V27798 n1_11771_16631 n3_11771_16631 0.0
V27799 n1_11771_16664 n3_11771_16664 0.0
V27800 n1_11771_16847 n3_11771_16847 0.0
V27801 n1_11771_16880 n3_11771_16880 0.0
V27802 n1_11771_17063 n3_11771_17063 0.0
V27803 n1_11771_17096 n3_11771_17096 0.0
V27804 n1_11771_17244 n3_11771_17244 0.0
V27805 n1_11771_17279 n3_11771_17279 0.0
V27806 n1_11771_17312 n3_11771_17312 0.0
V27807 n1_11771_17468 n3_11771_17468 0.0
V27808 n1_11771_17495 n3_11771_17495 0.0
V27809 n1_11771_17528 n3_11771_17528 0.0
V27810 n1_11771_17684 n3_11771_17684 0.0
V27811 n1_11771_17711 n3_11771_17711 0.0
V27812 n1_11771_17744 n3_11771_17744 0.0
V27813 n1_11771_17927 n3_11771_17927 0.0
V27814 n1_11771_17960 n3_11771_17960 0.0
V27815 n1_11771_18143 n3_11771_18143 0.0
V27816 n1_11771_18176 n3_11771_18176 0.0
V27817 n1_11771_18332 n3_11771_18332 0.0
V27818 n1_11771_18359 n3_11771_18359 0.0
V27819 n1_11771_18392 n3_11771_18392 0.0
V27820 n1_11771_18527 n3_11771_18527 0.0
V27821 n1_11771_18548 n3_11771_18548 0.0
V27822 n1_11771_18575 n3_11771_18575 0.0
V27823 n1_11771_18608 n3_11771_18608 0.0
V27824 n1_11771_18764 n3_11771_18764 0.0
V27825 n1_11771_18791 n3_11771_18791 0.0
V27826 n1_11771_18824 n3_11771_18824 0.0
V27827 n1_11771_19007 n3_11771_19007 0.0
V27828 n1_11771_19040 n3_11771_19040 0.0
V27829 n1_11771_19223 n3_11771_19223 0.0
V27830 n1_11771_19256 n3_11771_19256 0.0
V27831 n1_11771_19404 n3_11771_19404 0.0
V27832 n1_11771_19412 n3_11771_19412 0.0
V27833 n1_11771_19439 n3_11771_19439 0.0
V27834 n1_11771_19472 n3_11771_19472 0.0
V27835 n1_11771_19655 n3_11771_19655 0.0
V27836 n1_11771_19688 n3_11771_19688 0.0
V27837 n1_11771_19871 n3_11771_19871 0.0
V27838 n1_11771_19904 n3_11771_19904 0.0
V27839 n1_11771_20087 n3_11771_20087 0.0
V27840 n1_11771_20120 n3_11771_20120 0.0
V27841 n1_11771_20303 n3_11771_20303 0.0
V27842 n1_11771_20336 n3_11771_20336 0.0
V27843 n1_11771_20519 n3_11771_20519 0.0
V27844 n1_11771_20552 n3_11771_20552 0.0
V27845 n1_11771_20687 n3_11771_20687 0.0
V27846 n1_11771_20768 n3_11771_20768 0.0
V27847 n1_11771_20951 n3_11771_20951 0.0
V27848 n1_11771_20984 n3_11771_20984 0.0
V27849 n1_11864_215 n3_11864_215 0.0
V27850 n1_11864_248 n3_11864_248 0.0
V27851 n1_11864_383 n3_11864_383 0.0
V27852 n1_11864_431 n3_11864_431 0.0
V27853 n1_11864_464 n3_11864_464 0.0
V27854 n1_11864_647 n3_11864_647 0.0
V27855 n1_11864_680 n3_11864_680 0.0
V27856 n1_11864_863 n3_11864_863 0.0
V27857 n1_11864_896 n3_11864_896 0.0
V27858 n1_11864_1079 n3_11864_1079 0.0
V27859 n1_11864_1112 n3_11864_1112 0.0
V27860 n1_11864_1295 n3_11864_1295 0.0
V27861 n1_11864_1328 n3_11864_1328 0.0
V27862 n1_11864_1511 n3_11864_1511 0.0
V27863 n1_11864_1544 n3_11864_1544 0.0
V27864 n1_11864_1727 n3_11864_1727 0.0
V27865 n1_11864_1760 n3_11864_1760 0.0
V27866 n1_11864_1894 n3_11864_1894 0.0
V27867 n1_11864_1943 n3_11864_1943 0.0
V27868 n1_11864_1976 n3_11864_1976 0.0
V27869 n1_11864_2159 n3_11864_2159 0.0
V27870 n1_11864_2192 n3_11864_2192 0.0
V27871 n1_11864_2375 n3_11864_2375 0.0
V27872 n1_11864_2408 n3_11864_2408 0.0
V27873 n1_11864_2542 n3_11864_2542 0.0
V27874 n1_11864_2543 n3_11864_2543 0.0
V27875 n1_11864_2591 n3_11864_2591 0.0
V27876 n1_11864_2624 n3_11864_2624 0.0
V27877 n1_11864_18527 n3_11864_18527 0.0
V27878 n1_11864_18575 n3_11864_18575 0.0
V27879 n1_11864_18608 n3_11864_18608 0.0
V27880 n1_11864_18764 n3_11864_18764 0.0
V27881 n1_11864_18791 n3_11864_18791 0.0
V27882 n1_11864_18824 n3_11864_18824 0.0
V27883 n1_11864_19007 n3_11864_19007 0.0
V27884 n1_11864_19040 n3_11864_19040 0.0
V27885 n1_11864_19223 n3_11864_19223 0.0
V27886 n1_11864_19256 n3_11864_19256 0.0
V27887 n1_11864_19404 n3_11864_19404 0.0
V27888 n1_11864_19439 n3_11864_19439 0.0
V27889 n1_11864_19472 n3_11864_19472 0.0
V27890 n1_11864_19655 n3_11864_19655 0.0
V27891 n1_11864_19688 n3_11864_19688 0.0
V27892 n1_11864_19871 n3_11864_19871 0.0
V27893 n1_11864_19904 n3_11864_19904 0.0
V27894 n1_11864_20087 n3_11864_20087 0.0
V27895 n1_11864_20120 n3_11864_20120 0.0
V27896 n1_11864_20303 n3_11864_20303 0.0
V27897 n1_11864_20336 n3_11864_20336 0.0
V27898 n1_11864_20519 n3_11864_20519 0.0
V27899 n1_11864_20552 n3_11864_20552 0.0
V27900 n1_11864_20687 n3_11864_20687 0.0
V27901 n1_11864_20735 n3_11864_20735 0.0
V27902 n1_11864_20768 n3_11864_20768 0.0
V27903 n1_11864_20951 n3_11864_20951 0.0
V27904 n1_11864_20984 n3_11864_20984 0.0
V27905 n1_13650_215 n3_13650_215 0.0
V27906 n1_13650_248 n3_13650_248 0.0
V27907 n1_13650_383 n3_13650_383 0.0
V27908 n1_13650_431 n3_13650_431 0.0
V27909 n1_13650_464 n3_13650_464 0.0
V27910 n1_13650_647 n3_13650_647 0.0
V27911 n1_13650_680 n3_13650_680 0.0
V27912 n1_13650_863 n3_13650_863 0.0
V27913 n1_13650_896 n3_13650_896 0.0
V27914 n1_13650_1079 n3_13650_1079 0.0
V27915 n1_13650_1112 n3_13650_1112 0.0
V27916 n1_13650_1295 n3_13650_1295 0.0
V27917 n1_13650_1328 n3_13650_1328 0.0
V27918 n1_13650_1511 n3_13650_1511 0.0
V27919 n1_13650_1544 n3_13650_1544 0.0
V27920 n1_13650_1727 n3_13650_1727 0.0
V27921 n1_13650_1760 n3_13650_1760 0.0
V27922 n1_13650_1894 n3_13650_1894 0.0
V27923 n1_13650_1943 n3_13650_1943 0.0
V27924 n1_13650_1976 n3_13650_1976 0.0
V27925 n1_13650_2159 n3_13650_2159 0.0
V27926 n1_13650_2192 n3_13650_2192 0.0
V27927 n1_13650_2375 n3_13650_2375 0.0
V27928 n1_13650_2408 n3_13650_2408 0.0
V27929 n1_13650_2445 n3_13650_2445 0.0
V27930 n1_13650_2542 n3_13650_2542 0.0
V27931 n1_13650_2543 n3_13650_2543 0.0
V27932 n1_13650_2591 n3_13650_2591 0.0
V27933 n1_13650_2624 n3_13650_2624 0.0
V27934 n1_13650_18527 n3_13650_18527 0.0
V27935 n1_13650_18575 n3_13650_18575 0.0
V27936 n1_13650_18608 n3_13650_18608 0.0
V27937 n1_13650_18764 n3_13650_18764 0.0
V27938 n1_13650_18791 n3_13650_18791 0.0
V27939 n1_13650_18824 n3_13650_18824 0.0
V27940 n1_13650_19007 n3_13650_19007 0.0
V27941 n1_13650_19040 n3_13650_19040 0.0
V27942 n1_13650_19223 n3_13650_19223 0.0
V27943 n1_13650_19256 n3_13650_19256 0.0
V27944 n1_13650_19412 n3_13650_19412 0.0
V27945 n1_13650_19439 n3_13650_19439 0.0
V27946 n1_13650_19472 n3_13650_19472 0.0
V27947 n1_13650_19655 n3_13650_19655 0.0
V27948 n1_13650_19688 n3_13650_19688 0.0
V27949 n1_13650_19871 n3_13650_19871 0.0
V27950 n1_13650_19904 n3_13650_19904 0.0
V27951 n1_13650_20087 n3_13650_20087 0.0
V27952 n1_13650_20120 n3_13650_20120 0.0
V27953 n1_13650_20303 n3_13650_20303 0.0
V27954 n1_13650_20336 n3_13650_20336 0.0
V27955 n1_13650_20519 n3_13650_20519 0.0
V27956 n1_13650_20552 n3_13650_20552 0.0
V27957 n1_13650_20687 n3_13650_20687 0.0
V27958 n1_13650_20735 n3_13650_20735 0.0
V27959 n1_13650_20768 n3_13650_20768 0.0
V27960 n1_13650_20951 n3_13650_20951 0.0
V27961 n1_13650_20984 n3_13650_20984 0.0
V27962 n1_13833_215 n3_13833_215 0.0
V27963 n1_13833_248 n3_13833_248 0.0
V27964 n1_13833_383 n3_13833_383 0.0
V27965 n1_13833_431 n3_13833_431 0.0
V27966 n1_13833_464 n3_13833_464 0.0
V27967 n1_13833_647 n3_13833_647 0.0
V27968 n1_13833_680 n3_13833_680 0.0
V27969 n1_13833_863 n3_13833_863 0.0
V27970 n1_13833_896 n3_13833_896 0.0
V27971 n1_13833_1079 n3_13833_1079 0.0
V27972 n1_13833_1112 n3_13833_1112 0.0
V27973 n1_13833_1295 n3_13833_1295 0.0
V27974 n1_13833_1328 n3_13833_1328 0.0
V27975 n1_13833_1727 n3_13833_1727 0.0
V27976 n1_13833_1760 n3_13833_1760 0.0
V27977 n1_13833_1894 n3_13833_1894 0.0
V27978 n1_13833_1943 n3_13833_1943 0.0
V27979 n1_13833_1976 n3_13833_1976 0.0
V27980 n1_13833_2159 n3_13833_2159 0.0
V27981 n1_13833_2192 n3_13833_2192 0.0
V27982 n1_13833_2375 n3_13833_2375 0.0
V27983 n1_13833_2408 n3_13833_2408 0.0
V27984 n1_13833_2445 n3_13833_2445 0.0
V27985 n1_13833_2542 n3_13833_2542 0.0
V27986 n1_13833_2543 n3_13833_2543 0.0
V27987 n1_13833_2591 n3_13833_2591 0.0
V27988 n1_13833_2624 n3_13833_2624 0.0
V27989 n1_13833_2807 n3_13833_2807 0.0
V27990 n1_13833_2840 n3_13833_2840 0.0
V27991 n1_13833_2877 n3_13833_2877 0.0
V27992 n1_13833_2974 n3_13833_2974 0.0
V27993 n1_13833_3023 n3_13833_3023 0.0
V27994 n1_13833_3056 n3_13833_3056 0.0
V27995 n1_13833_3239 n3_13833_3239 0.0
V27996 n1_13833_3272 n3_13833_3272 0.0
V27997 n1_13833_3455 n3_13833_3455 0.0
V27998 n1_13833_3488 n3_13833_3488 0.0
V27999 n1_13833_3622 n3_13833_3622 0.0
V28000 n1_13833_3671 n3_13833_3671 0.0
V28001 n1_13833_3704 n3_13833_3704 0.0
V28002 n1_13833_4054 n3_13833_4054 0.0
V28003 n1_13833_4103 n3_13833_4103 0.0
V28004 n1_13833_4136 n3_13833_4136 0.0
V28005 n1_13833_4270 n3_13833_4270 0.0
V28006 n1_13833_4319 n3_13833_4319 0.0
V28007 n1_13833_4352 n3_13833_4352 0.0
V28008 n1_13833_4535 n3_13833_4535 0.0
V28009 n1_13833_4568 n3_13833_4568 0.0
V28010 n1_13833_4702 n3_13833_4702 0.0
V28011 n1_13833_4751 n3_13833_4751 0.0
V28012 n1_13833_4784 n3_13833_4784 0.0
V28013 n1_13833_4967 n3_13833_4967 0.0
V28014 n1_13833_5000 n3_13833_5000 0.0
V28015 n1_13833_5134 n3_13833_5134 0.0
V28016 n1_13833_5183 n3_13833_5183 0.0
V28017 n1_13833_5216 n3_13833_5216 0.0
V28018 n1_13833_5350 n3_13833_5350 0.0
V28019 n1_13833_5399 n3_13833_5399 0.0
V28020 n1_13833_5432 n3_13833_5432 0.0
V28021 n1_13833_5615 n3_13833_5615 0.0
V28022 n1_13833_5648 n3_13833_5648 0.0
V28023 n1_13833_5782 n3_13833_5782 0.0
V28024 n1_13833_5831 n3_13833_5831 0.0
V28025 n1_13833_5864 n3_13833_5864 0.0
V28026 n1_13833_6263 n3_13833_6263 0.0
V28027 n1_13833_6296 n3_13833_6296 0.0
V28028 n1_13833_6430 n3_13833_6430 0.0
V28029 n1_13833_6479 n3_13833_6479 0.0
V28030 n1_13833_6512 n3_13833_6512 0.0
V28031 n1_13833_6646 n3_13833_6646 0.0
V28032 n1_13833_6695 n3_13833_6695 0.0
V28033 n1_13833_6728 n3_13833_6728 0.0
V28034 n1_13833_6911 n3_13833_6911 0.0
V28035 n1_13833_6944 n3_13833_6944 0.0
V28036 n1_13833_7127 n3_13833_7127 0.0
V28037 n1_13833_7160 n3_13833_7160 0.0
V28038 n1_13833_7343 n3_13833_7343 0.0
V28039 n1_13833_7376 n3_13833_7376 0.0
V28040 n1_13833_7559 n3_13833_7559 0.0
V28041 n1_13833_7592 n3_13833_7592 0.0
V28042 n1_13833_7775 n3_13833_7775 0.0
V28043 n1_13833_7808 n3_13833_7808 0.0
V28044 n1_13833_7845 n3_13833_7845 0.0
V28045 n1_13833_7942 n3_13833_7942 0.0
V28046 n1_13833_7991 n3_13833_7991 0.0
V28047 n1_13833_8024 n3_13833_8024 0.0
V28048 n1_13833_8207 n3_13833_8207 0.0
V28049 n1_13833_8240 n3_13833_8240 0.0
V28050 n1_13833_8456 n3_13833_8456 0.0
V28051 n1_13833_8639 n3_13833_8639 0.0
V28052 n1_13833_8672 n3_13833_8672 0.0
V28053 n1_13833_8806 n3_13833_8806 0.0
V28054 n1_13833_8855 n3_13833_8855 0.0
V28055 n1_13833_8888 n3_13833_8888 0.0
V28056 n1_13833_8925 n3_13833_8925 0.0
V28057 n1_13833_9022 n3_13833_9022 0.0
V28058 n1_13833_9071 n3_13833_9071 0.0
V28059 n1_13833_9104 n3_13833_9104 0.0
V28060 n1_13833_9287 n3_13833_9287 0.0
V28061 n1_13833_9320 n3_13833_9320 0.0
V28062 n1_13833_9503 n3_13833_9503 0.0
V28063 n1_13833_9536 n3_13833_9536 0.0
V28064 n1_13833_9719 n3_13833_9719 0.0
V28065 n1_13833_9752 n3_13833_9752 0.0
V28066 n1_13833_9886 n3_13833_9886 0.0
V28067 n1_13833_9935 n3_13833_9935 0.0
V28068 n1_13833_9968 n3_13833_9968 0.0
V28069 n1_13833_10005 n3_13833_10005 0.0
V28070 n1_13833_10102 n3_13833_10102 0.0
V28071 n1_13833_10151 n3_13833_10151 0.0
V28072 n1_13833_10184 n3_13833_10184 0.0
V28073 n1_13833_10367 n3_13833_10367 0.0
V28074 n1_13833_10400 n3_13833_10400 0.0
V28075 n1_13833_10799 n3_13833_10799 0.0
V28076 n1_13833_10832 n3_13833_10832 0.0
V28077 n1_13833_10988 n3_13833_10988 0.0
V28078 n1_13833_11015 n3_13833_11015 0.0
V28079 n1_13833_11048 n3_13833_11048 0.0
V28080 n1_13833_11204 n3_13833_11204 0.0
V28081 n1_13833_11231 n3_13833_11231 0.0
V28082 n1_13833_11264 n3_13833_11264 0.0
V28083 n1_13833_11447 n3_13833_11447 0.0
V28084 n1_13833_11480 n3_13833_11480 0.0
V28085 n1_13833_11663 n3_13833_11663 0.0
V28086 n1_13833_11696 n3_13833_11696 0.0
V28087 n1_13833_11879 n3_13833_11879 0.0
V28088 n1_13833_11912 n3_13833_11912 0.0
V28089 n1_13833_12068 n3_13833_12068 0.0
V28090 n1_13833_12095 n3_13833_12095 0.0
V28091 n1_13833_12128 n3_13833_12128 0.0
V28092 n1_13833_12284 n3_13833_12284 0.0
V28093 n1_13833_12311 n3_13833_12311 0.0
V28094 n1_13833_12344 n3_13833_12344 0.0
V28095 n1_13833_12527 n3_13833_12527 0.0
V28096 n1_13833_12560 n3_13833_12560 0.0
V28097 n1_13833_12743 n3_13833_12743 0.0
V28098 n1_13833_12959 n3_13833_12959 0.0
V28099 n1_13833_12992 n3_13833_12992 0.0
V28100 n1_13833_13175 n3_13833_13175 0.0
V28101 n1_13833_13208 n3_13833_13208 0.0
V28102 n1_13833_13391 n3_13833_13391 0.0
V28103 n1_13833_13424 n3_13833_13424 0.0
V28104 n1_13833_13607 n3_13833_13607 0.0
V28105 n1_13833_13640 n3_13833_13640 0.0
V28106 n1_13833_13823 n3_13833_13823 0.0
V28107 n1_13833_13856 n3_13833_13856 0.0
V28108 n1_13833_14039 n3_13833_14039 0.0
V28109 n1_13833_14072 n3_13833_14072 0.0
V28110 n1_13833_14220 n3_13833_14220 0.0
V28111 n1_13833_14255 n3_13833_14255 0.0
V28112 n1_13833_14288 n3_13833_14288 0.0
V28113 n1_13833_14471 n3_13833_14471 0.0
V28114 n1_13833_14504 n3_13833_14504 0.0
V28115 n1_13833_14652 n3_13833_14652 0.0
V28116 n1_13833_14687 n3_13833_14687 0.0
V28117 n1_13833_14720 n3_13833_14720 0.0
V28118 n1_13833_14868 n3_13833_14868 0.0
V28119 n1_13833_14903 n3_13833_14903 0.0
V28120 n1_13833_14936 n3_13833_14936 0.0
V28121 n1_13833_15335 n3_13833_15335 0.0
V28122 n1_13833_15368 n3_13833_15368 0.0
V28123 n1_13833_15524 n3_13833_15524 0.0
V28124 n1_13833_15551 n3_13833_15551 0.0
V28125 n1_13833_15584 n3_13833_15584 0.0
V28126 n1_13833_15767 n3_13833_15767 0.0
V28127 n1_13833_15800 n3_13833_15800 0.0
V28128 n1_13833_15956 n3_13833_15956 0.0
V28129 n1_13833_15983 n3_13833_15983 0.0
V28130 n1_13833_16016 n3_13833_16016 0.0
V28131 n1_13833_16199 n3_13833_16199 0.0
V28132 n1_13833_16232 n3_13833_16232 0.0
V28133 n1_13833_16415 n3_13833_16415 0.0
V28134 n1_13833_16448 n3_13833_16448 0.0
V28135 n1_13833_16604 n3_13833_16604 0.0
V28136 n1_13833_16631 n3_13833_16631 0.0
V28137 n1_13833_16664 n3_13833_16664 0.0
V28138 n1_13833_16847 n3_13833_16847 0.0
V28139 n1_13833_16880 n3_13833_16880 0.0
V28140 n1_13833_17063 n3_13833_17063 0.0
V28141 n1_13833_17096 n3_13833_17096 0.0
V28142 n1_13833_17495 n3_13833_17495 0.0
V28143 n1_13833_17528 n3_13833_17528 0.0
V28144 n1_13833_17684 n3_13833_17684 0.0
V28145 n1_13833_17711 n3_13833_17711 0.0
V28146 n1_13833_17744 n3_13833_17744 0.0
V28147 n1_13833_17927 n3_13833_17927 0.0
V28148 n1_13833_17960 n3_13833_17960 0.0
V28149 n1_13833_18094 n3_13833_18094 0.0
V28150 n1_13833_18143 n3_13833_18143 0.0
V28151 n1_13833_18176 n3_13833_18176 0.0
V28152 n1_13833_18324 n3_13833_18324 0.0
V28153 n1_13833_18332 n3_13833_18332 0.0
V28154 n1_13833_18359 n3_13833_18359 0.0
V28155 n1_13833_18392 n3_13833_18392 0.0
V28156 n1_13833_18527 n3_13833_18527 0.0
V28157 n1_13833_18575 n3_13833_18575 0.0
V28158 n1_13833_18608 n3_13833_18608 0.0
V28159 n1_13833_18764 n3_13833_18764 0.0
V28160 n1_13833_18791 n3_13833_18791 0.0
V28161 n1_13833_18824 n3_13833_18824 0.0
V28162 n1_13833_19007 n3_13833_19007 0.0
V28163 n1_13833_19040 n3_13833_19040 0.0
V28164 n1_13833_19223 n3_13833_19223 0.0
V28165 n1_13833_19256 n3_13833_19256 0.0
V28166 n1_13833_19404 n3_13833_19404 0.0
V28167 n1_13833_19412 n3_13833_19412 0.0
V28168 n1_13833_19439 n3_13833_19439 0.0
V28169 n1_13833_19472 n3_13833_19472 0.0
V28170 n1_13833_19871 n3_13833_19871 0.0
V28171 n1_13833_19904 n3_13833_19904 0.0
V28172 n1_13833_20087 n3_13833_20087 0.0
V28173 n1_13833_20120 n3_13833_20120 0.0
V28174 n1_13833_20303 n3_13833_20303 0.0
V28175 n1_13833_20336 n3_13833_20336 0.0
V28176 n1_13833_20519 n3_13833_20519 0.0
V28177 n1_13833_20552 n3_13833_20552 0.0
V28178 n1_13833_20687 n3_13833_20687 0.0
V28179 n1_13833_20735 n3_13833_20735 0.0
V28180 n1_13833_20768 n3_13833_20768 0.0
V28181 n1_13833_20951 n3_13833_20951 0.0
V28182 n1_13833_20984 n3_13833_20984 0.0
V28183 n1_13880_431 n3_13880_431 0.0
V28184 n1_13880_464 n3_13880_464 0.0
V28185 n1_13880_4967 n3_13880_4967 0.0
V28186 n1_13880_5000 n3_13880_5000 0.0
V28187 n1_13880_7160 n3_13880_7160 0.0
V28188 n1_13880_9503 n3_13880_9503 0.0
V28189 n1_13880_9536 n3_13880_9536 0.0
V28190 n1_13880_11663 n3_13880_11663 0.0
V28191 n1_13880_11696 n3_13880_11696 0.0
V28192 n1_13880_14039 n3_13880_14039 0.0
V28193 n1_13880_16199 n3_13880_16199 0.0
V28194 n1_13880_16232 n3_13880_16232 0.0
V28195 n1_13880_18392 n3_13880_18392 0.0
V28196 n1_13880_18527 n3_13880_18527 0.0
V28197 n1_13880_20687 n3_13880_20687 0.0
V28198 n1_13880_20735 n3_13880_20735 0.0
V28199 n1_13880_20768 n3_13880_20768 0.0
V28200 n1_14021_215 n3_14021_215 0.0
V28201 n1_14021_248 n3_14021_248 0.0
V28202 n1_14021_383 n3_14021_383 0.0
V28203 n1_14021_431 n3_14021_431 0.0
V28204 n1_14021_647 n3_14021_647 0.0
V28205 n1_14021_680 n3_14021_680 0.0
V28206 n1_14021_863 n3_14021_863 0.0
V28207 n1_14021_896 n3_14021_896 0.0
V28208 n1_14021_1079 n3_14021_1079 0.0
V28209 n1_14021_1112 n3_14021_1112 0.0
V28210 n1_14021_1295 n3_14021_1295 0.0
V28211 n1_14021_1328 n3_14021_1328 0.0
V28212 n1_14021_1511 n3_14021_1511 0.0
V28213 n1_14021_1544 n3_14021_1544 0.0
V28214 n1_14021_1727 n3_14021_1727 0.0
V28215 n1_14021_1760 n3_14021_1760 0.0
V28216 n1_14021_1894 n3_14021_1894 0.0
V28217 n1_14021_1943 n3_14021_1943 0.0
V28218 n1_14021_1976 n3_14021_1976 0.0
V28219 n1_14021_2159 n3_14021_2159 0.0
V28220 n1_14021_2192 n3_14021_2192 0.0
V28221 n1_14021_2375 n3_14021_2375 0.0
V28222 n1_14021_2408 n3_14021_2408 0.0
V28223 n1_14021_2445 n3_14021_2445 0.0
V28224 n1_14021_2542 n3_14021_2542 0.0
V28225 n1_14021_2543 n3_14021_2543 0.0
V28226 n1_14021_2591 n3_14021_2591 0.0
V28227 n1_14021_2624 n3_14021_2624 0.0
V28228 n1_14021_2807 n3_14021_2807 0.0
V28229 n1_14021_2840 n3_14021_2840 0.0
V28230 n1_14021_2877 n3_14021_2877 0.0
V28231 n1_14021_2974 n3_14021_2974 0.0
V28232 n1_14021_3023 n3_14021_3023 0.0
V28233 n1_14021_3056 n3_14021_3056 0.0
V28234 n1_14021_3239 n3_14021_3239 0.0
V28235 n1_14021_3272 n3_14021_3272 0.0
V28236 n1_14021_3455 n3_14021_3455 0.0
V28237 n1_14021_3488 n3_14021_3488 0.0
V28238 n1_14021_3622 n3_14021_3622 0.0
V28239 n1_14021_3671 n3_14021_3671 0.0
V28240 n1_14021_3704 n3_14021_3704 0.0
V28241 n1_14021_3887 n3_14021_3887 0.0
V28242 n1_14021_3920 n3_14021_3920 0.0
V28243 n1_14021_4054 n3_14021_4054 0.0
V28244 n1_14021_4103 n3_14021_4103 0.0
V28245 n1_14021_4136 n3_14021_4136 0.0
V28246 n1_14021_4270 n3_14021_4270 0.0
V28247 n1_14021_4319 n3_14021_4319 0.0
V28248 n1_14021_4352 n3_14021_4352 0.0
V28249 n1_14021_4535 n3_14021_4535 0.0
V28250 n1_14021_4568 n3_14021_4568 0.0
V28251 n1_14021_4702 n3_14021_4702 0.0
V28252 n1_14021_4751 n3_14021_4751 0.0
V28253 n1_14021_4784 n3_14021_4784 0.0
V28254 n1_14021_5000 n3_14021_5000 0.0
V28255 n1_14021_5134 n3_14021_5134 0.0
V28256 n1_14021_5183 n3_14021_5183 0.0
V28257 n1_14021_5216 n3_14021_5216 0.0
V28258 n1_14021_5350 n3_14021_5350 0.0
V28259 n1_14021_5399 n3_14021_5399 0.0
V28260 n1_14021_5432 n3_14021_5432 0.0
V28261 n1_14021_5615 n3_14021_5615 0.0
V28262 n1_14021_5648 n3_14021_5648 0.0
V28263 n1_14021_5782 n3_14021_5782 0.0
V28264 n1_14021_5831 n3_14021_5831 0.0
V28265 n1_14021_5864 n3_14021_5864 0.0
V28266 n1_14021_6047 n3_14021_6047 0.0
V28267 n1_14021_6080 n3_14021_6080 0.0
V28268 n1_14021_6263 n3_14021_6263 0.0
V28269 n1_14021_6296 n3_14021_6296 0.0
V28270 n1_14021_6430 n3_14021_6430 0.0
V28271 n1_14021_6479 n3_14021_6479 0.0
V28272 n1_14021_6512 n3_14021_6512 0.0
V28273 n1_14021_6646 n3_14021_6646 0.0
V28274 n1_14021_6695 n3_14021_6695 0.0
V28275 n1_14021_6728 n3_14021_6728 0.0
V28276 n1_14021_6911 n3_14021_6911 0.0
V28277 n1_14021_6944 n3_14021_6944 0.0
V28278 n1_14021_7127 n3_14021_7127 0.0
V28279 n1_14021_7160 n3_14021_7160 0.0
V28280 n1_14021_7343 n3_14021_7343 0.0
V28281 n1_14021_7376 n3_14021_7376 0.0
V28282 n1_14021_7559 n3_14021_7559 0.0
V28283 n1_14021_7592 n3_14021_7592 0.0
V28284 n1_14021_7775 n3_14021_7775 0.0
V28285 n1_14021_7808 n3_14021_7808 0.0
V28286 n1_14021_7845 n3_14021_7845 0.0
V28287 n1_14021_7942 n3_14021_7942 0.0
V28288 n1_14021_7991 n3_14021_7991 0.0
V28289 n1_14021_8024 n3_14021_8024 0.0
V28290 n1_14021_8207 n3_14021_8207 0.0
V28291 n1_14021_8240 n3_14021_8240 0.0
V28292 n1_14021_8423 n3_14021_8423 0.0
V28293 n1_14021_8456 n3_14021_8456 0.0
V28294 n1_14021_8639 n3_14021_8639 0.0
V28295 n1_14021_8672 n3_14021_8672 0.0
V28296 n1_14021_8806 n3_14021_8806 0.0
V28297 n1_14021_8855 n3_14021_8855 0.0
V28298 n1_14021_8888 n3_14021_8888 0.0
V28299 n1_14021_8925 n3_14021_8925 0.0
V28300 n1_14021_9022 n3_14021_9022 0.0
V28301 n1_14021_9071 n3_14021_9071 0.0
V28302 n1_14021_9104 n3_14021_9104 0.0
V28303 n1_14021_9287 n3_14021_9287 0.0
V28304 n1_14021_9320 n3_14021_9320 0.0
V28305 n1_14021_9503 n3_14021_9503 0.0
V28306 n1_14021_9536 n3_14021_9536 0.0
V28307 n1_14021_9719 n3_14021_9719 0.0
V28308 n1_14021_9752 n3_14021_9752 0.0
V28309 n1_14021_9886 n3_14021_9886 0.0
V28310 n1_14021_9935 n3_14021_9935 0.0
V28311 n1_14021_9968 n3_14021_9968 0.0
V28312 n1_14021_10005 n3_14021_10005 0.0
V28313 n1_14021_10102 n3_14021_10102 0.0
V28314 n1_14021_10151 n3_14021_10151 0.0
V28315 n1_14021_10184 n3_14021_10184 0.0
V28316 n1_14021_10367 n3_14021_10367 0.0
V28317 n1_14021_10400 n3_14021_10400 0.0
V28318 n1_14021_10616 n3_14021_10616 0.0
V28319 n1_14021_10799 n3_14021_10799 0.0
V28320 n1_14021_10832 n3_14021_10832 0.0
V28321 n1_14021_10988 n3_14021_10988 0.0
V28322 n1_14021_11015 n3_14021_11015 0.0
V28323 n1_14021_11048 n3_14021_11048 0.0
V28324 n1_14021_11204 n3_14021_11204 0.0
V28325 n1_14021_11231 n3_14021_11231 0.0
V28326 n1_14021_11264 n3_14021_11264 0.0
V28327 n1_14021_11447 n3_14021_11447 0.0
V28328 n1_14021_11480 n3_14021_11480 0.0
V28329 n1_14021_11663 n3_14021_11663 0.0
V28330 n1_14021_11696 n3_14021_11696 0.0
V28331 n1_14021_11879 n3_14021_11879 0.0
V28332 n1_14021_11912 n3_14021_11912 0.0
V28333 n1_14021_12068 n3_14021_12068 0.0
V28334 n1_14021_12095 n3_14021_12095 0.0
V28335 n1_14021_12128 n3_14021_12128 0.0
V28336 n1_14021_12284 n3_14021_12284 0.0
V28337 n1_14021_12311 n3_14021_12311 0.0
V28338 n1_14021_12344 n3_14021_12344 0.0
V28339 n1_14021_12527 n3_14021_12527 0.0
V28340 n1_14021_12560 n3_14021_12560 0.0
V28341 n1_14021_12743 n3_14021_12743 0.0
V28342 n1_14021_12776 n3_14021_12776 0.0
V28343 n1_14021_12959 n3_14021_12959 0.0
V28344 n1_14021_12992 n3_14021_12992 0.0
V28345 n1_14021_13175 n3_14021_13175 0.0
V28346 n1_14021_13208 n3_14021_13208 0.0
V28347 n1_14021_13391 n3_14021_13391 0.0
V28348 n1_14021_13424 n3_14021_13424 0.0
V28349 n1_14021_13607 n3_14021_13607 0.0
V28350 n1_14021_13640 n3_14021_13640 0.0
V28351 n1_14021_13823 n3_14021_13823 0.0
V28352 n1_14021_13856 n3_14021_13856 0.0
V28353 n1_14021_14039 n3_14021_14039 0.0
V28354 n1_14021_14072 n3_14021_14072 0.0
V28355 n1_14021_14220 n3_14021_14220 0.0
V28356 n1_14021_14255 n3_14021_14255 0.0
V28357 n1_14021_14288 n3_14021_14288 0.0
V28358 n1_14021_14471 n3_14021_14471 0.0
V28359 n1_14021_14504 n3_14021_14504 0.0
V28360 n1_14021_14652 n3_14021_14652 0.0
V28361 n1_14021_14687 n3_14021_14687 0.0
V28362 n1_14021_14720 n3_14021_14720 0.0
V28363 n1_14021_14868 n3_14021_14868 0.0
V28364 n1_14021_14903 n3_14021_14903 0.0
V28365 n1_14021_14936 n3_14021_14936 0.0
V28366 n1_14021_15119 n3_14021_15119 0.0
V28367 n1_14021_15152 n3_14021_15152 0.0
V28368 n1_14021_15335 n3_14021_15335 0.0
V28369 n1_14021_15368 n3_14021_15368 0.0
V28370 n1_14021_15524 n3_14021_15524 0.0
V28371 n1_14021_15551 n3_14021_15551 0.0
V28372 n1_14021_15584 n3_14021_15584 0.0
V28373 n1_14021_15767 n3_14021_15767 0.0
V28374 n1_14021_15800 n3_14021_15800 0.0
V28375 n1_14021_15956 n3_14021_15956 0.0
V28376 n1_14021_15983 n3_14021_15983 0.0
V28377 n1_14021_16016 n3_14021_16016 0.0
V28378 n1_14021_16199 n3_14021_16199 0.0
V28379 n1_14021_16415 n3_14021_16415 0.0
V28380 n1_14021_16448 n3_14021_16448 0.0
V28381 n1_14021_16604 n3_14021_16604 0.0
V28382 n1_14021_16631 n3_14021_16631 0.0
V28383 n1_14021_16664 n3_14021_16664 0.0
V28384 n1_14021_16847 n3_14021_16847 0.0
V28385 n1_14021_16880 n3_14021_16880 0.0
V28386 n1_14021_17063 n3_14021_17063 0.0
V28387 n1_14021_17096 n3_14021_17096 0.0
V28388 n1_14021_17252 n3_14021_17252 0.0
V28389 n1_14021_17279 n3_14021_17279 0.0
V28390 n1_14021_17312 n3_14021_17312 0.0
V28391 n1_14021_17495 n3_14021_17495 0.0
V28392 n1_14021_17528 n3_14021_17528 0.0
V28393 n1_14021_17684 n3_14021_17684 0.0
V28394 n1_14021_17711 n3_14021_17711 0.0
V28395 n1_14021_17744 n3_14021_17744 0.0
V28396 n1_14021_17927 n3_14021_17927 0.0
V28397 n1_14021_17960 n3_14021_17960 0.0
V28398 n1_14021_18094 n3_14021_18094 0.0
V28399 n1_14021_18143 n3_14021_18143 0.0
V28400 n1_14021_18176 n3_14021_18176 0.0
V28401 n1_14021_18324 n3_14021_18324 0.0
V28402 n1_14021_18332 n3_14021_18332 0.0
V28403 n1_14021_18359 n3_14021_18359 0.0
V28404 n1_14021_18392 n3_14021_18392 0.0
V28405 n1_14021_18527 n3_14021_18527 0.0
V28406 n1_14021_18575 n3_14021_18575 0.0
V28407 n1_14021_18608 n3_14021_18608 0.0
V28408 n1_14021_18764 n3_14021_18764 0.0
V28409 n1_14021_18791 n3_14021_18791 0.0
V28410 n1_14021_18824 n3_14021_18824 0.0
V28411 n1_14021_19007 n3_14021_19007 0.0
V28412 n1_14021_19040 n3_14021_19040 0.0
V28413 n1_14021_19223 n3_14021_19223 0.0
V28414 n1_14021_19256 n3_14021_19256 0.0
V28415 n1_14021_19404 n3_14021_19404 0.0
V28416 n1_14021_19412 n3_14021_19412 0.0
V28417 n1_14021_19439 n3_14021_19439 0.0
V28418 n1_14021_19472 n3_14021_19472 0.0
V28419 n1_14021_19655 n3_14021_19655 0.0
V28420 n1_14021_19688 n3_14021_19688 0.0
V28421 n1_14021_19871 n3_14021_19871 0.0
V28422 n1_14021_19904 n3_14021_19904 0.0
V28423 n1_14021_20087 n3_14021_20087 0.0
V28424 n1_14021_20120 n3_14021_20120 0.0
V28425 n1_14021_20303 n3_14021_20303 0.0
V28426 n1_14021_20336 n3_14021_20336 0.0
V28427 n1_14021_20519 n3_14021_20519 0.0
V28428 n1_14021_20552 n3_14021_20552 0.0
V28429 n1_14021_20687 n3_14021_20687 0.0
V28430 n1_14021_20768 n3_14021_20768 0.0
V28431 n1_14021_20951 n3_14021_20951 0.0
V28432 n1_14021_20984 n3_14021_20984 0.0
V28433 n1_14114_215 n3_14114_215 0.0
V28434 n1_14114_248 n3_14114_248 0.0
V28435 n1_14114_383 n3_14114_383 0.0
V28436 n1_14114_431 n3_14114_431 0.0
V28437 n1_14114_464 n3_14114_464 0.0
V28438 n1_14114_647 n3_14114_647 0.0
V28439 n1_14114_680 n3_14114_680 0.0
V28440 n1_14114_863 n3_14114_863 0.0
V28441 n1_14114_896 n3_14114_896 0.0
V28442 n1_14114_1079 n3_14114_1079 0.0
V28443 n1_14114_1112 n3_14114_1112 0.0
V28444 n1_14114_1295 n3_14114_1295 0.0
V28445 n1_14114_1328 n3_14114_1328 0.0
V28446 n1_14114_1511 n3_14114_1511 0.0
V28447 n1_14114_1544 n3_14114_1544 0.0
V28448 n1_14114_1727 n3_14114_1727 0.0
V28449 n1_14114_1760 n3_14114_1760 0.0
V28450 n1_14114_1894 n3_14114_1894 0.0
V28451 n1_14114_1943 n3_14114_1943 0.0
V28452 n1_14114_1976 n3_14114_1976 0.0
V28453 n1_14114_2159 n3_14114_2159 0.0
V28454 n1_14114_2192 n3_14114_2192 0.0
V28455 n1_14114_2375 n3_14114_2375 0.0
V28456 n1_14114_2408 n3_14114_2408 0.0
V28457 n1_14114_2445 n3_14114_2445 0.0
V28458 n1_14114_2542 n3_14114_2542 0.0
V28459 n1_14114_2543 n3_14114_2543 0.0
V28460 n1_14114_2591 n3_14114_2591 0.0
V28461 n1_14114_2624 n3_14114_2624 0.0
V28462 n1_14114_18527 n3_14114_18527 0.0
V28463 n1_14114_18575 n3_14114_18575 0.0
V28464 n1_14114_18608 n3_14114_18608 0.0
V28465 n1_14114_18764 n3_14114_18764 0.0
V28466 n1_14114_18791 n3_14114_18791 0.0
V28467 n1_14114_18824 n3_14114_18824 0.0
V28468 n1_14114_19007 n3_14114_19007 0.0
V28469 n1_14114_19040 n3_14114_19040 0.0
V28470 n1_14114_19223 n3_14114_19223 0.0
V28471 n1_14114_19256 n3_14114_19256 0.0
V28472 n1_14114_19404 n3_14114_19404 0.0
V28473 n1_14114_19439 n3_14114_19439 0.0
V28474 n1_14114_19472 n3_14114_19472 0.0
V28475 n1_14114_19655 n3_14114_19655 0.0
V28476 n1_14114_19688 n3_14114_19688 0.0
V28477 n1_14114_19871 n3_14114_19871 0.0
V28478 n1_14114_19904 n3_14114_19904 0.0
V28479 n1_14114_20087 n3_14114_20087 0.0
V28480 n1_14114_20120 n3_14114_20120 0.0
V28481 n1_14114_20303 n3_14114_20303 0.0
V28482 n1_14114_20336 n3_14114_20336 0.0
V28483 n1_14114_20519 n3_14114_20519 0.0
V28484 n1_14114_20552 n3_14114_20552 0.0
V28485 n1_14114_20687 n3_14114_20687 0.0
V28486 n1_14114_20735 n3_14114_20735 0.0
V28487 n1_14114_20768 n3_14114_20768 0.0
V28488 n1_14114_20951 n3_14114_20951 0.0
V28489 n1_14114_20984 n3_14114_20984 0.0
V28490 n1_15900_215 n3_15900_215 0.0
V28491 n1_15900_248 n3_15900_248 0.0
V28492 n1_15900_383 n3_15900_383 0.0
V28493 n1_15900_431 n3_15900_431 0.0
V28494 n1_15900_464 n3_15900_464 0.0
V28495 n1_15900_647 n3_15900_647 0.0
V28496 n1_15900_680 n3_15900_680 0.0
V28497 n1_15900_863 n3_15900_863 0.0
V28498 n1_15900_896 n3_15900_896 0.0
V28499 n1_15900_1079 n3_15900_1079 0.0
V28500 n1_15900_1112 n3_15900_1112 0.0
V28501 n1_15900_1295 n3_15900_1295 0.0
V28502 n1_15900_1328 n3_15900_1328 0.0
V28503 n1_15900_1511 n3_15900_1511 0.0
V28504 n1_15900_1544 n3_15900_1544 0.0
V28505 n1_15900_1727 n3_15900_1727 0.0
V28506 n1_15900_1760 n3_15900_1760 0.0
V28507 n1_15900_1894 n3_15900_1894 0.0
V28508 n1_15900_1943 n3_15900_1943 0.0
V28509 n1_15900_1976 n3_15900_1976 0.0
V28510 n1_15900_2159 n3_15900_2159 0.0
V28511 n1_15900_2192 n3_15900_2192 0.0
V28512 n1_15900_2375 n3_15900_2375 0.0
V28513 n1_15900_2408 n3_15900_2408 0.0
V28514 n1_15900_2445 n3_15900_2445 0.0
V28515 n1_15900_2542 n3_15900_2542 0.0
V28516 n1_15900_2543 n3_15900_2543 0.0
V28517 n1_15900_2591 n3_15900_2591 0.0
V28518 n1_15900_2624 n3_15900_2624 0.0
V28519 n1_15900_18527 n3_15900_18527 0.0
V28520 n1_15900_18575 n3_15900_18575 0.0
V28521 n1_15900_18608 n3_15900_18608 0.0
V28522 n1_15900_18764 n3_15900_18764 0.0
V28523 n1_15900_18791 n3_15900_18791 0.0
V28524 n1_15900_18824 n3_15900_18824 0.0
V28525 n1_15900_19007 n3_15900_19007 0.0
V28526 n1_15900_19040 n3_15900_19040 0.0
V28527 n1_15900_19223 n3_15900_19223 0.0
V28528 n1_15900_19256 n3_15900_19256 0.0
V28529 n1_15900_19412 n3_15900_19412 0.0
V28530 n1_15900_19439 n3_15900_19439 0.0
V28531 n1_15900_19472 n3_15900_19472 0.0
V28532 n1_15900_19655 n3_15900_19655 0.0
V28533 n1_15900_19688 n3_15900_19688 0.0
V28534 n1_15900_19871 n3_15900_19871 0.0
V28535 n1_15900_19904 n3_15900_19904 0.0
V28536 n1_15900_20087 n3_15900_20087 0.0
V28537 n1_15900_20120 n3_15900_20120 0.0
V28538 n1_15900_20303 n3_15900_20303 0.0
V28539 n1_15900_20336 n3_15900_20336 0.0
V28540 n1_15900_20519 n3_15900_20519 0.0
V28541 n1_15900_20552 n3_15900_20552 0.0
V28542 n1_15900_20687 n3_15900_20687 0.0
V28543 n1_15900_20735 n3_15900_20735 0.0
V28544 n1_15900_20768 n3_15900_20768 0.0
V28545 n1_15900_20951 n3_15900_20951 0.0
V28546 n1_15900_20984 n3_15900_20984 0.0
V28547 n1_16083_215 n3_16083_215 0.0
V28548 n1_16083_248 n3_16083_248 0.0
V28549 n1_16083_383 n3_16083_383 0.0
V28550 n1_16083_431 n3_16083_431 0.0
V28551 n1_16083_464 n3_16083_464 0.0
V28552 n1_16083_647 n3_16083_647 0.0
V28553 n1_16083_680 n3_16083_680 0.0
V28554 n1_16083_863 n3_16083_863 0.0
V28555 n1_16083_896 n3_16083_896 0.0
V28556 n1_16083_1079 n3_16083_1079 0.0
V28557 n1_16083_1112 n3_16083_1112 0.0
V28558 n1_16083_1295 n3_16083_1295 0.0
V28559 n1_16083_1328 n3_16083_1328 0.0
V28560 n1_16083_1727 n3_16083_1727 0.0
V28561 n1_16083_1760 n3_16083_1760 0.0
V28562 n1_16083_1894 n3_16083_1894 0.0
V28563 n1_16083_1943 n3_16083_1943 0.0
V28564 n1_16083_1976 n3_16083_1976 0.0
V28565 n1_16083_2159 n3_16083_2159 0.0
V28566 n1_16083_2192 n3_16083_2192 0.0
V28567 n1_16083_2375 n3_16083_2375 0.0
V28568 n1_16083_2408 n3_16083_2408 0.0
V28569 n1_16083_2445 n3_16083_2445 0.0
V28570 n1_16083_2542 n3_16083_2542 0.0
V28571 n1_16083_2543 n3_16083_2543 0.0
V28572 n1_16083_2591 n3_16083_2591 0.0
V28573 n1_16083_2624 n3_16083_2624 0.0
V28574 n1_16083_2807 n3_16083_2807 0.0
V28575 n1_16083_2840 n3_16083_2840 0.0
V28576 n1_16083_2877 n3_16083_2877 0.0
V28577 n1_16083_2974 n3_16083_2974 0.0
V28578 n1_16083_3023 n3_16083_3023 0.0
V28579 n1_16083_3056 n3_16083_3056 0.0
V28580 n1_16083_3239 n3_16083_3239 0.0
V28581 n1_16083_3272 n3_16083_3272 0.0
V28582 n1_16083_3406 n3_16083_3406 0.0
V28583 n1_16083_3455 n3_16083_3455 0.0
V28584 n1_16083_3488 n3_16083_3488 0.0
V28585 n1_16083_3671 n3_16083_3671 0.0
V28586 n1_16083_3704 n3_16083_3704 0.0
V28587 n1_16083_4103 n3_16083_4103 0.0
V28588 n1_16083_4136 n3_16083_4136 0.0
V28589 n1_16083_4319 n3_16083_4319 0.0
V28590 n1_16083_4352 n3_16083_4352 0.0
V28591 n1_16083_4486 n3_16083_4486 0.0
V28592 n1_16083_4535 n3_16083_4535 0.0
V28593 n1_16083_4568 n3_16083_4568 0.0
V28594 n1_16083_4702 n3_16083_4702 0.0
V28595 n1_16083_4751 n3_16083_4751 0.0
V28596 n1_16083_4784 n3_16083_4784 0.0
V28597 n1_16083_4919 n3_16083_4919 0.0
V28598 n1_16083_4967 n3_16083_4967 0.0
V28599 n1_16083_5000 n3_16083_5000 0.0
V28600 n1_16083_5134 n3_16083_5134 0.0
V28601 n1_16083_5183 n3_16083_5183 0.0
V28602 n1_16083_5216 n3_16083_5216 0.0
V28603 n1_16083_5253 n3_16083_5253 0.0
V28604 n1_16083_5350 n3_16083_5350 0.0
V28605 n1_16083_5399 n3_16083_5399 0.0
V28606 n1_16083_5432 n3_16083_5432 0.0
V28607 n1_16083_5566 n3_16083_5566 0.0
V28608 n1_16083_5615 n3_16083_5615 0.0
V28609 n1_16083_5648 n3_16083_5648 0.0
V28610 n1_16083_5831 n3_16083_5831 0.0
V28611 n1_16083_5864 n3_16083_5864 0.0
V28612 n1_16083_6263 n3_16083_6263 0.0
V28613 n1_16083_6296 n3_16083_6296 0.0
V28614 n1_16083_6333 n3_16083_6333 0.0
V28615 n1_16083_6430 n3_16083_6430 0.0
V28616 n1_16083_6479 n3_16083_6479 0.0
V28617 n1_16083_6512 n3_16083_6512 0.0
V28618 n1_16083_6695 n3_16083_6695 0.0
V28619 n1_16083_6728 n3_16083_6728 0.0
V28620 n1_16083_6911 n3_16083_6911 0.0
V28621 n1_16083_6944 n3_16083_6944 0.0
V28622 n1_16083_7127 n3_16083_7127 0.0
V28623 n1_16083_7160 n3_16083_7160 0.0
V28624 n1_16083_7343 n3_16083_7343 0.0
V28625 n1_16083_7376 n3_16083_7376 0.0
V28626 n1_16083_7559 n3_16083_7559 0.0
V28627 n1_16083_7592 n3_16083_7592 0.0
V28628 n1_16083_7775 n3_16083_7775 0.0
V28629 n1_16083_7808 n3_16083_7808 0.0
V28630 n1_16083_7845 n3_16083_7845 0.0
V28631 n1_16083_7942 n3_16083_7942 0.0
V28632 n1_16083_7991 n3_16083_7991 0.0
V28633 n1_16083_8024 n3_16083_8024 0.0
V28634 n1_16083_8207 n3_16083_8207 0.0
V28635 n1_16083_8240 n3_16083_8240 0.0
V28636 n1_16083_8456 n3_16083_8456 0.0
V28637 n1_16083_8639 n3_16083_8639 0.0
V28638 n1_16083_8672 n3_16083_8672 0.0
V28639 n1_16083_8855 n3_16083_8855 0.0
V28640 n1_16083_8888 n3_16083_8888 0.0
V28641 n1_16083_8925 n3_16083_8925 0.0
V28642 n1_16083_9022 n3_16083_9022 0.0
V28643 n1_16083_9071 n3_16083_9071 0.0
V28644 n1_16083_9104 n3_16083_9104 0.0
V28645 n1_16083_9287 n3_16083_9287 0.0
V28646 n1_16083_9320 n3_16083_9320 0.0
V28647 n1_16083_9503 n3_16083_9503 0.0
V28648 n1_16083_9536 n3_16083_9536 0.0
V28649 n1_16083_9719 n3_16083_9719 0.0
V28650 n1_16083_9752 n3_16083_9752 0.0
V28651 n1_16083_9935 n3_16083_9935 0.0
V28652 n1_16083_9968 n3_16083_9968 0.0
V28653 n1_16083_10005 n3_16083_10005 0.0
V28654 n1_16083_10102 n3_16083_10102 0.0
V28655 n1_16083_10151 n3_16083_10151 0.0
V28656 n1_16083_10184 n3_16083_10184 0.0
V28657 n1_16083_10367 n3_16083_10367 0.0
V28658 n1_16083_10400 n3_16083_10400 0.0
V28659 n1_16083_10799 n3_16083_10799 0.0
V28660 n1_16083_10832 n3_16083_10832 0.0
V28661 n1_16083_11015 n3_16083_11015 0.0
V28662 n1_16083_11048 n3_16083_11048 0.0
V28663 n1_16083_11196 n3_16083_11196 0.0
V28664 n1_16083_11204 n3_16083_11204 0.0
V28665 n1_16083_11231 n3_16083_11231 0.0
V28666 n1_16083_11264 n3_16083_11264 0.0
V28667 n1_16083_11447 n3_16083_11447 0.0
V28668 n1_16083_11480 n3_16083_11480 0.0
V28669 n1_16083_11663 n3_16083_11663 0.0
V28670 n1_16083_11696 n3_16083_11696 0.0
V28671 n1_16083_11879 n3_16083_11879 0.0
V28672 n1_16083_11912 n3_16083_11912 0.0
V28673 n1_16083_12095 n3_16083_12095 0.0
V28674 n1_16083_12128 n3_16083_12128 0.0
V28675 n1_16083_12276 n3_16083_12276 0.0
V28676 n1_16083_12284 n3_16083_12284 0.0
V28677 n1_16083_12311 n3_16083_12311 0.0
V28678 n1_16083_12344 n3_16083_12344 0.0
V28679 n1_16083_12527 n3_16083_12527 0.0
V28680 n1_16083_12560 n3_16083_12560 0.0
V28681 n1_16083_12743 n3_16083_12743 0.0
V28682 n1_16083_12959 n3_16083_12959 0.0
V28683 n1_16083_12992 n3_16083_12992 0.0
V28684 n1_16083_13175 n3_16083_13175 0.0
V28685 n1_16083_13208 n3_16083_13208 0.0
V28686 n1_16083_13391 n3_16083_13391 0.0
V28687 n1_16083_13424 n3_16083_13424 0.0
V28688 n1_16083_13607 n3_16083_13607 0.0
V28689 n1_16083_13640 n3_16083_13640 0.0
V28690 n1_16083_13788 n3_16083_13788 0.0
V28691 n1_16083_13823 n3_16083_13823 0.0
V28692 n1_16083_13856 n3_16083_13856 0.0
V28693 n1_16083_14039 n3_16083_14039 0.0
V28694 n1_16083_14072 n3_16083_14072 0.0
V28695 n1_16083_14255 n3_16083_14255 0.0
V28696 n1_16083_14288 n3_16083_14288 0.0
V28697 n1_16083_14471 n3_16083_14471 0.0
V28698 n1_16083_14504 n3_16083_14504 0.0
V28699 n1_16083_14652 n3_16083_14652 0.0
V28700 n1_16083_14687 n3_16083_14687 0.0
V28701 n1_16083_14720 n3_16083_14720 0.0
V28702 n1_16083_14903 n3_16083_14903 0.0
V28703 n1_16083_14936 n3_16083_14936 0.0
V28704 n1_16083_15300 n3_16083_15300 0.0
V28705 n1_16083_15335 n3_16083_15335 0.0
V28706 n1_16083_15368 n3_16083_15368 0.0
V28707 n1_16083_15551 n3_16083_15551 0.0
V28708 n1_16083_15584 n3_16083_15584 0.0
V28709 n1_16083_15740 n3_16083_15740 0.0
V28710 n1_16083_15767 n3_16083_15767 0.0
V28711 n1_16083_15800 n3_16083_15800 0.0
V28712 n1_16083_15983 n3_16083_15983 0.0
V28713 n1_16083_16016 n3_16083_16016 0.0
V28714 n1_16083_16199 n3_16083_16199 0.0
V28715 n1_16083_16232 n3_16083_16232 0.0
V28716 n1_16083_16415 n3_16083_16415 0.0
V28717 n1_16083_16448 n3_16083_16448 0.0
V28718 n1_16083_16604 n3_16083_16604 0.0
V28719 n1_16083_16631 n3_16083_16631 0.0
V28720 n1_16083_16664 n3_16083_16664 0.0
V28721 n1_16083_16798 n3_16083_16798 0.0
V28722 n1_16083_16820 n3_16083_16820 0.0
V28723 n1_16083_16847 n3_16083_16847 0.0
V28724 n1_16083_16880 n3_16083_16880 0.0
V28725 n1_16083_17063 n3_16083_17063 0.0
V28726 n1_16083_17096 n3_16083_17096 0.0
V28727 n1_16083_17495 n3_16083_17495 0.0
V28728 n1_16083_17528 n3_16083_17528 0.0
V28729 n1_16083_17676 n3_16083_17676 0.0
V28730 n1_16083_17684 n3_16083_17684 0.0
V28731 n1_16083_17711 n3_16083_17711 0.0
V28732 n1_16083_17744 n3_16083_17744 0.0
V28733 n1_16083_17927 n3_16083_17927 0.0
V28734 n1_16083_17960 n3_16083_17960 0.0
V28735 n1_16083_18143 n3_16083_18143 0.0
V28736 n1_16083_18176 n3_16083_18176 0.0
V28737 n1_16083_18332 n3_16083_18332 0.0
V28738 n1_16083_18359 n3_16083_18359 0.0
V28739 n1_16083_18392 n3_16083_18392 0.0
V28740 n1_16083_18527 n3_16083_18527 0.0
V28741 n1_16083_18575 n3_16083_18575 0.0
V28742 n1_16083_18608 n3_16083_18608 0.0
V28743 n1_16083_18764 n3_16083_18764 0.0
V28744 n1_16083_18791 n3_16083_18791 0.0
V28745 n1_16083_18824 n3_16083_18824 0.0
V28746 n1_16083_19007 n3_16083_19007 0.0
V28747 n1_16083_19040 n3_16083_19040 0.0
V28748 n1_16083_19196 n3_16083_19196 0.0
V28749 n1_16083_19223 n3_16083_19223 0.0
V28750 n1_16083_19256 n3_16083_19256 0.0
V28751 n1_16083_19412 n3_16083_19412 0.0
V28752 n1_16083_19439 n3_16083_19439 0.0
V28753 n1_16083_19472 n3_16083_19472 0.0
V28754 n1_16083_19871 n3_16083_19871 0.0
V28755 n1_16083_19904 n3_16083_19904 0.0
V28756 n1_16083_20087 n3_16083_20087 0.0
V28757 n1_16083_20120 n3_16083_20120 0.0
V28758 n1_16083_20303 n3_16083_20303 0.0
V28759 n1_16083_20336 n3_16083_20336 0.0
V28760 n1_16083_20519 n3_16083_20519 0.0
V28761 n1_16083_20552 n3_16083_20552 0.0
V28762 n1_16083_20687 n3_16083_20687 0.0
V28763 n1_16083_20735 n3_16083_20735 0.0
V28764 n1_16083_20768 n3_16083_20768 0.0
V28765 n1_16083_20951 n3_16083_20951 0.0
V28766 n1_16083_20984 n3_16083_20984 0.0
V28767 n1_16130_431 n3_16130_431 0.0
V28768 n1_16130_464 n3_16130_464 0.0
V28769 n1_16130_4919 n3_16130_4919 0.0
V28770 n1_16130_4967 n3_16130_4967 0.0
V28771 n1_16130_5000 n3_16130_5000 0.0
V28772 n1_16130_7160 n3_16130_7160 0.0
V28773 n1_16130_9503 n3_16130_9503 0.0
V28774 n1_16130_9536 n3_16130_9536 0.0
V28775 n1_16130_11663 n3_16130_11663 0.0
V28776 n1_16130_11696 n3_16130_11696 0.0
V28777 n1_16130_14039 n3_16130_14039 0.0
V28778 n1_16130_16199 n3_16130_16199 0.0
V28779 n1_16130_16232 n3_16130_16232 0.0
V28780 n1_16130_18392 n3_16130_18392 0.0
V28781 n1_16130_18527 n3_16130_18527 0.0
V28782 n1_16130_20687 n3_16130_20687 0.0
V28783 n1_16130_20735 n3_16130_20735 0.0
V28784 n1_16130_20768 n3_16130_20768 0.0
V28785 n1_16271_215 n3_16271_215 0.0
V28786 n1_16271_248 n3_16271_248 0.0
V28787 n1_16271_383 n3_16271_383 0.0
V28788 n1_16271_431 n3_16271_431 0.0
V28789 n1_16271_647 n3_16271_647 0.0
V28790 n1_16271_680 n3_16271_680 0.0
V28791 n1_16271_863 n3_16271_863 0.0
V28792 n1_16271_896 n3_16271_896 0.0
V28793 n1_16271_1079 n3_16271_1079 0.0
V28794 n1_16271_1112 n3_16271_1112 0.0
V28795 n1_16271_1295 n3_16271_1295 0.0
V28796 n1_16271_1328 n3_16271_1328 0.0
V28797 n1_16271_1511 n3_16271_1511 0.0
V28798 n1_16271_1544 n3_16271_1544 0.0
V28799 n1_16271_1727 n3_16271_1727 0.0
V28800 n1_16271_1760 n3_16271_1760 0.0
V28801 n1_16271_1894 n3_16271_1894 0.0
V28802 n1_16271_1943 n3_16271_1943 0.0
V28803 n1_16271_1976 n3_16271_1976 0.0
V28804 n1_16271_2159 n3_16271_2159 0.0
V28805 n1_16271_2192 n3_16271_2192 0.0
V28806 n1_16271_2375 n3_16271_2375 0.0
V28807 n1_16271_2408 n3_16271_2408 0.0
V28808 n1_16271_2445 n3_16271_2445 0.0
V28809 n1_16271_2542 n3_16271_2542 0.0
V28810 n1_16271_2543 n3_16271_2543 0.0
V28811 n1_16271_2591 n3_16271_2591 0.0
V28812 n1_16271_2624 n3_16271_2624 0.0
V28813 n1_16271_2807 n3_16271_2807 0.0
V28814 n1_16271_2840 n3_16271_2840 0.0
V28815 n1_16271_2877 n3_16271_2877 0.0
V28816 n1_16271_2974 n3_16271_2974 0.0
V28817 n1_16271_3023 n3_16271_3023 0.0
V28818 n1_16271_3056 n3_16271_3056 0.0
V28819 n1_16271_3239 n3_16271_3239 0.0
V28820 n1_16271_3272 n3_16271_3272 0.0
V28821 n1_16271_3406 n3_16271_3406 0.0
V28822 n1_16271_3455 n3_16271_3455 0.0
V28823 n1_16271_3488 n3_16271_3488 0.0
V28824 n1_16271_3671 n3_16271_3671 0.0
V28825 n1_16271_3704 n3_16271_3704 0.0
V28826 n1_16271_3887 n3_16271_3887 0.0
V28827 n1_16271_3920 n3_16271_3920 0.0
V28828 n1_16271_4103 n3_16271_4103 0.0
V28829 n1_16271_4136 n3_16271_4136 0.0
V28830 n1_16271_4319 n3_16271_4319 0.0
V28831 n1_16271_4352 n3_16271_4352 0.0
V28832 n1_16271_4486 n3_16271_4486 0.0
V28833 n1_16271_4535 n3_16271_4535 0.0
V28834 n1_16271_4568 n3_16271_4568 0.0
V28835 n1_16271_4702 n3_16271_4702 0.0
V28836 n1_16271_4751 n3_16271_4751 0.0
V28837 n1_16271_4784 n3_16271_4784 0.0
V28838 n1_16271_4919 n3_16271_4919 0.0
V28839 n1_16271_5000 n3_16271_5000 0.0
V28840 n1_16271_5134 n3_16271_5134 0.0
V28841 n1_16271_5183 n3_16271_5183 0.0
V28842 n1_16271_5216 n3_16271_5216 0.0
V28843 n1_16271_5253 n3_16271_5253 0.0
V28844 n1_16271_5350 n3_16271_5350 0.0
V28845 n1_16271_5399 n3_16271_5399 0.0
V28846 n1_16271_5432 n3_16271_5432 0.0
V28847 n1_16271_5566 n3_16271_5566 0.0
V28848 n1_16271_5615 n3_16271_5615 0.0
V28849 n1_16271_5648 n3_16271_5648 0.0
V28850 n1_16271_5831 n3_16271_5831 0.0
V28851 n1_16271_5864 n3_16271_5864 0.0
V28852 n1_16271_6047 n3_16271_6047 0.0
V28853 n1_16271_6080 n3_16271_6080 0.0
V28854 n1_16271_6263 n3_16271_6263 0.0
V28855 n1_16271_6296 n3_16271_6296 0.0
V28856 n1_16271_6333 n3_16271_6333 0.0
V28857 n1_16271_6430 n3_16271_6430 0.0
V28858 n1_16271_6479 n3_16271_6479 0.0
V28859 n1_16271_6512 n3_16271_6512 0.0
V28860 n1_16271_6695 n3_16271_6695 0.0
V28861 n1_16271_6728 n3_16271_6728 0.0
V28862 n1_16271_6911 n3_16271_6911 0.0
V28863 n1_16271_6944 n3_16271_6944 0.0
V28864 n1_16271_7127 n3_16271_7127 0.0
V28865 n1_16271_7160 n3_16271_7160 0.0
V28866 n1_16271_7343 n3_16271_7343 0.0
V28867 n1_16271_7376 n3_16271_7376 0.0
V28868 n1_16271_7559 n3_16271_7559 0.0
V28869 n1_16271_7592 n3_16271_7592 0.0
V28870 n1_16271_7775 n3_16271_7775 0.0
V28871 n1_16271_7808 n3_16271_7808 0.0
V28872 n1_16271_7845 n3_16271_7845 0.0
V28873 n1_16271_7942 n3_16271_7942 0.0
V28874 n1_16271_7991 n3_16271_7991 0.0
V28875 n1_16271_8024 n3_16271_8024 0.0
V28876 n1_16271_8207 n3_16271_8207 0.0
V28877 n1_16271_8240 n3_16271_8240 0.0
V28878 n1_16271_8423 n3_16271_8423 0.0
V28879 n1_16271_8456 n3_16271_8456 0.0
V28880 n1_16271_8639 n3_16271_8639 0.0
V28881 n1_16271_8672 n3_16271_8672 0.0
V28882 n1_16271_8855 n3_16271_8855 0.0
V28883 n1_16271_8888 n3_16271_8888 0.0
V28884 n1_16271_8925 n3_16271_8925 0.0
V28885 n1_16271_9022 n3_16271_9022 0.0
V28886 n1_16271_9071 n3_16271_9071 0.0
V28887 n1_16271_9104 n3_16271_9104 0.0
V28888 n1_16271_9287 n3_16271_9287 0.0
V28889 n1_16271_9320 n3_16271_9320 0.0
V28890 n1_16271_9503 n3_16271_9503 0.0
V28891 n1_16271_9536 n3_16271_9536 0.0
V28892 n1_16271_9719 n3_16271_9719 0.0
V28893 n1_16271_9752 n3_16271_9752 0.0
V28894 n1_16271_9935 n3_16271_9935 0.0
V28895 n1_16271_9968 n3_16271_9968 0.0
V28896 n1_16271_10005 n3_16271_10005 0.0
V28897 n1_16271_10102 n3_16271_10102 0.0
V28898 n1_16271_10151 n3_16271_10151 0.0
V28899 n1_16271_10184 n3_16271_10184 0.0
V28900 n1_16271_10367 n3_16271_10367 0.0
V28901 n1_16271_10400 n3_16271_10400 0.0
V28902 n1_16271_10616 n3_16271_10616 0.0
V28903 n1_16271_10799 n3_16271_10799 0.0
V28904 n1_16271_10832 n3_16271_10832 0.0
V28905 n1_16271_11015 n3_16271_11015 0.0
V28906 n1_16271_11048 n3_16271_11048 0.0
V28907 n1_16271_11196 n3_16271_11196 0.0
V28908 n1_16271_11204 n3_16271_11204 0.0
V28909 n1_16271_11231 n3_16271_11231 0.0
V28910 n1_16271_11264 n3_16271_11264 0.0
V28911 n1_16271_11447 n3_16271_11447 0.0
V28912 n1_16271_11480 n3_16271_11480 0.0
V28913 n1_16271_11663 n3_16271_11663 0.0
V28914 n1_16271_11696 n3_16271_11696 0.0
V28915 n1_16271_11879 n3_16271_11879 0.0
V28916 n1_16271_11912 n3_16271_11912 0.0
V28917 n1_16271_12095 n3_16271_12095 0.0
V28918 n1_16271_12128 n3_16271_12128 0.0
V28919 n1_16271_12276 n3_16271_12276 0.0
V28920 n1_16271_12284 n3_16271_12284 0.0
V28921 n1_16271_12311 n3_16271_12311 0.0
V28922 n1_16271_12344 n3_16271_12344 0.0
V28923 n1_16271_12527 n3_16271_12527 0.0
V28924 n1_16271_12560 n3_16271_12560 0.0
V28925 n1_16271_12743 n3_16271_12743 0.0
V28926 n1_16271_12776 n3_16271_12776 0.0
V28927 n1_16271_12959 n3_16271_12959 0.0
V28928 n1_16271_12992 n3_16271_12992 0.0
V28929 n1_16271_13175 n3_16271_13175 0.0
V28930 n1_16271_13208 n3_16271_13208 0.0
V28931 n1_16271_13391 n3_16271_13391 0.0
V28932 n1_16271_13424 n3_16271_13424 0.0
V28933 n1_16271_13607 n3_16271_13607 0.0
V28934 n1_16271_13640 n3_16271_13640 0.0
V28935 n1_16271_13788 n3_16271_13788 0.0
V28936 n1_16271_13823 n3_16271_13823 0.0
V28937 n1_16271_13856 n3_16271_13856 0.0
V28938 n1_16271_14039 n3_16271_14039 0.0
V28939 n1_16271_14072 n3_16271_14072 0.0
V28940 n1_16271_14255 n3_16271_14255 0.0
V28941 n1_16271_14288 n3_16271_14288 0.0
V28942 n1_16271_14471 n3_16271_14471 0.0
V28943 n1_16271_14504 n3_16271_14504 0.0
V28944 n1_16271_14652 n3_16271_14652 0.0
V28945 n1_16271_14687 n3_16271_14687 0.0
V28946 n1_16271_14720 n3_16271_14720 0.0
V28947 n1_16271_14903 n3_16271_14903 0.0
V28948 n1_16271_14936 n3_16271_14936 0.0
V28949 n1_16271_15084 n3_16271_15084 0.0
V28950 n1_16271_15119 n3_16271_15119 0.0
V28951 n1_16271_15152 n3_16271_15152 0.0
V28952 n1_16271_15300 n3_16271_15300 0.0
V28953 n1_16271_15335 n3_16271_15335 0.0
V28954 n1_16271_15368 n3_16271_15368 0.0
V28955 n1_16271_15551 n3_16271_15551 0.0
V28956 n1_16271_15584 n3_16271_15584 0.0
V28957 n1_16271_15740 n3_16271_15740 0.0
V28958 n1_16271_15767 n3_16271_15767 0.0
V28959 n1_16271_15800 n3_16271_15800 0.0
V28960 n1_16271_15983 n3_16271_15983 0.0
V28961 n1_16271_16016 n3_16271_16016 0.0
V28962 n1_16271_16199 n3_16271_16199 0.0
V28963 n1_16271_16415 n3_16271_16415 0.0
V28964 n1_16271_16448 n3_16271_16448 0.0
V28965 n1_16271_16604 n3_16271_16604 0.0
V28966 n1_16271_16631 n3_16271_16631 0.0
V28967 n1_16271_16664 n3_16271_16664 0.0
V28968 n1_16271_16798 n3_16271_16798 0.0
V28969 n1_16271_16820 n3_16271_16820 0.0
V28970 n1_16271_16847 n3_16271_16847 0.0
V28971 n1_16271_16880 n3_16271_16880 0.0
V28972 n1_16271_17063 n3_16271_17063 0.0
V28973 n1_16271_17096 n3_16271_17096 0.0
V28974 n1_16271_17252 n3_16271_17252 0.0
V28975 n1_16271_17279 n3_16271_17279 0.0
V28976 n1_16271_17312 n3_16271_17312 0.0
V28977 n1_16271_17495 n3_16271_17495 0.0
V28978 n1_16271_17528 n3_16271_17528 0.0
V28979 n1_16271_17676 n3_16271_17676 0.0
V28980 n1_16271_17684 n3_16271_17684 0.0
V28981 n1_16271_17711 n3_16271_17711 0.0
V28982 n1_16271_17744 n3_16271_17744 0.0
V28983 n1_16271_17927 n3_16271_17927 0.0
V28984 n1_16271_17960 n3_16271_17960 0.0
V28985 n1_16271_18143 n3_16271_18143 0.0
V28986 n1_16271_18176 n3_16271_18176 0.0
V28987 n1_16271_18332 n3_16271_18332 0.0
V28988 n1_16271_18359 n3_16271_18359 0.0
V28989 n1_16271_18392 n3_16271_18392 0.0
V28990 n1_16271_18527 n3_16271_18527 0.0
V28991 n1_16271_18575 n3_16271_18575 0.0
V28992 n1_16271_18608 n3_16271_18608 0.0
V28993 n1_16271_18764 n3_16271_18764 0.0
V28994 n1_16271_18791 n3_16271_18791 0.0
V28995 n1_16271_18824 n3_16271_18824 0.0
V28996 n1_16271_19007 n3_16271_19007 0.0
V28997 n1_16271_19040 n3_16271_19040 0.0
V28998 n1_16271_19196 n3_16271_19196 0.0
V28999 n1_16271_19223 n3_16271_19223 0.0
V29000 n1_16271_19256 n3_16271_19256 0.0
V29001 n1_16271_19412 n3_16271_19412 0.0
V29002 n1_16271_19439 n3_16271_19439 0.0
V29003 n1_16271_19472 n3_16271_19472 0.0
V29004 n1_16271_19655 n3_16271_19655 0.0
V29005 n1_16271_19688 n3_16271_19688 0.0
V29006 n1_16271_19871 n3_16271_19871 0.0
V29007 n1_16271_19904 n3_16271_19904 0.0
V29008 n1_16271_20087 n3_16271_20087 0.0
V29009 n1_16271_20120 n3_16271_20120 0.0
V29010 n1_16271_20303 n3_16271_20303 0.0
V29011 n1_16271_20336 n3_16271_20336 0.0
V29012 n1_16271_20519 n3_16271_20519 0.0
V29013 n1_16271_20552 n3_16271_20552 0.0
V29014 n1_16271_20687 n3_16271_20687 0.0
V29015 n1_16271_20768 n3_16271_20768 0.0
V29016 n1_16271_20951 n3_16271_20951 0.0
V29017 n1_16271_20984 n3_16271_20984 0.0
V29018 n1_16364_215 n3_16364_215 0.0
V29019 n1_16364_248 n3_16364_248 0.0
V29020 n1_16364_383 n3_16364_383 0.0
V29021 n1_16364_431 n3_16364_431 0.0
V29022 n1_16364_464 n3_16364_464 0.0
V29023 n1_16364_647 n3_16364_647 0.0
V29024 n1_16364_680 n3_16364_680 0.0
V29025 n1_16364_863 n3_16364_863 0.0
V29026 n1_16364_896 n3_16364_896 0.0
V29027 n1_16364_1079 n3_16364_1079 0.0
V29028 n1_16364_1112 n3_16364_1112 0.0
V29029 n1_16364_1295 n3_16364_1295 0.0
V29030 n1_16364_1328 n3_16364_1328 0.0
V29031 n1_16364_1511 n3_16364_1511 0.0
V29032 n1_16364_1544 n3_16364_1544 0.0
V29033 n1_16364_1727 n3_16364_1727 0.0
V29034 n1_16364_1760 n3_16364_1760 0.0
V29035 n1_16364_1894 n3_16364_1894 0.0
V29036 n1_16364_1943 n3_16364_1943 0.0
V29037 n1_16364_1976 n3_16364_1976 0.0
V29038 n1_16364_2159 n3_16364_2159 0.0
V29039 n1_16364_2192 n3_16364_2192 0.0
V29040 n1_16364_2375 n3_16364_2375 0.0
V29041 n1_16364_2408 n3_16364_2408 0.0
V29042 n1_16364_2445 n3_16364_2445 0.0
V29043 n1_16364_2542 n3_16364_2542 0.0
V29044 n1_16364_2543 n3_16364_2543 0.0
V29045 n1_16364_2591 n3_16364_2591 0.0
V29046 n1_16364_2624 n3_16364_2624 0.0
V29047 n1_16364_18527 n3_16364_18527 0.0
V29048 n1_16364_18575 n3_16364_18575 0.0
V29049 n1_16364_18608 n3_16364_18608 0.0
V29050 n1_16364_18791 n3_16364_18791 0.0
V29051 n1_16364_18824 n3_16364_18824 0.0
V29052 n1_16364_19007 n3_16364_19007 0.0
V29053 n1_16364_19040 n3_16364_19040 0.0
V29054 n1_16364_19196 n3_16364_19196 0.0
V29055 n1_16364_19223 n3_16364_19223 0.0
V29056 n1_16364_19256 n3_16364_19256 0.0
V29057 n1_16364_19439 n3_16364_19439 0.0
V29058 n1_16364_19472 n3_16364_19472 0.0
V29059 n1_16364_19655 n3_16364_19655 0.0
V29060 n1_16364_19688 n3_16364_19688 0.0
V29061 n1_16364_19871 n3_16364_19871 0.0
V29062 n1_16364_19904 n3_16364_19904 0.0
V29063 n1_16364_20087 n3_16364_20087 0.0
V29064 n1_16364_20120 n3_16364_20120 0.0
V29065 n1_16364_20303 n3_16364_20303 0.0
V29066 n1_16364_20336 n3_16364_20336 0.0
V29067 n1_16364_20519 n3_16364_20519 0.0
V29068 n1_16364_20552 n3_16364_20552 0.0
V29069 n1_16364_20687 n3_16364_20687 0.0
V29070 n1_16364_20735 n3_16364_20735 0.0
V29071 n1_16364_20768 n3_16364_20768 0.0
V29072 n1_16364_20951 n3_16364_20951 0.0
V29073 n1_16364_20984 n3_16364_20984 0.0
V29074 n1_18150_215 n3_18150_215 0.0
V29075 n1_18150_248 n3_18150_248 0.0
V29076 n1_18150_383 n3_18150_383 0.0
V29077 n1_18150_431 n3_18150_431 0.0
V29078 n1_18150_464 n3_18150_464 0.0
V29079 n1_18150_647 n3_18150_647 0.0
V29080 n1_18150_680 n3_18150_680 0.0
V29081 n1_18150_863 n3_18150_863 0.0
V29082 n1_18150_896 n3_18150_896 0.0
V29083 n1_18150_1079 n3_18150_1079 0.0
V29084 n1_18150_1112 n3_18150_1112 0.0
V29085 n1_18150_1295 n3_18150_1295 0.0
V29086 n1_18150_1328 n3_18150_1328 0.0
V29087 n1_18150_1511 n3_18150_1511 0.0
V29088 n1_18150_1544 n3_18150_1544 0.0
V29089 n1_18150_1727 n3_18150_1727 0.0
V29090 n1_18150_1760 n3_18150_1760 0.0
V29091 n1_18150_1894 n3_18150_1894 0.0
V29092 n1_18150_1943 n3_18150_1943 0.0
V29093 n1_18150_1976 n3_18150_1976 0.0
V29094 n1_18150_2159 n3_18150_2159 0.0
V29095 n1_18150_2192 n3_18150_2192 0.0
V29096 n1_18150_2375 n3_18150_2375 0.0
V29097 n1_18150_2408 n3_18150_2408 0.0
V29098 n1_18150_2542 n3_18150_2542 0.0
V29099 n1_18150_2543 n3_18150_2543 0.0
V29100 n1_18150_2591 n3_18150_2591 0.0
V29101 n1_18150_2624 n3_18150_2624 0.0
V29102 n1_18150_18527 n3_18150_18527 0.0
V29103 n1_18150_18575 n3_18150_18575 0.0
V29104 n1_18150_18608 n3_18150_18608 0.0
V29105 n1_18150_18791 n3_18150_18791 0.0
V29106 n1_18150_18824 n3_18150_18824 0.0
V29107 n1_18150_19007 n3_18150_19007 0.0
V29108 n1_18150_19040 n3_18150_19040 0.0
V29109 n1_18150_19223 n3_18150_19223 0.0
V29110 n1_18150_19256 n3_18150_19256 0.0
V29111 n1_18150_19439 n3_18150_19439 0.0
V29112 n1_18150_19472 n3_18150_19472 0.0
V29113 n1_18150_19655 n3_18150_19655 0.0
V29114 n1_18150_19688 n3_18150_19688 0.0
V29115 n1_18150_19871 n3_18150_19871 0.0
V29116 n1_18150_19904 n3_18150_19904 0.0
V29117 n1_18150_20087 n3_18150_20087 0.0
V29118 n1_18150_20120 n3_18150_20120 0.0
V29119 n1_18150_20303 n3_18150_20303 0.0
V29120 n1_18150_20336 n3_18150_20336 0.0
V29121 n1_18150_20519 n3_18150_20519 0.0
V29122 n1_18150_20552 n3_18150_20552 0.0
V29123 n1_18150_20687 n3_18150_20687 0.0
V29124 n1_18150_20735 n3_18150_20735 0.0
V29125 n1_18150_20768 n3_18150_20768 0.0
V29126 n1_18150_20951 n3_18150_20951 0.0
V29127 n1_18150_20984 n3_18150_20984 0.0
V29128 n1_18333_215 n3_18333_215 0.0
V29129 n1_18333_248 n3_18333_248 0.0
V29130 n1_18333_383 n3_18333_383 0.0
V29131 n1_18333_431 n3_18333_431 0.0
V29132 n1_18333_464 n3_18333_464 0.0
V29133 n1_18333_647 n3_18333_647 0.0
V29134 n1_18333_680 n3_18333_680 0.0
V29135 n1_18333_863 n3_18333_863 0.0
V29136 n1_18333_896 n3_18333_896 0.0
V29137 n1_18333_1079 n3_18333_1079 0.0
V29138 n1_18333_1112 n3_18333_1112 0.0
V29139 n1_18333_1295 n3_18333_1295 0.0
V29140 n1_18333_1328 n3_18333_1328 0.0
V29141 n1_18333_1727 n3_18333_1727 0.0
V29142 n1_18333_1760 n3_18333_1760 0.0
V29143 n1_18333_1894 n3_18333_1894 0.0
V29144 n1_18333_1943 n3_18333_1943 0.0
V29145 n1_18333_1976 n3_18333_1976 0.0
V29146 n1_18333_2110 n3_18333_2110 0.0
V29147 n1_18333_2159 n3_18333_2159 0.0
V29148 n1_18333_2192 n3_18333_2192 0.0
V29149 n1_18333_2375 n3_18333_2375 0.0
V29150 n1_18333_2408 n3_18333_2408 0.0
V29151 n1_18333_2542 n3_18333_2542 0.0
V29152 n1_18333_2543 n3_18333_2543 0.0
V29153 n1_18333_2591 n3_18333_2591 0.0
V29154 n1_18333_2624 n3_18333_2624 0.0
V29155 n1_18333_2807 n3_18333_2807 0.0
V29156 n1_18333_2840 n3_18333_2840 0.0
V29157 n1_18333_3023 n3_18333_3023 0.0
V29158 n1_18333_3056 n3_18333_3056 0.0
V29159 n1_18333_3239 n3_18333_3239 0.0
V29160 n1_18333_3272 n3_18333_3272 0.0
V29161 n1_18333_3406 n3_18333_3406 0.0
V29162 n1_18333_3455 n3_18333_3455 0.0
V29163 n1_18333_3488 n3_18333_3488 0.0
V29164 n1_18333_3671 n3_18333_3671 0.0
V29165 n1_18333_3704 n3_18333_3704 0.0
V29166 n1_18333_4103 n3_18333_4103 0.0
V29167 n1_18333_4136 n3_18333_4136 0.0
V29168 n1_18333_4319 n3_18333_4319 0.0
V29169 n1_18333_4352 n3_18333_4352 0.0
V29170 n1_18333_4486 n3_18333_4486 0.0
V29171 n1_18333_4535 n3_18333_4535 0.0
V29172 n1_18333_4568 n3_18333_4568 0.0
V29173 n1_18333_4702 n3_18333_4702 0.0
V29174 n1_18333_4751 n3_18333_4751 0.0
V29175 n1_18333_4784 n3_18333_4784 0.0
V29176 n1_18333_4920 n3_18333_4920 0.0
V29177 n1_18333_4967 n3_18333_4967 0.0
V29178 n1_18333_5000 n3_18333_5000 0.0
V29179 n1_18333_5134 n3_18333_5134 0.0
V29180 n1_18333_5183 n3_18333_5183 0.0
V29181 n1_18333_5216 n3_18333_5216 0.0
V29182 n1_18333_5253 n3_18333_5253 0.0
V29183 n1_18333_5350 n3_18333_5350 0.0
V29184 n1_18333_5399 n3_18333_5399 0.0
V29185 n1_18333_5432 n3_18333_5432 0.0
V29186 n1_18333_5566 n3_18333_5566 0.0
V29187 n1_18333_5615 n3_18333_5615 0.0
V29188 n1_18333_5648 n3_18333_5648 0.0
V29189 n1_18333_5831 n3_18333_5831 0.0
V29190 n1_18333_5864 n3_18333_5864 0.0
V29191 n1_18333_6263 n3_18333_6263 0.0
V29192 n1_18333_6296 n3_18333_6296 0.0
V29193 n1_18333_6333 n3_18333_6333 0.0
V29194 n1_18333_6430 n3_18333_6430 0.0
V29195 n1_18333_6479 n3_18333_6479 0.0
V29196 n1_18333_6512 n3_18333_6512 0.0
V29197 n1_18333_6695 n3_18333_6695 0.0
V29198 n1_18333_6728 n3_18333_6728 0.0
V29199 n1_18333_6911 n3_18333_6911 0.0
V29200 n1_18333_6944 n3_18333_6944 0.0
V29201 n1_18333_7127 n3_18333_7127 0.0
V29202 n1_18333_7160 n3_18333_7160 0.0
V29203 n1_18333_7343 n3_18333_7343 0.0
V29204 n1_18333_7376 n3_18333_7376 0.0
V29205 n1_18333_7559 n3_18333_7559 0.0
V29206 n1_18333_7592 n3_18333_7592 0.0
V29207 n1_18333_7775 n3_18333_7775 0.0
V29208 n1_18333_7808 n3_18333_7808 0.0
V29209 n1_18333_7845 n3_18333_7845 0.0
V29210 n1_18333_7942 n3_18333_7942 0.0
V29211 n1_18333_7991 n3_18333_7991 0.0
V29212 n1_18333_8024 n3_18333_8024 0.0
V29213 n1_18333_8207 n3_18333_8207 0.0
V29214 n1_18333_8240 n3_18333_8240 0.0
V29215 n1_18333_8456 n3_18333_8456 0.0
V29216 n1_18333_8639 n3_18333_8639 0.0
V29217 n1_18333_8672 n3_18333_8672 0.0
V29218 n1_18333_8855 n3_18333_8855 0.0
V29219 n1_18333_8888 n3_18333_8888 0.0
V29220 n1_18333_8925 n3_18333_8925 0.0
V29221 n1_18333_9022 n3_18333_9022 0.0
V29222 n1_18333_9071 n3_18333_9071 0.0
V29223 n1_18333_9104 n3_18333_9104 0.0
V29224 n1_18333_9287 n3_18333_9287 0.0
V29225 n1_18333_9320 n3_18333_9320 0.0
V29226 n1_18333_9503 n3_18333_9503 0.0
V29227 n1_18333_9536 n3_18333_9536 0.0
V29228 n1_18333_9719 n3_18333_9719 0.0
V29229 n1_18333_9752 n3_18333_9752 0.0
V29230 n1_18333_9935 n3_18333_9935 0.0
V29231 n1_18333_9968 n3_18333_9968 0.0
V29232 n1_18333_10005 n3_18333_10005 0.0
V29233 n1_18333_10102 n3_18333_10102 0.0
V29234 n1_18333_10151 n3_18333_10151 0.0
V29235 n1_18333_10184 n3_18333_10184 0.0
V29236 n1_18333_10367 n3_18333_10367 0.0
V29237 n1_18333_10400 n3_18333_10400 0.0
V29238 n1_18333_10799 n3_18333_10799 0.0
V29239 n1_18333_10832 n3_18333_10832 0.0
V29240 n1_18333_11015 n3_18333_11015 0.0
V29241 n1_18333_11048 n3_18333_11048 0.0
V29242 n1_18333_11196 n3_18333_11196 0.0
V29243 n1_18333_11231 n3_18333_11231 0.0
V29244 n1_18333_11264 n3_18333_11264 0.0
V29245 n1_18333_11447 n3_18333_11447 0.0
V29246 n1_18333_11480 n3_18333_11480 0.0
V29247 n1_18333_11663 n3_18333_11663 0.0
V29248 n1_18333_11696 n3_18333_11696 0.0
V29249 n1_18333_11879 n3_18333_11879 0.0
V29250 n1_18333_11912 n3_18333_11912 0.0
V29251 n1_18333_12095 n3_18333_12095 0.0
V29252 n1_18333_12128 n3_18333_12128 0.0
V29253 n1_18333_12284 n3_18333_12284 0.0
V29254 n1_18333_12311 n3_18333_12311 0.0
V29255 n1_18333_12344 n3_18333_12344 0.0
V29256 n1_18333_12527 n3_18333_12527 0.0
V29257 n1_18333_12560 n3_18333_12560 0.0
V29258 n1_18333_12743 n3_18333_12743 0.0
V29259 n1_18333_12959 n3_18333_12959 0.0
V29260 n1_18333_12992 n3_18333_12992 0.0
V29261 n1_18333_13175 n3_18333_13175 0.0
V29262 n1_18333_13208 n3_18333_13208 0.0
V29263 n1_18333_13391 n3_18333_13391 0.0
V29264 n1_18333_13424 n3_18333_13424 0.0
V29265 n1_18333_13607 n3_18333_13607 0.0
V29266 n1_18333_13640 n3_18333_13640 0.0
V29267 n1_18333_13788 n3_18333_13788 0.0
V29268 n1_18333_13796 n3_18333_13796 0.0
V29269 n1_18333_13823 n3_18333_13823 0.0
V29270 n1_18333_13856 n3_18333_13856 0.0
V29271 n1_18333_14039 n3_18333_14039 0.0
V29272 n1_18333_14072 n3_18333_14072 0.0
V29273 n1_18333_14255 n3_18333_14255 0.0
V29274 n1_18333_14288 n3_18333_14288 0.0
V29275 n1_18333_14471 n3_18333_14471 0.0
V29276 n1_18333_14504 n3_18333_14504 0.0
V29277 n1_18333_14652 n3_18333_14652 0.0
V29278 n1_18333_14660 n3_18333_14660 0.0
V29279 n1_18333_14687 n3_18333_14687 0.0
V29280 n1_18333_14720 n3_18333_14720 0.0
V29281 n1_18333_14903 n3_18333_14903 0.0
V29282 n1_18333_14936 n3_18333_14936 0.0
V29283 n1_18333_15308 n3_18333_15308 0.0
V29284 n1_18333_15335 n3_18333_15335 0.0
V29285 n1_18333_15368 n3_18333_15368 0.0
V29286 n1_18333_15551 n3_18333_15551 0.0
V29287 n1_18333_15584 n3_18333_15584 0.0
V29288 n1_18333_15740 n3_18333_15740 0.0
V29289 n1_18333_15767 n3_18333_15767 0.0
V29290 n1_18333_15800 n3_18333_15800 0.0
V29291 n1_18333_15983 n3_18333_15983 0.0
V29292 n1_18333_16016 n3_18333_16016 0.0
V29293 n1_18333_16199 n3_18333_16199 0.0
V29294 n1_18333_16232 n3_18333_16232 0.0
V29295 n1_18333_16415 n3_18333_16415 0.0
V29296 n1_18333_16448 n3_18333_16448 0.0
V29297 n1_18333_16631 n3_18333_16631 0.0
V29298 n1_18333_16664 n3_18333_16664 0.0
V29299 n1_18333_16812 n3_18333_16812 0.0
V29300 n1_18333_16820 n3_18333_16820 0.0
V29301 n1_18333_16847 n3_18333_16847 0.0
V29302 n1_18333_16880 n3_18333_16880 0.0
V29303 n1_18333_17063 n3_18333_17063 0.0
V29304 n1_18333_17096 n3_18333_17096 0.0
V29305 n1_18333_17230 n3_18333_17230 0.0
V29306 n1_18333_17495 n3_18333_17495 0.0
V29307 n1_18333_17528 n3_18333_17528 0.0
V29308 n1_18333_17711 n3_18333_17711 0.0
V29309 n1_18333_17744 n3_18333_17744 0.0
V29310 n1_18333_17900 n3_18333_17900 0.0
V29311 n1_18333_17927 n3_18333_17927 0.0
V29312 n1_18333_17960 n3_18333_17960 0.0
V29313 n1_18333_18143 n3_18333_18143 0.0
V29314 n1_18333_18176 n3_18333_18176 0.0
V29315 n1_18333_18359 n3_18333_18359 0.0
V29316 n1_18333_18392 n3_18333_18392 0.0
V29317 n1_18333_18527 n3_18333_18527 0.0
V29318 n1_18333_18575 n3_18333_18575 0.0
V29319 n1_18333_18608 n3_18333_18608 0.0
V29320 n1_18333_18791 n3_18333_18791 0.0
V29321 n1_18333_18824 n3_18333_18824 0.0
V29322 n1_18333_19007 n3_18333_19007 0.0
V29323 n1_18333_19040 n3_18333_19040 0.0
V29324 n1_18333_19223 n3_18333_19223 0.0
V29325 n1_18333_19256 n3_18333_19256 0.0
V29326 n1_18333_19439 n3_18333_19439 0.0
V29327 n1_18333_19472 n3_18333_19472 0.0
V29328 n1_18333_19871 n3_18333_19871 0.0
V29329 n1_18333_19904 n3_18333_19904 0.0
V29330 n1_18333_20087 n3_18333_20087 0.0
V29331 n1_18333_20120 n3_18333_20120 0.0
V29332 n1_18333_20303 n3_18333_20303 0.0
V29333 n1_18333_20336 n3_18333_20336 0.0
V29334 n1_18333_20519 n3_18333_20519 0.0
V29335 n1_18333_20552 n3_18333_20552 0.0
V29336 n1_18333_20687 n3_18333_20687 0.0
V29337 n1_18333_20735 n3_18333_20735 0.0
V29338 n1_18333_20768 n3_18333_20768 0.0
V29339 n1_18333_20951 n3_18333_20951 0.0
V29340 n1_18333_20984 n3_18333_20984 0.0
V29341 n1_18380_431 n3_18380_431 0.0
V29342 n1_18380_464 n3_18380_464 0.0
V29343 n1_18380_4920 n3_18380_4920 0.0
V29344 n1_18380_4967 n3_18380_4967 0.0
V29345 n1_18380_5000 n3_18380_5000 0.0
V29346 n1_18380_7160 n3_18380_7160 0.0
V29347 n1_18380_9503 n3_18380_9503 0.0
V29348 n1_18380_9536 n3_18380_9536 0.0
V29349 n1_18380_11663 n3_18380_11663 0.0
V29350 n1_18380_11696 n3_18380_11696 0.0
V29351 n1_18380_14039 n3_18380_14039 0.0
V29352 n1_18380_16199 n3_18380_16199 0.0
V29353 n1_18380_16232 n3_18380_16232 0.0
V29354 n1_18380_18392 n3_18380_18392 0.0
V29355 n1_18380_18527 n3_18380_18527 0.0
V29356 n1_18380_20687 n3_18380_20687 0.0
V29357 n1_18380_20735 n3_18380_20735 0.0
V29358 n1_18380_20768 n3_18380_20768 0.0
V29359 n1_18521_215 n3_18521_215 0.0
V29360 n1_18521_248 n3_18521_248 0.0
V29361 n1_18521_383 n3_18521_383 0.0
V29362 n1_18521_431 n3_18521_431 0.0
V29363 n1_18521_647 n3_18521_647 0.0
V29364 n1_18521_680 n3_18521_680 0.0
V29365 n1_18521_863 n3_18521_863 0.0
V29366 n1_18521_896 n3_18521_896 0.0
V29367 n1_18521_1079 n3_18521_1079 0.0
V29368 n1_18521_1112 n3_18521_1112 0.0
V29369 n1_18521_1295 n3_18521_1295 0.0
V29370 n1_18521_1328 n3_18521_1328 0.0
V29371 n1_18521_1511 n3_18521_1511 0.0
V29372 n1_18521_1544 n3_18521_1544 0.0
V29373 n1_18521_1727 n3_18521_1727 0.0
V29374 n1_18521_1760 n3_18521_1760 0.0
V29375 n1_18521_1894 n3_18521_1894 0.0
V29376 n1_18521_1943 n3_18521_1943 0.0
V29377 n1_18521_1976 n3_18521_1976 0.0
V29378 n1_18521_2110 n3_18521_2110 0.0
V29379 n1_18521_2159 n3_18521_2159 0.0
V29380 n1_18521_2192 n3_18521_2192 0.0
V29381 n1_18521_2375 n3_18521_2375 0.0
V29382 n1_18521_2408 n3_18521_2408 0.0
V29383 n1_18521_2542 n3_18521_2542 0.0
V29384 n1_18521_2543 n3_18521_2543 0.0
V29385 n1_18521_2591 n3_18521_2591 0.0
V29386 n1_18521_2624 n3_18521_2624 0.0
V29387 n1_18521_2807 n3_18521_2807 0.0
V29388 n1_18521_2840 n3_18521_2840 0.0
V29389 n1_18521_3023 n3_18521_3023 0.0
V29390 n1_18521_3056 n3_18521_3056 0.0
V29391 n1_18521_3239 n3_18521_3239 0.0
V29392 n1_18521_3272 n3_18521_3272 0.0
V29393 n1_18521_3406 n3_18521_3406 0.0
V29394 n1_18521_3455 n3_18521_3455 0.0
V29395 n1_18521_3488 n3_18521_3488 0.0
V29396 n1_18521_3671 n3_18521_3671 0.0
V29397 n1_18521_3704 n3_18521_3704 0.0
V29398 n1_18521_3887 n3_18521_3887 0.0
V29399 n1_18521_3920 n3_18521_3920 0.0
V29400 n1_18521_4103 n3_18521_4103 0.0
V29401 n1_18521_4136 n3_18521_4136 0.0
V29402 n1_18521_4319 n3_18521_4319 0.0
V29403 n1_18521_4352 n3_18521_4352 0.0
V29404 n1_18521_4486 n3_18521_4486 0.0
V29405 n1_18521_4535 n3_18521_4535 0.0
V29406 n1_18521_4568 n3_18521_4568 0.0
V29407 n1_18521_4702 n3_18521_4702 0.0
V29408 n1_18521_4751 n3_18521_4751 0.0
V29409 n1_18521_4784 n3_18521_4784 0.0
V29410 n1_18521_4920 n3_18521_4920 0.0
V29411 n1_18521_5000 n3_18521_5000 0.0
V29412 n1_18521_5134 n3_18521_5134 0.0
V29413 n1_18521_5183 n3_18521_5183 0.0
V29414 n1_18521_5216 n3_18521_5216 0.0
V29415 n1_18521_5253 n3_18521_5253 0.0
V29416 n1_18521_5350 n3_18521_5350 0.0
V29417 n1_18521_5399 n3_18521_5399 0.0
V29418 n1_18521_5432 n3_18521_5432 0.0
V29419 n1_18521_5566 n3_18521_5566 0.0
V29420 n1_18521_5615 n3_18521_5615 0.0
V29421 n1_18521_5648 n3_18521_5648 0.0
V29422 n1_18521_5831 n3_18521_5831 0.0
V29423 n1_18521_5864 n3_18521_5864 0.0
V29424 n1_18521_6047 n3_18521_6047 0.0
V29425 n1_18521_6080 n3_18521_6080 0.0
V29426 n1_18521_6263 n3_18521_6263 0.0
V29427 n1_18521_6296 n3_18521_6296 0.0
V29428 n1_18521_6333 n3_18521_6333 0.0
V29429 n1_18521_6430 n3_18521_6430 0.0
V29430 n1_18521_6479 n3_18521_6479 0.0
V29431 n1_18521_6512 n3_18521_6512 0.0
V29432 n1_18521_6695 n3_18521_6695 0.0
V29433 n1_18521_6728 n3_18521_6728 0.0
V29434 n1_18521_6911 n3_18521_6911 0.0
V29435 n1_18521_6944 n3_18521_6944 0.0
V29436 n1_18521_7127 n3_18521_7127 0.0
V29437 n1_18521_7160 n3_18521_7160 0.0
V29438 n1_18521_7343 n3_18521_7343 0.0
V29439 n1_18521_7376 n3_18521_7376 0.0
V29440 n1_18521_7559 n3_18521_7559 0.0
V29441 n1_18521_7592 n3_18521_7592 0.0
V29442 n1_18521_7775 n3_18521_7775 0.0
V29443 n1_18521_7808 n3_18521_7808 0.0
V29444 n1_18521_7845 n3_18521_7845 0.0
V29445 n1_18521_7942 n3_18521_7942 0.0
V29446 n1_18521_7991 n3_18521_7991 0.0
V29447 n1_18521_8024 n3_18521_8024 0.0
V29448 n1_18521_8207 n3_18521_8207 0.0
V29449 n1_18521_8240 n3_18521_8240 0.0
V29450 n1_18521_8423 n3_18521_8423 0.0
V29451 n1_18521_8456 n3_18521_8456 0.0
V29452 n1_18521_8639 n3_18521_8639 0.0
V29453 n1_18521_8672 n3_18521_8672 0.0
V29454 n1_18521_8855 n3_18521_8855 0.0
V29455 n1_18521_8888 n3_18521_8888 0.0
V29456 n1_18521_8925 n3_18521_8925 0.0
V29457 n1_18521_9022 n3_18521_9022 0.0
V29458 n1_18521_9071 n3_18521_9071 0.0
V29459 n1_18521_9104 n3_18521_9104 0.0
V29460 n1_18521_9287 n3_18521_9287 0.0
V29461 n1_18521_9320 n3_18521_9320 0.0
V29462 n1_18521_9503 n3_18521_9503 0.0
V29463 n1_18521_9536 n3_18521_9536 0.0
V29464 n1_18521_9719 n3_18521_9719 0.0
V29465 n1_18521_9752 n3_18521_9752 0.0
V29466 n1_18521_9935 n3_18521_9935 0.0
V29467 n1_18521_9968 n3_18521_9968 0.0
V29468 n1_18521_10005 n3_18521_10005 0.0
V29469 n1_18521_10102 n3_18521_10102 0.0
V29470 n1_18521_10151 n3_18521_10151 0.0
V29471 n1_18521_10184 n3_18521_10184 0.0
V29472 n1_18521_10367 n3_18521_10367 0.0
V29473 n1_18521_10400 n3_18521_10400 0.0
V29474 n1_18521_10616 n3_18521_10616 0.0
V29475 n1_18521_10799 n3_18521_10799 0.0
V29476 n1_18521_10832 n3_18521_10832 0.0
V29477 n1_18521_11015 n3_18521_11015 0.0
V29478 n1_18521_11048 n3_18521_11048 0.0
V29479 n1_18521_11196 n3_18521_11196 0.0
V29480 n1_18521_11231 n3_18521_11231 0.0
V29481 n1_18521_11264 n3_18521_11264 0.0
V29482 n1_18521_11447 n3_18521_11447 0.0
V29483 n1_18521_11480 n3_18521_11480 0.0
V29484 n1_18521_11663 n3_18521_11663 0.0
V29485 n1_18521_11696 n3_18521_11696 0.0
V29486 n1_18521_11879 n3_18521_11879 0.0
V29487 n1_18521_11912 n3_18521_11912 0.0
V29488 n1_18521_12095 n3_18521_12095 0.0
V29489 n1_18521_12128 n3_18521_12128 0.0
V29490 n1_18521_12284 n3_18521_12284 0.0
V29491 n1_18521_12311 n3_18521_12311 0.0
V29492 n1_18521_12344 n3_18521_12344 0.0
V29493 n1_18521_12527 n3_18521_12527 0.0
V29494 n1_18521_12560 n3_18521_12560 0.0
V29495 n1_18521_12743 n3_18521_12743 0.0
V29496 n1_18521_12776 n3_18521_12776 0.0
V29497 n1_18521_12959 n3_18521_12959 0.0
V29498 n1_18521_12992 n3_18521_12992 0.0
V29499 n1_18521_13175 n3_18521_13175 0.0
V29500 n1_18521_13208 n3_18521_13208 0.0
V29501 n1_18521_13391 n3_18521_13391 0.0
V29502 n1_18521_13424 n3_18521_13424 0.0
V29503 n1_18521_13607 n3_18521_13607 0.0
V29504 n1_18521_13640 n3_18521_13640 0.0
V29505 n1_18521_13788 n3_18521_13788 0.0
V29506 n1_18521_13796 n3_18521_13796 0.0
V29507 n1_18521_13823 n3_18521_13823 0.0
V29508 n1_18521_13856 n3_18521_13856 0.0
V29509 n1_18521_14039 n3_18521_14039 0.0
V29510 n1_18521_14072 n3_18521_14072 0.0
V29511 n1_18521_14255 n3_18521_14255 0.0
V29512 n1_18521_14288 n3_18521_14288 0.0
V29513 n1_18521_14471 n3_18521_14471 0.0
V29514 n1_18521_14504 n3_18521_14504 0.0
V29515 n1_18521_14652 n3_18521_14652 0.0
V29516 n1_18521_14660 n3_18521_14660 0.0
V29517 n1_18521_14687 n3_18521_14687 0.0
V29518 n1_18521_14720 n3_18521_14720 0.0
V29519 n1_18521_14903 n3_18521_14903 0.0
V29520 n1_18521_14936 n3_18521_14936 0.0
V29521 n1_18521_15092 n3_18521_15092 0.0
V29522 n1_18521_15119 n3_18521_15119 0.0
V29523 n1_18521_15152 n3_18521_15152 0.0
V29524 n1_18521_15308 n3_18521_15308 0.0
V29525 n1_18521_15335 n3_18521_15335 0.0
V29526 n1_18521_15368 n3_18521_15368 0.0
V29527 n1_18521_15551 n3_18521_15551 0.0
V29528 n1_18521_15584 n3_18521_15584 0.0
V29529 n1_18521_15740 n3_18521_15740 0.0
V29530 n1_18521_15767 n3_18521_15767 0.0
V29531 n1_18521_15800 n3_18521_15800 0.0
V29532 n1_18521_15983 n3_18521_15983 0.0
V29533 n1_18521_16016 n3_18521_16016 0.0
V29534 n1_18521_16199 n3_18521_16199 0.0
V29535 n1_18521_16415 n3_18521_16415 0.0
V29536 n1_18521_16448 n3_18521_16448 0.0
V29537 n1_18521_16631 n3_18521_16631 0.0
V29538 n1_18521_16664 n3_18521_16664 0.0
V29539 n1_18521_16812 n3_18521_16812 0.0
V29540 n1_18521_16820 n3_18521_16820 0.0
V29541 n1_18521_16847 n3_18521_16847 0.0
V29542 n1_18521_16880 n3_18521_16880 0.0
V29543 n1_18521_17063 n3_18521_17063 0.0
V29544 n1_18521_17096 n3_18521_17096 0.0
V29545 n1_18521_17230 n3_18521_17230 0.0
V29546 n1_18521_17279 n3_18521_17279 0.0
V29547 n1_18521_17312 n3_18521_17312 0.0
V29548 n1_18521_17495 n3_18521_17495 0.0
V29549 n1_18521_17528 n3_18521_17528 0.0
V29550 n1_18521_17711 n3_18521_17711 0.0
V29551 n1_18521_17744 n3_18521_17744 0.0
V29552 n1_18521_17900 n3_18521_17900 0.0
V29553 n1_18521_17927 n3_18521_17927 0.0
V29554 n1_18521_17960 n3_18521_17960 0.0
V29555 n1_18521_18143 n3_18521_18143 0.0
V29556 n1_18521_18176 n3_18521_18176 0.0
V29557 n1_18521_18359 n3_18521_18359 0.0
V29558 n1_18521_18392 n3_18521_18392 0.0
V29559 n1_18521_18527 n3_18521_18527 0.0
V29560 n1_18521_18575 n3_18521_18575 0.0
V29561 n1_18521_18608 n3_18521_18608 0.0
V29562 n1_18521_18791 n3_18521_18791 0.0
V29563 n1_18521_18824 n3_18521_18824 0.0
V29564 n1_18521_19007 n3_18521_19007 0.0
V29565 n1_18521_19040 n3_18521_19040 0.0
V29566 n1_18521_19223 n3_18521_19223 0.0
V29567 n1_18521_19256 n3_18521_19256 0.0
V29568 n1_18521_19439 n3_18521_19439 0.0
V29569 n1_18521_19472 n3_18521_19472 0.0
V29570 n1_18521_19655 n3_18521_19655 0.0
V29571 n1_18521_19688 n3_18521_19688 0.0
V29572 n1_18521_19871 n3_18521_19871 0.0
V29573 n1_18521_19904 n3_18521_19904 0.0
V29574 n1_18521_20087 n3_18521_20087 0.0
V29575 n1_18521_20120 n3_18521_20120 0.0
V29576 n1_18521_20303 n3_18521_20303 0.0
V29577 n1_18521_20336 n3_18521_20336 0.0
V29578 n1_18521_20519 n3_18521_20519 0.0
V29579 n1_18521_20552 n3_18521_20552 0.0
V29580 n1_18521_20687 n3_18521_20687 0.0
V29581 n1_18521_20768 n3_18521_20768 0.0
V29582 n1_18521_20951 n3_18521_20951 0.0
V29583 n1_18521_20984 n3_18521_20984 0.0
V29584 n1_18614_215 n3_18614_215 0.0
V29585 n1_18614_248 n3_18614_248 0.0
V29586 n1_18614_383 n3_18614_383 0.0
V29587 n1_18614_431 n3_18614_431 0.0
V29588 n1_18614_464 n3_18614_464 0.0
V29589 n1_18614_647 n3_18614_647 0.0
V29590 n1_18614_680 n3_18614_680 0.0
V29591 n1_18614_863 n3_18614_863 0.0
V29592 n1_18614_896 n3_18614_896 0.0
V29593 n1_18614_1079 n3_18614_1079 0.0
V29594 n1_18614_1112 n3_18614_1112 0.0
V29595 n1_18614_1295 n3_18614_1295 0.0
V29596 n1_18614_1328 n3_18614_1328 0.0
V29597 n1_18614_1511 n3_18614_1511 0.0
V29598 n1_18614_1544 n3_18614_1544 0.0
V29599 n1_18614_1727 n3_18614_1727 0.0
V29600 n1_18614_1760 n3_18614_1760 0.0
V29601 n1_18614_1943 n3_18614_1943 0.0
V29602 n1_18614_1976 n3_18614_1976 0.0
V29603 n1_18614_2110 n3_18614_2110 0.0
V29604 n1_18614_2159 n3_18614_2159 0.0
V29605 n1_18614_2192 n3_18614_2192 0.0
V29606 n1_18614_2375 n3_18614_2375 0.0
V29607 n1_18614_2408 n3_18614_2408 0.0
V29608 n1_18614_2543 n3_18614_2543 0.0
V29609 n1_18614_2591 n3_18614_2591 0.0
V29610 n1_18614_2624 n3_18614_2624 0.0
V29611 n1_18614_18527 n3_18614_18527 0.0
V29612 n1_18614_18575 n3_18614_18575 0.0
V29613 n1_18614_18608 n3_18614_18608 0.0
V29614 n1_18614_18791 n3_18614_18791 0.0
V29615 n1_18614_18824 n3_18614_18824 0.0
V29616 n1_18614_19007 n3_18614_19007 0.0
V29617 n1_18614_19040 n3_18614_19040 0.0
V29618 n1_18614_19223 n3_18614_19223 0.0
V29619 n1_18614_19256 n3_18614_19256 0.0
V29620 n1_18614_19439 n3_18614_19439 0.0
V29621 n1_18614_19472 n3_18614_19472 0.0
V29622 n1_18614_19655 n3_18614_19655 0.0
V29623 n1_18614_19688 n3_18614_19688 0.0
V29624 n1_18614_19871 n3_18614_19871 0.0
V29625 n1_18614_19904 n3_18614_19904 0.0
V29626 n1_18614_20087 n3_18614_20087 0.0
V29627 n1_18614_20120 n3_18614_20120 0.0
V29628 n1_18614_20303 n3_18614_20303 0.0
V29629 n1_18614_20336 n3_18614_20336 0.0
V29630 n1_18614_20519 n3_18614_20519 0.0
V29631 n1_18614_20552 n3_18614_20552 0.0
V29632 n1_18614_20687 n3_18614_20687 0.0
V29633 n1_18614_20735 n3_18614_20735 0.0
V29634 n1_18614_20768 n3_18614_20768 0.0
V29635 n1_18614_20951 n3_18614_20951 0.0
V29636 n1_18614_20984 n3_18614_20984 0.0
V29637 n1_20583_215 n3_20583_215 0.0
V29638 n1_20583_248 n3_20583_248 0.0
V29639 n1_20583_383 n3_20583_383 0.0
V29640 n1_20583_431 n3_20583_431 0.0
V29641 n1_20583_464 n3_20583_464 0.0
V29642 n1_20583_647 n3_20583_647 0.0
V29643 n1_20583_680 n3_20583_680 0.0
V29644 n1_20583_863 n3_20583_863 0.0
V29645 n1_20583_896 n3_20583_896 0.0
V29646 n1_20583_1079 n3_20583_1079 0.0
V29647 n1_20583_1112 n3_20583_1112 0.0
V29648 n1_20583_1295 n3_20583_1295 0.0
V29649 n1_20583_1328 n3_20583_1328 0.0
V29650 n1_20583_1727 n3_20583_1727 0.0
V29651 n1_20583_1760 n3_20583_1760 0.0
V29652 n1_20583_1943 n3_20583_1943 0.0
V29653 n1_20583_1976 n3_20583_1976 0.0
V29654 n1_20583_2159 n3_20583_2159 0.0
V29655 n1_20583_2192 n3_20583_2192 0.0
V29656 n1_20583_2375 n3_20583_2375 0.0
V29657 n1_20583_2408 n3_20583_2408 0.0
V29658 n1_20583_2543 n3_20583_2543 0.0
V29659 n1_20583_2591 n3_20583_2591 0.0
V29660 n1_20583_2624 n3_20583_2624 0.0
V29661 n1_20583_2807 n3_20583_2807 0.0
V29662 n1_20583_2840 n3_20583_2840 0.0
V29663 n1_20583_3023 n3_20583_3023 0.0
V29664 n1_20583_3056 n3_20583_3056 0.0
V29665 n1_20583_3239 n3_20583_3239 0.0
V29666 n1_20583_3272 n3_20583_3272 0.0
V29667 n1_20583_3455 n3_20583_3455 0.0
V29668 n1_20583_3488 n3_20583_3488 0.0
V29669 n1_20583_3671 n3_20583_3671 0.0
V29670 n1_20583_3704 n3_20583_3704 0.0
V29671 n1_20583_4103 n3_20583_4103 0.0
V29672 n1_20583_4136 n3_20583_4136 0.0
V29673 n1_20583_4319 n3_20583_4319 0.0
V29674 n1_20583_4352 n3_20583_4352 0.0
V29675 n1_20583_4535 n3_20583_4535 0.0
V29676 n1_20583_4568 n3_20583_4568 0.0
V29677 n1_20583_4751 n3_20583_4751 0.0
V29678 n1_20583_4784 n3_20583_4784 0.0
V29679 n1_20583_4967 n3_20583_4967 0.0
V29680 n1_20583_5000 n3_20583_5000 0.0
V29681 n1_20583_5183 n3_20583_5183 0.0
V29682 n1_20583_5216 n3_20583_5216 0.0
V29683 n1_20583_5399 n3_20583_5399 0.0
V29684 n1_20583_5432 n3_20583_5432 0.0
V29685 n1_20583_5615 n3_20583_5615 0.0
V29686 n1_20583_5648 n3_20583_5648 0.0
V29687 n1_20583_5782 n3_20583_5782 0.0
V29688 n1_20583_5831 n3_20583_5831 0.0
V29689 n1_20583_5864 n3_20583_5864 0.0
V29690 n1_20583_6263 n3_20583_6263 0.0
V29691 n1_20583_6296 n3_20583_6296 0.0
V29692 n1_20583_6333 n3_20583_6333 0.0
V29693 n1_20583_6479 n3_20583_6479 0.0
V29694 n1_20583_6512 n3_20583_6512 0.0
V29695 n1_20583_6695 n3_20583_6695 0.0
V29696 n1_20583_6728 n3_20583_6728 0.0
V29697 n1_20583_6911 n3_20583_6911 0.0
V29698 n1_20583_6944 n3_20583_6944 0.0
V29699 n1_20583_7127 n3_20583_7127 0.0
V29700 n1_20583_7160 n3_20583_7160 0.0
V29701 n1_20583_7343 n3_20583_7343 0.0
V29702 n1_20583_7376 n3_20583_7376 0.0
V29703 n1_20583_7559 n3_20583_7559 0.0
V29704 n1_20583_7592 n3_20583_7592 0.0
V29705 n1_20583_7775 n3_20583_7775 0.0
V29706 n1_20583_7808 n3_20583_7808 0.0
V29707 n1_20583_7991 n3_20583_7991 0.0
V29708 n1_20583_8024 n3_20583_8024 0.0
V29709 n1_20583_8207 n3_20583_8207 0.0
V29710 n1_20583_8240 n3_20583_8240 0.0
V29711 n1_20583_8456 n3_20583_8456 0.0
V29712 n1_20583_8639 n3_20583_8639 0.0
V29713 n1_20583_8672 n3_20583_8672 0.0
V29714 n1_20583_8855 n3_20583_8855 0.0
V29715 n1_20583_8888 n3_20583_8888 0.0
V29716 n1_20583_9071 n3_20583_9071 0.0
V29717 n1_20583_9104 n3_20583_9104 0.0
V29718 n1_20583_9287 n3_20583_9287 0.0
V29719 n1_20583_9320 n3_20583_9320 0.0
V29720 n1_20583_9503 n3_20583_9503 0.0
V29721 n1_20583_9536 n3_20583_9536 0.0
V29722 n1_20583_9719 n3_20583_9719 0.0
V29723 n1_20583_9752 n3_20583_9752 0.0
V29724 n1_20583_9935 n3_20583_9935 0.0
V29725 n1_20583_9968 n3_20583_9968 0.0
V29726 n1_20583_10151 n3_20583_10151 0.0
V29727 n1_20583_10184 n3_20583_10184 0.0
V29728 n1_20583_10367 n3_20583_10367 0.0
V29729 n1_20583_10400 n3_20583_10400 0.0
V29730 n1_20583_10799 n3_20583_10799 0.0
V29731 n1_20583_10832 n3_20583_10832 0.0
V29732 n1_20583_11015 n3_20583_11015 0.0
V29733 n1_20583_11048 n3_20583_11048 0.0
V29734 n1_20583_11231 n3_20583_11231 0.0
V29735 n1_20583_11264 n3_20583_11264 0.0
V29736 n1_20583_11447 n3_20583_11447 0.0
V29737 n1_20583_11480 n3_20583_11480 0.0
V29738 n1_20583_11663 n3_20583_11663 0.0
V29739 n1_20583_11696 n3_20583_11696 0.0
V29740 n1_20583_11879 n3_20583_11879 0.0
V29741 n1_20583_11912 n3_20583_11912 0.0
V29742 n1_20583_12095 n3_20583_12095 0.0
V29743 n1_20583_12128 n3_20583_12128 0.0
V29744 n1_20583_12311 n3_20583_12311 0.0
V29745 n1_20583_12344 n3_20583_12344 0.0
V29746 n1_20583_12527 n3_20583_12527 0.0
V29747 n1_20583_12560 n3_20583_12560 0.0
V29748 n1_20583_12743 n3_20583_12743 0.0
V29749 n1_20583_12959 n3_20583_12959 0.0
V29750 n1_20583_12992 n3_20583_12992 0.0
V29751 n1_20583_13175 n3_20583_13175 0.0
V29752 n1_20583_13208 n3_20583_13208 0.0
V29753 n1_20583_13391 n3_20583_13391 0.0
V29754 n1_20583_13424 n3_20583_13424 0.0
V29755 n1_20583_13607 n3_20583_13607 0.0
V29756 n1_20583_13640 n3_20583_13640 0.0
V29757 n1_20583_13823 n3_20583_13823 0.0
V29758 n1_20583_13856 n3_20583_13856 0.0
V29759 n1_20583_14039 n3_20583_14039 0.0
V29760 n1_20583_14072 n3_20583_14072 0.0
V29761 n1_20583_14255 n3_20583_14255 0.0
V29762 n1_20583_14288 n3_20583_14288 0.0
V29763 n1_20583_14471 n3_20583_14471 0.0
V29764 n1_20583_14504 n3_20583_14504 0.0
V29765 n1_20583_14687 n3_20583_14687 0.0
V29766 n1_20583_14720 n3_20583_14720 0.0
V29767 n1_20583_14903 n3_20583_14903 0.0
V29768 n1_20583_14936 n3_20583_14936 0.0
V29769 n1_20583_15308 n3_20583_15308 0.0
V29770 n1_20583_15335 n3_20583_15335 0.0
V29771 n1_20583_15368 n3_20583_15368 0.0
V29772 n1_20583_15551 n3_20583_15551 0.0
V29773 n1_20583_15584 n3_20583_15584 0.0
V29774 n1_20583_15767 n3_20583_15767 0.0
V29775 n1_20583_15800 n3_20583_15800 0.0
V29776 n1_20583_15983 n3_20583_15983 0.0
V29777 n1_20583_16016 n3_20583_16016 0.0
V29778 n1_20583_16199 n3_20583_16199 0.0
V29779 n1_20583_16232 n3_20583_16232 0.0
V29780 n1_20583_16415 n3_20583_16415 0.0
V29781 n1_20583_16448 n3_20583_16448 0.0
V29782 n1_20583_16631 n3_20583_16631 0.0
V29783 n1_20583_16664 n3_20583_16664 0.0
V29784 n1_20583_16798 n3_20583_16798 0.0
V29785 n1_20583_16847 n3_20583_16847 0.0
V29786 n1_20583_16880 n3_20583_16880 0.0
V29787 n1_20583_17063 n3_20583_17063 0.0
V29788 n1_20583_17096 n3_20583_17096 0.0
V29789 n1_20583_17495 n3_20583_17495 0.0
V29790 n1_20583_17528 n3_20583_17528 0.0
V29791 n1_20583_17711 n3_20583_17711 0.0
V29792 n1_20583_17744 n3_20583_17744 0.0
V29793 n1_20583_17927 n3_20583_17927 0.0
V29794 n1_20583_17960 n3_20583_17960 0.0
V29795 n1_20583_18143 n3_20583_18143 0.0
V29796 n1_20583_18176 n3_20583_18176 0.0
V29797 n1_20583_18359 n3_20583_18359 0.0
V29798 n1_20583_18392 n3_20583_18392 0.0
V29799 n1_20583_18527 n3_20583_18527 0.0
V29800 n1_20583_18575 n3_20583_18575 0.0
V29801 n1_20583_18608 n3_20583_18608 0.0
V29802 n1_20583_18791 n3_20583_18791 0.0
V29803 n1_20583_18824 n3_20583_18824 0.0
V29804 n1_20583_19007 n3_20583_19007 0.0
V29805 n1_20583_19040 n3_20583_19040 0.0
V29806 n1_20583_19223 n3_20583_19223 0.0
V29807 n1_20583_19256 n3_20583_19256 0.0
V29808 n1_20583_19439 n3_20583_19439 0.0
V29809 n1_20583_19472 n3_20583_19472 0.0
V29810 n1_20583_19871 n3_20583_19871 0.0
V29811 n1_20583_19904 n3_20583_19904 0.0
V29812 n1_20583_20087 n3_20583_20087 0.0
V29813 n1_20583_20120 n3_20583_20120 0.0
V29814 n1_20583_20303 n3_20583_20303 0.0
V29815 n1_20583_20336 n3_20583_20336 0.0
V29816 n1_20583_20519 n3_20583_20519 0.0
V29817 n1_20583_20552 n3_20583_20552 0.0
V29818 n1_20583_20687 n3_20583_20687 0.0
V29819 n1_20583_20735 n3_20583_20735 0.0
V29820 n1_20583_20768 n3_20583_20768 0.0
V29821 n1_20583_20951 n3_20583_20951 0.0
V29822 n1_20583_20984 n3_20583_20984 0.0
V29823 n1_20630_431 n3_20630_431 0.0
V29824 n1_20630_464 n3_20630_464 0.0
V29825 n1_20630_4967 n3_20630_4967 0.0
V29826 n1_20630_5000 n3_20630_5000 0.0
V29827 n1_20630_7160 n3_20630_7160 0.0
V29828 n1_20630_9503 n3_20630_9503 0.0
V29829 n1_20630_9536 n3_20630_9536 0.0
V29830 n1_20630_11663 n3_20630_11663 0.0
V29831 n1_20630_11696 n3_20630_11696 0.0
V29832 n1_20630_14039 n3_20630_14039 0.0
V29833 n1_20630_16199 n3_20630_16199 0.0
V29834 n1_20630_16232 n3_20630_16232 0.0
V29835 n1_20630_18392 n3_20630_18392 0.0
V29836 n1_20630_18527 n3_20630_18527 0.0
V29837 n1_20630_20687 n3_20630_20687 0.0
V29838 n1_20630_20735 n3_20630_20735 0.0
V29839 n1_20630_20768 n3_20630_20768 0.0
V29840 n1_20771_647 n3_20771_647 0.0
V29841 n1_20771_680 n3_20771_680 0.0
V29842 n1_20771_863 n3_20771_863 0.0
V29843 n1_20771_896 n3_20771_896 0.0
V29844 n1_20771_1079 n3_20771_1079 0.0
V29845 n1_20771_1112 n3_20771_1112 0.0
V29846 n1_20771_1295 n3_20771_1295 0.0
V29847 n1_20771_1328 n3_20771_1328 0.0
V29848 n1_20771_1511 n3_20771_1511 0.0
V29849 n1_20771_1544 n3_20771_1544 0.0
V29850 n1_20771_1727 n3_20771_1727 0.0
V29851 n1_20771_1760 n3_20771_1760 0.0
V29852 n1_20771_1943 n3_20771_1943 0.0
V29853 n1_20771_1976 n3_20771_1976 0.0
V29854 n1_20771_2159 n3_20771_2159 0.0
V29855 n1_20771_2192 n3_20771_2192 0.0
V29856 n1_20771_2375 n3_20771_2375 0.0
V29857 n1_20771_2408 n3_20771_2408 0.0
V29858 n1_20771_2543 n3_20771_2543 0.0
V29859 n1_20771_2591 n3_20771_2591 0.0
V29860 n1_20771_2624 n3_20771_2624 0.0
V29861 n1_20771_2807 n3_20771_2807 0.0
V29862 n1_20771_2840 n3_20771_2840 0.0
V29863 n1_20771_3023 n3_20771_3023 0.0
V29864 n1_20771_3056 n3_20771_3056 0.0
V29865 n1_20771_3239 n3_20771_3239 0.0
V29866 n1_20771_3272 n3_20771_3272 0.0
V29867 n1_20771_3455 n3_20771_3455 0.0
V29868 n1_20771_3488 n3_20771_3488 0.0
V29869 n1_20771_3671 n3_20771_3671 0.0
V29870 n1_20771_3704 n3_20771_3704 0.0
V29871 n1_20771_3887 n3_20771_3887 0.0
V29872 n1_20771_3920 n3_20771_3920 0.0
V29873 n1_20771_4103 n3_20771_4103 0.0
V29874 n1_20771_4136 n3_20771_4136 0.0
V29875 n1_20771_4319 n3_20771_4319 0.0
V29876 n1_20771_4352 n3_20771_4352 0.0
V29877 n1_20771_4535 n3_20771_4535 0.0
V29878 n1_20771_4568 n3_20771_4568 0.0
V29879 n1_20771_4751 n3_20771_4751 0.0
V29880 n1_20771_4784 n3_20771_4784 0.0
V29881 n1_20771_5000 n3_20771_5000 0.0
V29882 n1_20771_5183 n3_20771_5183 0.0
V29883 n1_20771_5216 n3_20771_5216 0.0
V29884 n1_20771_5399 n3_20771_5399 0.0
V29885 n1_20771_5432 n3_20771_5432 0.0
V29886 n1_20771_5615 n3_20771_5615 0.0
V29887 n1_20771_5648 n3_20771_5648 0.0
V29888 n1_20771_5782 n3_20771_5782 0.0
V29889 n1_20771_5831 n3_20771_5831 0.0
V29890 n1_20771_5864 n3_20771_5864 0.0
V29891 n1_20771_6047 n3_20771_6047 0.0
V29892 n1_20771_6080 n3_20771_6080 0.0
V29893 n1_20771_6263 n3_20771_6263 0.0
V29894 n1_20771_6296 n3_20771_6296 0.0
V29895 n1_20771_6479 n3_20771_6479 0.0
V29896 n1_20771_6512 n3_20771_6512 0.0
V29897 n1_20771_6695 n3_20771_6695 0.0
V29898 n1_20771_6728 n3_20771_6728 0.0
V29899 n1_20771_6911 n3_20771_6911 0.0
V29900 n1_20771_6944 n3_20771_6944 0.0
V29901 n1_20771_7127 n3_20771_7127 0.0
V29902 n1_20771_7160 n3_20771_7160 0.0
V29903 n1_20771_7343 n3_20771_7343 0.0
V29904 n1_20771_7376 n3_20771_7376 0.0
V29905 n1_20771_7559 n3_20771_7559 0.0
V29906 n1_20771_7592 n3_20771_7592 0.0
V29907 n1_20771_7775 n3_20771_7775 0.0
V29908 n1_20771_7808 n3_20771_7808 0.0
V29909 n1_20771_7991 n3_20771_7991 0.0
V29910 n1_20771_8024 n3_20771_8024 0.0
V29911 n1_20771_8207 n3_20771_8207 0.0
V29912 n1_20771_8240 n3_20771_8240 0.0
V29913 n1_20771_8423 n3_20771_8423 0.0
V29914 n1_20771_8456 n3_20771_8456 0.0
V29915 n1_20771_8639 n3_20771_8639 0.0
V29916 n1_20771_8672 n3_20771_8672 0.0
V29917 n1_20771_8855 n3_20771_8855 0.0
V29918 n1_20771_8888 n3_20771_8888 0.0
V29919 n1_20771_9071 n3_20771_9071 0.0
V29920 n1_20771_9104 n3_20771_9104 0.0
V29921 n1_20771_9287 n3_20771_9287 0.0
V29922 n1_20771_9320 n3_20771_9320 0.0
V29923 n1_20771_9503 n3_20771_9503 0.0
V29924 n1_20771_9536 n3_20771_9536 0.0
V29925 n1_20771_9719 n3_20771_9719 0.0
V29926 n1_20771_9752 n3_20771_9752 0.0
V29927 n1_20771_9935 n3_20771_9935 0.0
V29928 n1_20771_9968 n3_20771_9968 0.0
V29929 n1_20771_10151 n3_20771_10151 0.0
V29930 n1_20771_10184 n3_20771_10184 0.0
V29931 n1_20771_10367 n3_20771_10367 0.0
V29932 n1_20771_10400 n3_20771_10400 0.0
V29933 n1_20771_10616 n3_20771_10616 0.0
V29934 n1_20771_10799 n3_20771_10799 0.0
V29935 n1_20771_10832 n3_20771_10832 0.0
V29936 n1_20771_11015 n3_20771_11015 0.0
V29937 n1_20771_11048 n3_20771_11048 0.0
V29938 n1_20771_11231 n3_20771_11231 0.0
V29939 n1_20771_11264 n3_20771_11264 0.0
V29940 n1_20771_11447 n3_20771_11447 0.0
V29941 n1_20771_11480 n3_20771_11480 0.0
V29942 n1_20771_11663 n3_20771_11663 0.0
V29943 n1_20771_11696 n3_20771_11696 0.0
V29944 n1_20771_11879 n3_20771_11879 0.0
V29945 n1_20771_11912 n3_20771_11912 0.0
V29946 n1_20771_12095 n3_20771_12095 0.0
V29947 n1_20771_12128 n3_20771_12128 0.0
V29948 n1_20771_12311 n3_20771_12311 0.0
V29949 n1_20771_12344 n3_20771_12344 0.0
V29950 n1_20771_12527 n3_20771_12527 0.0
V29951 n1_20771_12560 n3_20771_12560 0.0
V29952 n1_20771_12743 n3_20771_12743 0.0
V29953 n1_20771_12776 n3_20771_12776 0.0
V29954 n1_20771_12959 n3_20771_12959 0.0
V29955 n1_20771_12992 n3_20771_12992 0.0
V29956 n1_20771_13175 n3_20771_13175 0.0
V29957 n1_20771_13208 n3_20771_13208 0.0
V29958 n1_20771_13391 n3_20771_13391 0.0
V29959 n1_20771_13424 n3_20771_13424 0.0
V29960 n1_20771_13607 n3_20771_13607 0.0
V29961 n1_20771_13640 n3_20771_13640 0.0
V29962 n1_20771_13823 n3_20771_13823 0.0
V29963 n1_20771_13856 n3_20771_13856 0.0
V29964 n1_20771_14039 n3_20771_14039 0.0
V29965 n1_20771_14072 n3_20771_14072 0.0
V29966 n1_20771_14255 n3_20771_14255 0.0
V29967 n1_20771_14288 n3_20771_14288 0.0
V29968 n1_20771_14471 n3_20771_14471 0.0
V29969 n1_20771_14504 n3_20771_14504 0.0
V29970 n1_20771_14687 n3_20771_14687 0.0
V29971 n1_20771_14720 n3_20771_14720 0.0
V29972 n1_20771_14903 n3_20771_14903 0.0
V29973 n1_20771_14936 n3_20771_14936 0.0
V29974 n1_20771_15092 n3_20771_15092 0.0
V29975 n1_20771_15119 n3_20771_15119 0.0
V29976 n1_20771_15152 n3_20771_15152 0.0
V29977 n1_20771_15308 n3_20771_15308 0.0
V29978 n1_20771_15335 n3_20771_15335 0.0
V29979 n1_20771_15368 n3_20771_15368 0.0
V29980 n1_20771_15551 n3_20771_15551 0.0
V29981 n1_20771_15584 n3_20771_15584 0.0
V29982 n1_20771_15767 n3_20771_15767 0.0
V29983 n1_20771_15800 n3_20771_15800 0.0
V29984 n1_20771_15983 n3_20771_15983 0.0
V29985 n1_20771_16016 n3_20771_16016 0.0
V29986 n1_20771_16199 n3_20771_16199 0.0
V29987 n1_20771_16415 n3_20771_16415 0.0
V29988 n1_20771_16448 n3_20771_16448 0.0
V29989 n1_20771_16631 n3_20771_16631 0.0
V29990 n1_20771_16664 n3_20771_16664 0.0
V29991 n1_20771_16798 n3_20771_16798 0.0
V29992 n1_20771_16847 n3_20771_16847 0.0
V29993 n1_20771_16880 n3_20771_16880 0.0
V29994 n1_20771_17063 n3_20771_17063 0.0
V29995 n1_20771_17096 n3_20771_17096 0.0
V29996 n1_20771_17279 n3_20771_17279 0.0
V29997 n1_20771_17312 n3_20771_17312 0.0
V29998 n1_20771_17495 n3_20771_17495 0.0
V29999 n1_20771_17528 n3_20771_17528 0.0
V30000 n1_20771_17711 n3_20771_17711 0.0
V30001 n1_20771_17744 n3_20771_17744 0.0
V30002 n1_20771_17927 n3_20771_17927 0.0
V30003 n1_20771_17960 n3_20771_17960 0.0
V30004 n1_20771_18143 n3_20771_18143 0.0
V30005 n1_20771_18176 n3_20771_18176 0.0
V30006 n1_20771_18359 n3_20771_18359 0.0
V30007 n1_20771_18392 n3_20771_18392 0.0
V30008 n1_20771_18527 n3_20771_18527 0.0
V30009 n1_20771_18575 n3_20771_18575 0.0
V30010 n1_20771_18608 n3_20771_18608 0.0
V30011 n1_20771_18791 n3_20771_18791 0.0
V30012 n1_20771_18824 n3_20771_18824 0.0
V30013 n1_20771_19007 n3_20771_19007 0.0
V30014 n1_20771_19040 n3_20771_19040 0.0
V30015 n1_20771_19223 n3_20771_19223 0.0
V30016 n1_20771_19256 n3_20771_19256 0.0
V30017 n1_20771_19439 n3_20771_19439 0.0
V30018 n1_20771_19472 n3_20771_19472 0.0
V30019 n1_20771_19655 n3_20771_19655 0.0
V30020 n1_20771_19688 n3_20771_19688 0.0
V30021 n1_20771_19871 n3_20771_19871 0.0
V30022 n1_20771_19904 n3_20771_19904 0.0
V30023 n1_20771_20087 n3_20771_20087 0.0
V30024 n1_20771_20120 n3_20771_20120 0.0
V30025 n1_20771_20303 n3_20771_20303 0.0
V30026 n1_20771_20336 n3_20771_20336 0.0
V30027 n1_20771_20519 n3_20771_20519 0.0
V30028 n1_20771_20552 n3_20771_20552 0.0
V30029 n1_20771_20687 n3_20771_20687 0.0
rr1b4 n3_2630_9471 _X_n3_2630_9471 2.500000e-01
v219 _X_n3_13880_20721 0 1.8
v15f _X_n2_2630_3846 0 0
rrd4 n2_19505_3846 _X_n2_19505_3846 2.500000e-01
v221 _X_n3_11630_20721 0 1.8
rr1b6 n3_4880_9471 _X_n3_4880_9471 2.500000e-01
rrd6 n2_18380_3846 _X_n2_18380_3846 2.500000e-01
v223 _X_n3_11630_18471 0 1.8
rr1b8 n3_7130_9471 _X_n3_7130_9471 2.500000e-01
rr1c0 n3_380_4971 _X_n3_380_4971 2.500000e-01
rrd8 n2_17255_3846 _X_n2_17255_3846 2.500000e-01
v225 _X_n3_11630_16221 0 1.8
v16b _X_n3_7130_20721 0 1.8
rre0 n2_17255_6096 _X_n2_17255_6096 2.500000e-01
rr1c2 n3_2630_4971 _X_n3_2630_4971 2.500000e-01
v227 _X_n3_11630_13971 0 1.8
v16d _X_n3_7130_18471 0 1.8
rre2 n2_16130_6096 _X_n2_16130_6096 2.500000e-01
rr1c4 n3_380_2721 _X_n3_380_2721 2.500000e-01
v229 _X_n3_11630_11721 0 1.8
v16f _X_n3_7130_16221 0 1.8
rre4 n2_15005_6096 _X_n2_15005_6096 2.500000e-01
rr1c6 n3_11630_471 _X_n3_11630_471 2.500000e-01
rre6 n2_20630_8346 _X_n2_20630_8346 2.500000e-01
rr1c8 n3_11630_2721 _X_n3_11630_2721 2.500000e-01
rr1d0 n3_13880_2721 _X_n3_13880_2721 2.500000e-01
rre8 n2_19505_8346 _X_n2_19505_8346 2.500000e-01
v17b _X_n3_2630_18471 0 1.8
rrf0 n2_15005_8346 _X_n2_15005_8346 2.500000e-01
rr1d2 n3_13880_4971 _X_n3_13880_4971 2.500000e-01
v17d _X_n3_380_16221 0 1.8
rrf2 n2_13880_8346 _X_n2_13880_8346 2.500000e-01
rr1d4 n3_16130_471 _X_n3_16130_471 2.500000e-01
v17f _X_n3_2630_16221 0 1.8
rrf4 n2_12755_8346 _X_n2_12755_8346 2.500000e-01
rraa n2_7130_10596 _X_n2_7130_10596 2.500000e-01
rr1d6 n3_16130_2721 _X_n3_16130_2721 2.500000e-01
rrf6 n2_20630_10596 _X_n2_20630_10596 2.500000e-01
rrac n2_8255_10596 _X_n2_8255_10596 2.500000e-01
rr1d8 n3_18380_471 _X_n3_18380_471 2.500000e-01
rr1e0 n3_20630_4971 _X_n3_20630_4971 2.500000e-01
rrf8 n2_19505_10596 _X_n2_19505_10596 2.500000e-01
rrae n2_9380_10596 _X_n2_9380_10596 2.500000e-01
v18b _X_n3_380_11721 0 1.8
rr1e2 n3_18380_4971 _X_n3_18380_4971 2.500000e-01
v18d _X_n3_2630_11721 0 1.8
rr1e4 n3_16130_4971 _X_n3_16130_4971 2.500000e-01
v18f _X_n3_4880_11721 0 1.8
rrba n2_12755_6096 _X_n2_12755_6096 2.500000e-01
rr1e6 n3_20630_7221 _X_n3_20630_7221 2.500000e-01
rrbc n2_12755_7221 _X_n2_12755_7221 2.500000e-01
rr1e8 n3_18380_7221 _X_n3_18380_7221 2.500000e-01
rr1f0 n3_18380_9471 _X_n3_18380_9471 2.500000e-01
rrbe n2_15005_471 _X_n2_15005_471 2.500000e-01
v20b _X_n3_20630_18471 0 1.8
v19b _X_n3_4880_471 0 1.8
rr1f2 n3_16130_9471 _X_n3_16130_9471 2.500000e-01
v20d _X_n3_20630_20721 0 1.8
v19d _X_n3_4880_2721 0 1.8
rr1f4 n3_13880_9471 _X_n3_13880_9471 2.500000e-01
rr1aa n3_9380_2721 _X_n3_9380_2721 2.500000e-01
v20f _X_n3_18380_20721 0 1.8
v19f _X_n3_4880_4971 0 1.8
rrca n2_17255_1596 _X_n2_17255_1596 2.500000e-01
rr1f6 n3_11630_9471 _X_n3_11630_9471 2.500000e-01
rr1ac n3_9380_4971 _X_n3_9380_4971 2.500000e-01
* layer: M5,GND net: 0
R30030 n0_241_1065 n0_429_1065 1.074286e+00
R30031 n0_429_1065 n0_1366_1065 5.354286e+00
R30032 n0_1366_1065 n0_1458_1065 5.257143e-01
R30033 n0_1458_1065 n0_1554_1065 5.485714e-01
R30034 n0_1554_1065 n0_1646_1065 5.257143e-01
R30035 n0_1646_1065 n0_3616_1065 1.125714e+01
R30036 n0_3616_1065 n0_3708_1065 5.257143e-01
R30037 n0_3708_1065 n0_3804_1065 5.485714e-01
R30038 n0_3804_1065 n0_3896_1065 5.257143e-01
R30039 n0_3896_1065 n0_5866_1065 1.125714e+01
R30040 n0_5866_1065 n0_5958_1065 5.257143e-01
R30041 n0_5958_1065 n0_6054_1065 5.485714e-01
R30042 n0_6054_1065 n0_6146_1065 5.257143e-01
R30043 n0_6146_1065 n0_8116_1065 1.125714e+01
R30044 n0_8116_1065 n0_8208_1065 5.257143e-01
R30045 n0_8208_1065 n0_8304_1065 5.485714e-01
R30046 n0_8304_1065 n0_8396_1065 5.257143e-01
R30047 n0_1366_417 n0_1458_417 5.257143e-01
R30048 n0_1458_417 n0_1505_417 2.685714e-01
R30049 n0_1505_417 n0_1554_417 2.800000e-01
R30050 n0_1554_417 n0_1646_417 5.257143e-01
R30051 n0_1646_417 n0_3616_417 1.125714e+01
R30052 n0_3616_417 n0_3708_417 5.257143e-01
R30053 n0_3708_417 n0_3755_417 2.685714e-01
R30054 n0_3755_417 n0_3804_417 2.800000e-01
R30055 n0_3804_417 n0_3896_417 5.257143e-01
R30056 n0_3896_417 n0_5866_417 1.125714e+01
R30057 n0_5866_417 n0_5958_417 5.257143e-01
R30058 n0_5958_417 n0_6005_417 2.685714e-01
R30059 n0_6005_417 n0_6054_417 2.800000e-01
R30060 n0_6054_417 n0_6146_417 5.257143e-01
R30061 n0_6146_417 n0_8116_417 1.125714e+01
R30062 n0_8116_417 n0_8208_417 5.257143e-01
R30063 n0_8208_417 n0_8255_417 2.685714e-01
R30064 n0_8255_417 n0_8304_417 2.800000e-01
R30065 n0_8304_417 n0_8396_417 5.257143e-01
R30066 n0_1366_450 n0_1458_450 5.257143e-01
R30067 n0_1458_450 n0_1505_450 2.685714e-01
R30068 n0_1505_450 n0_1554_450 2.800000e-01
R30069 n0_1554_450 n0_1646_450 5.257143e-01
R30070 n0_1646_450 n0_3616_450 1.125714e+01
R30071 n0_3616_450 n0_3708_450 5.257143e-01
R30072 n0_3708_450 n0_3755_450 2.685714e-01
R30073 n0_3755_450 n0_3804_450 2.800000e-01
R30074 n0_3804_450 n0_3896_450 5.257143e-01
R30075 n0_3896_450 n0_5866_450 1.125714e+01
R30076 n0_5866_450 n0_5958_450 5.257143e-01
R30077 n0_5958_450 n0_6005_450 2.685714e-01
R30078 n0_6005_450 n0_6054_450 2.800000e-01
R30079 n0_6054_450 n0_6146_450 5.257143e-01
R30080 n0_6146_450 n0_8116_450 1.125714e+01
R30081 n0_8116_450 n0_8208_450 5.257143e-01
R30082 n0_8208_450 n0_8255_450 2.685714e-01
R30083 n0_8255_450 n0_8304_450 2.800000e-01
R30084 n0_8304_450 n0_8396_450 5.257143e-01
R30085 n0_241_633 n0_429_633 1.074286e+00
R30086 n0_429_633 n0_1366_633 5.354286e+00
R30087 n0_1366_633 n0_1458_633 5.257143e-01
R30088 n0_1458_633 n0_1554_633 5.485714e-01
R30089 n0_1554_633 n0_1646_633 5.257143e-01
R30090 n0_1646_633 n0_3616_633 1.125714e+01
R30091 n0_3616_633 n0_3708_633 5.257143e-01
R30092 n0_3708_633 n0_3804_633 5.485714e-01
R30093 n0_3804_633 n0_3896_633 5.257143e-01
R30094 n0_3896_633 n0_5866_633 1.125714e+01
R30095 n0_5866_633 n0_5958_633 5.257143e-01
R30096 n0_5958_633 n0_6054_633 5.485714e-01
R30097 n0_6054_633 n0_6146_633 5.257143e-01
R30098 n0_6146_633 n0_8116_633 1.125714e+01
R30099 n0_8116_633 n0_8208_633 5.257143e-01
R30100 n0_8208_633 n0_8304_633 5.485714e-01
R30101 n0_8304_633 n0_8396_633 5.257143e-01
R30102 n0_241_666 n0_429_666 1.074286e+00
R30103 n0_429_666 n0_1366_666 5.354286e+00
R30104 n0_1366_666 n0_1458_666 5.257143e-01
R30105 n0_1458_666 n0_1554_666 5.485714e-01
R30106 n0_1554_666 n0_1646_666 5.257143e-01
R30107 n0_1646_666 n0_3616_666 1.125714e+01
R30108 n0_3616_666 n0_3708_666 5.257143e-01
R30109 n0_3708_666 n0_3804_666 5.485714e-01
R30110 n0_3804_666 n0_3896_666 5.257143e-01
R30111 n0_3896_666 n0_5866_666 1.125714e+01
R30112 n0_5866_666 n0_5958_666 5.257143e-01
R30113 n0_5958_666 n0_6054_666 5.485714e-01
R30114 n0_6054_666 n0_6146_666 5.257143e-01
R30115 n0_6146_666 n0_8116_666 1.125714e+01
R30116 n0_8116_666 n0_8208_666 5.257143e-01
R30117 n0_8208_666 n0_8304_666 5.485714e-01
R30118 n0_8304_666 n0_8396_666 5.257143e-01
R30119 n0_241_849 n0_429_849 1.074286e+00
R30120 n0_429_849 n0_1366_849 5.354286e+00
R30121 n0_1366_849 n0_1458_849 5.257143e-01
R30122 n0_1458_849 n0_1554_849 5.485714e-01
R30123 n0_1554_849 n0_1646_849 5.257143e-01
R30124 n0_1646_849 n0_3616_849 1.125714e+01
R30125 n0_3616_849 n0_3708_849 5.257143e-01
R30126 n0_3708_849 n0_3804_849 5.485714e-01
R30127 n0_3804_849 n0_3896_849 5.257143e-01
R30128 n0_3896_849 n0_5866_849 1.125714e+01
R30129 n0_5866_849 n0_5958_849 5.257143e-01
R30130 n0_5958_849 n0_6054_849 5.485714e-01
R30131 n0_6054_849 n0_6146_849 5.257143e-01
R30132 n0_6146_849 n0_8116_849 1.125714e+01
R30133 n0_8116_849 n0_8208_849 5.257143e-01
R30134 n0_8208_849 n0_8304_849 5.485714e-01
R30135 n0_8304_849 n0_8396_849 5.257143e-01
R30136 n0_241_882 n0_429_882 1.074286e+00
R30137 n0_429_882 n0_1366_882 5.354286e+00
R30138 n0_1366_882 n0_1458_882 5.257143e-01
R30139 n0_1458_882 n0_1554_882 5.485714e-01
R30140 n0_1554_882 n0_1646_882 5.257143e-01
R30141 n0_1646_882 n0_3616_882 1.125714e+01
R30142 n0_3616_882 n0_3708_882 5.257143e-01
R30143 n0_3708_882 n0_3804_882 5.485714e-01
R30144 n0_3804_882 n0_3896_882 5.257143e-01
R30145 n0_3896_882 n0_5866_882 1.125714e+01
R30146 n0_5866_882 n0_5958_882 5.257143e-01
R30147 n0_5958_882 n0_6054_882 5.485714e-01
R30148 n0_6054_882 n0_6146_882 5.257143e-01
R30149 n0_6146_882 n0_8116_882 1.125714e+01
R30150 n0_8116_882 n0_8208_882 5.257143e-01
R30151 n0_8208_882 n0_8304_882 5.485714e-01
R30152 n0_8304_882 n0_8396_882 5.257143e-01
R30153 n0_241_9273 n0_429_9273 1.074286e+00
R30154 n0_429_9273 n0_1366_9273 5.354286e+00
R30155 n0_1366_9273 n0_1554_9273 1.074286e+00
R30156 n0_1554_9273 n0_2491_9273 5.354286e+00
R30157 n0_2491_9273 n0_2679_9273 1.074286e+00
R30158 n0_2679_9273 n0_3616_9273 5.354286e+00
R30159 n0_3616_9273 n0_3804_9273 1.074286e+00
R30160 n0_3804_9273 n0_4741_9273 5.354286e+00
R30161 n0_4741_9273 n0_4929_9273 1.074286e+00
R30162 n0_4929_9273 n0_5866_9273 5.354286e+00
R30163 n0_5866_9273 n0_6054_9273 1.074286e+00
R30164 n0_6054_9273 n0_6991_9273 5.354286e+00
R30165 n0_6991_9273 n0_7179_9273 1.074286e+00
R30166 n0_7179_9273 n0_8116_9273 5.354286e+00
R30167 n0_8116_9273 n0_8304_9273 1.074286e+00
R30168 n0_8304_9273 n0_10366_9273 1.178286e+01
R30169 n0_10366_9273 n0_10458_9273 5.257143e-01
R30170 n0_10458_9273 n0_10554_9273 5.485714e-01
R30171 n0_10554_9273 n0_10646_9273 5.257143e-01
R30172 n0_10646_9273 n0_12616_9273 1.125714e+01
R30173 n0_12616_9273 n0_12804_9273 1.074286e+00
R30174 n0_12804_9273 n0_13741_9273 5.354286e+00
R30175 n0_13741_9273 n0_13929_9273 1.074286e+00
R30176 n0_13929_9273 n0_14866_9273 5.354286e+00
R30177 n0_14866_9273 n0_15054_9273 1.074286e+00
R30178 n0_15054_9273 n0_15991_9273 5.354286e+00
R30179 n0_15991_9273 n0_16179_9273 1.074286e+00
R30180 n0_16179_9273 n0_17116_9273 5.354286e+00
R30181 n0_17116_9273 n0_17304_9273 1.074286e+00
R30182 n0_17304_9273 n0_18241_9273 5.354286e+00
R30183 n0_18241_9273 n0_18429_9273 1.074286e+00
R30184 n0_18429_9273 n0_19366_9273 5.354286e+00
R30185 n0_19366_9273 n0_19554_9273 1.074286e+00
R30186 n0_241_9306 n0_429_9306 1.074286e+00
R30187 n0_429_9306 n0_1366_9306 5.354286e+00
R30188 n0_1366_9306 n0_1554_9306 1.074286e+00
R30189 n0_1554_9306 n0_2491_9306 5.354286e+00
R30190 n0_2491_9306 n0_2679_9306 1.074286e+00
R30191 n0_2679_9306 n0_3616_9306 5.354286e+00
R30192 n0_3616_9306 n0_3804_9306 1.074286e+00
R30193 n0_3804_9306 n0_4741_9306 5.354286e+00
R30194 n0_4741_9306 n0_4929_9306 1.074286e+00
R30195 n0_4929_9306 n0_5866_9306 5.354286e+00
R30196 n0_5866_9306 n0_6054_9306 1.074286e+00
R30197 n0_6054_9306 n0_6991_9306 5.354286e+00
R30198 n0_6991_9306 n0_7179_9306 1.074286e+00
R30199 n0_7179_9306 n0_8116_9306 5.354286e+00
R30200 n0_8116_9306 n0_8304_9306 1.074286e+00
R30201 n0_8304_9306 n0_10366_9306 1.178286e+01
R30202 n0_10366_9306 n0_10458_9306 5.257143e-01
R30203 n0_10458_9306 n0_10554_9306 5.485714e-01
R30204 n0_10554_9306 n0_10646_9306 5.257143e-01
R30205 n0_10646_9306 n0_12616_9306 1.125714e+01
R30206 n0_12616_9306 n0_12804_9306 1.074286e+00
R30207 n0_12804_9306 n0_13741_9306 5.354286e+00
R30208 n0_13741_9306 n0_13929_9306 1.074286e+00
R30209 n0_13929_9306 n0_14866_9306 5.354286e+00
R30210 n0_14866_9306 n0_15054_9306 1.074286e+00
R30211 n0_15054_9306 n0_15991_9306 5.354286e+00
R30212 n0_15991_9306 n0_16179_9306 1.074286e+00
R30213 n0_16179_9306 n0_17116_9306 5.354286e+00
R30214 n0_17116_9306 n0_17304_9306 1.074286e+00
R30215 n0_17304_9306 n0_18241_9306 5.354286e+00
R30216 n0_18241_9306 n0_18429_9306 1.074286e+00
R30217 n0_18429_9306 n0_19366_9306 5.354286e+00
R30218 n0_19366_9306 n0_19554_9306 1.074286e+00
R30219 n0_241_9489 n0_1366_9489 6.428571e+00
R30220 n0_1366_9489 n0_2491_9489 6.428571e+00
R30221 n0_2491_9489 n0_3616_9489 6.428571e+00
R30222 n0_3616_9489 n0_4741_9489 6.428571e+00
R30223 n0_4741_9489 n0_5866_9489 6.428571e+00
R30224 n0_5866_9489 n0_6991_9489 6.428571e+00
R30225 n0_6991_9489 n0_8116_9489 6.428571e+00
R30226 n0_8116_9489 n0_9241_9489 6.428571e+00
R30227 n0_9241_9489 n0_10366_9489 6.428571e+00
R30228 n0_10366_9489 n0_10458_9489 5.257143e-01
R30229 n0_10458_9489 n0_10505_9489 2.685714e-01
R30230 n0_10505_9489 n0_10554_9489 2.800000e-01
R30231 n0_10554_9489 n0_10646_9489 5.257143e-01
R30232 n0_10646_9489 n0_11491_9489 4.828571e+00
R30233 n0_11491_9489 n0_12616_9489 6.428571e+00
R30234 n0_12616_9489 n0_13741_9489 6.428571e+00
R30235 n0_13741_9489 n0_14866_9489 6.428571e+00
R30236 n0_14866_9489 n0_15991_9489 6.428571e+00
R30237 n0_15991_9489 n0_17116_9489 6.428571e+00
R30238 n0_17116_9489 n0_18241_9489 6.428571e+00
R30239 n0_18241_9489 n0_19366_9489 6.428571e+00
R30240 n0_241_9522 n0_1366_9522 6.428571e+00
R30241 n0_1366_9522 n0_2491_9522 6.428571e+00
R30242 n0_2491_9522 n0_3616_9522 6.428571e+00
R30243 n0_3616_9522 n0_4741_9522 6.428571e+00
R30244 n0_4741_9522 n0_5866_9522 6.428571e+00
R30245 n0_5866_9522 n0_6991_9522 6.428571e+00
R30246 n0_6991_9522 n0_8116_9522 6.428571e+00
R30247 n0_8116_9522 n0_9241_9522 6.428571e+00
R30248 n0_9241_9522 n0_10366_9522 6.428571e+00
R30249 n0_10366_9522 n0_10458_9522 5.257143e-01
R30250 n0_10458_9522 n0_10505_9522 2.685714e-01
R30251 n0_10505_9522 n0_10554_9522 2.800000e-01
R30252 n0_10554_9522 n0_10646_9522 5.257143e-01
R30253 n0_10646_9522 n0_11491_9522 4.828571e+00
R30254 n0_11491_9522 n0_12616_9522 6.428571e+00
R30255 n0_12616_9522 n0_13741_9522 6.428571e+00
R30256 n0_13741_9522 n0_14866_9522 6.428571e+00
R30257 n0_14866_9522 n0_15991_9522 6.428571e+00
R30258 n0_15991_9522 n0_17116_9522 6.428571e+00
R30259 n0_17116_9522 n0_18241_9522 6.428571e+00
R30260 n0_18241_9522 n0_19366_9522 6.428571e+00
R30261 n0_241_9705 n0_429_9705 1.074286e+00
R30262 n0_429_9705 n0_1366_9705 5.354286e+00
R30263 n0_1366_9705 n0_1554_9705 1.074286e+00
R30264 n0_1554_9705 n0_2491_9705 5.354286e+00
R30265 n0_2491_9705 n0_2679_9705 1.074286e+00
R30266 n0_2679_9705 n0_3616_9705 5.354286e+00
R30267 n0_3616_9705 n0_3804_9705 1.074286e+00
R30268 n0_3804_9705 n0_4741_9705 5.354286e+00
R30269 n0_4741_9705 n0_4929_9705 1.074286e+00
R30270 n0_4929_9705 n0_5866_9705 5.354286e+00
R30271 n0_5866_9705 n0_6054_9705 1.074286e+00
R30272 n0_6054_9705 n0_6991_9705 5.354286e+00
R30273 n0_6991_9705 n0_7179_9705 1.074286e+00
R30274 n0_7179_9705 n0_8116_9705 5.354286e+00
R30275 n0_8116_9705 n0_8304_9705 1.074286e+00
R30276 n0_8304_9705 n0_9241_9705 5.354286e+00
R30277 n0_9241_9705 n0_9429_9705 1.074286e+00
R30278 n0_9429_9705 n0_10366_9705 5.354286e+00
R30279 n0_10366_9705 n0_10458_9705 5.257143e-01
R30280 n0_10458_9705 n0_10554_9705 5.485714e-01
R30281 n0_10554_9705 n0_10646_9705 5.257143e-01
R30282 n0_10646_9705 n0_11491_9705 4.828571e+00
R30283 n0_11491_9705 n0_11679_9705 1.074286e+00
R30284 n0_11679_9705 n0_12616_9705 5.354286e+00
R30285 n0_12616_9705 n0_12804_9705 1.074286e+00
R30286 n0_12804_9705 n0_13741_9705 5.354286e+00
R30287 n0_13741_9705 n0_13929_9705 1.074286e+00
R30288 n0_13929_9705 n0_14866_9705 5.354286e+00
R30289 n0_14866_9705 n0_15054_9705 1.074286e+00
R30290 n0_15054_9705 n0_15991_9705 5.354286e+00
R30291 n0_15991_9705 n0_16179_9705 1.074286e+00
R30292 n0_16179_9705 n0_17116_9705 5.354286e+00
R30293 n0_17116_9705 n0_17304_9705 1.074286e+00
R30294 n0_17304_9705 n0_18241_9705 5.354286e+00
R30295 n0_18241_9705 n0_18429_9705 1.074286e+00
R30296 n0_18429_9705 n0_19366_9705 5.354286e+00
R30297 n0_19366_9705 n0_19554_9705 1.074286e+00
R30298 n0_241_9738 n0_429_9738 1.074286e+00
R30299 n0_429_9738 n0_1366_9738 5.354286e+00
R30300 n0_1366_9738 n0_1554_9738 1.074286e+00
R30301 n0_1554_9738 n0_2491_9738 5.354286e+00
R30302 n0_2491_9738 n0_2679_9738 1.074286e+00
R30303 n0_2679_9738 n0_3616_9738 5.354286e+00
R30304 n0_3616_9738 n0_3804_9738 1.074286e+00
R30305 n0_3804_9738 n0_4741_9738 5.354286e+00
R30306 n0_4741_9738 n0_4929_9738 1.074286e+00
R30307 n0_4929_9738 n0_5866_9738 5.354286e+00
R30308 n0_5866_9738 n0_6054_9738 1.074286e+00
R30309 n0_6054_9738 n0_6991_9738 5.354286e+00
R30310 n0_6991_9738 n0_7179_9738 1.074286e+00
R30311 n0_7179_9738 n0_8116_9738 5.354286e+00
R30312 n0_8116_9738 n0_8304_9738 1.074286e+00
R30313 n0_8304_9738 n0_9241_9738 5.354286e+00
R30314 n0_9241_9738 n0_9429_9738 1.074286e+00
R30315 n0_9429_9738 n0_10366_9738 5.354286e+00
R30316 n0_10366_9738 n0_10458_9738 5.257143e-01
R30317 n0_10458_9738 n0_10554_9738 5.485714e-01
R30318 n0_10554_9738 n0_10646_9738 5.257143e-01
R30319 n0_10646_9738 n0_11491_9738 4.828571e+00
R30320 n0_11491_9738 n0_11679_9738 1.074286e+00
R30321 n0_11679_9738 n0_12616_9738 5.354286e+00
R30322 n0_12616_9738 n0_12804_9738 1.074286e+00
R30323 n0_12804_9738 n0_13741_9738 5.354286e+00
R30324 n0_13741_9738 n0_13929_9738 1.074286e+00
R30325 n0_13929_9738 n0_14866_9738 5.354286e+00
R30326 n0_14866_9738 n0_15054_9738 1.074286e+00
R30327 n0_15054_9738 n0_15991_9738 5.354286e+00
R30328 n0_15991_9738 n0_16179_9738 1.074286e+00
R30329 n0_16179_9738 n0_17116_9738 5.354286e+00
R30330 n0_17116_9738 n0_17304_9738 1.074286e+00
R30331 n0_17304_9738 n0_18241_9738 5.354286e+00
R30332 n0_18241_9738 n0_18429_9738 1.074286e+00
R30333 n0_18429_9738 n0_19366_9738 5.354286e+00
R30334 n0_19366_9738 n0_19554_9738 1.074286e+00
R30335 n0_241_9921 n0_429_9921 1.074286e+00
R30336 n0_429_9921 n0_1366_9921 5.354286e+00
R30337 n0_1366_9921 n0_1554_9921 1.074286e+00
R30338 n0_1554_9921 n0_2491_9921 5.354286e+00
R30339 n0_2491_9921 n0_2679_9921 1.074286e+00
R30340 n0_2679_9921 n0_3616_9921 5.354286e+00
R30341 n0_3616_9921 n0_3804_9921 1.074286e+00
R30342 n0_3804_9921 n0_4741_9921 5.354286e+00
R30343 n0_4741_9921 n0_4929_9921 1.074286e+00
R30344 n0_4929_9921 n0_5866_9921 5.354286e+00
R30345 n0_5866_9921 n0_6054_9921 1.074286e+00
R30346 n0_6054_9921 n0_6991_9921 5.354286e+00
R30347 n0_6991_9921 n0_7179_9921 1.074286e+00
R30348 n0_7179_9921 n0_8116_9921 5.354286e+00
R30349 n0_8116_9921 n0_8304_9921 1.074286e+00
R30350 n0_8304_9921 n0_9241_9921 5.354286e+00
R30351 n0_9241_9921 n0_9429_9921 1.074286e+00
R30352 n0_9429_9921 n0_10366_9921 5.354286e+00
R30353 n0_10366_9921 n0_10458_9921 5.257143e-01
R30354 n0_10458_9921 n0_10554_9921 5.485714e-01
R30355 n0_10554_9921 n0_10646_9921 5.257143e-01
R30356 n0_10646_9921 n0_11491_9921 4.828571e+00
R30357 n0_11491_9921 n0_11679_9921 1.074286e+00
R30358 n0_11679_9921 n0_12616_9921 5.354286e+00
R30359 n0_12616_9921 n0_12804_9921 1.074286e+00
R30360 n0_12804_9921 n0_13741_9921 5.354286e+00
R30361 n0_13741_9921 n0_13929_9921 1.074286e+00
R30362 n0_13929_9921 n0_14866_9921 5.354286e+00
R30363 n0_14866_9921 n0_15054_9921 1.074286e+00
R30364 n0_15054_9921 n0_15991_9921 5.354286e+00
R30365 n0_15991_9921 n0_16179_9921 1.074286e+00
R30366 n0_16179_9921 n0_17116_9921 5.354286e+00
R30367 n0_17116_9921 n0_17304_9921 1.074286e+00
R30368 n0_17304_9921 n0_18241_9921 5.354286e+00
R30369 n0_18241_9921 n0_18429_9921 1.074286e+00
R30370 n0_18429_9921 n0_19366_9921 5.354286e+00
R30371 n0_19366_9921 n0_19554_9921 1.074286e+00
R30372 n0_241_9954 n0_429_9954 1.074286e+00
R30373 n0_429_9954 n0_1366_9954 5.354286e+00
R30374 n0_1366_9954 n0_1554_9954 1.074286e+00
R30375 n0_1554_9954 n0_2491_9954 5.354286e+00
R30376 n0_2491_9954 n0_2679_9954 1.074286e+00
R30377 n0_2679_9954 n0_3616_9954 5.354286e+00
R30378 n0_3616_9954 n0_3804_9954 1.074286e+00
R30379 n0_3804_9954 n0_4741_9954 5.354286e+00
R30380 n0_4741_9954 n0_4929_9954 1.074286e+00
R30381 n0_4929_9954 n0_5866_9954 5.354286e+00
R30382 n0_5866_9954 n0_6054_9954 1.074286e+00
R30383 n0_6054_9954 n0_6991_9954 5.354286e+00
R30384 n0_6991_9954 n0_7179_9954 1.074286e+00
R30385 n0_7179_9954 n0_8116_9954 5.354286e+00
R30386 n0_8116_9954 n0_8304_9954 1.074286e+00
R30387 n0_8304_9954 n0_9241_9954 5.354286e+00
R30388 n0_9241_9954 n0_9429_9954 1.074286e+00
R30389 n0_9429_9954 n0_10366_9954 5.354286e+00
R30390 n0_10366_9954 n0_10458_9954 5.257143e-01
R30391 n0_10458_9954 n0_10554_9954 5.485714e-01
R30392 n0_10554_9954 n0_10646_9954 5.257143e-01
R30393 n0_10646_9954 n0_11491_9954 4.828571e+00
R30394 n0_11491_9954 n0_11679_9954 1.074286e+00
R30395 n0_11679_9954 n0_12616_9954 5.354286e+00
R30396 n0_12616_9954 n0_12804_9954 1.074286e+00
R30397 n0_12804_9954 n0_13741_9954 5.354286e+00
R30398 n0_13741_9954 n0_13929_9954 1.074286e+00
R30399 n0_13929_9954 n0_14866_9954 5.354286e+00
R30400 n0_14866_9954 n0_15054_9954 1.074286e+00
R30401 n0_15054_9954 n0_15991_9954 5.354286e+00
R30402 n0_15991_9954 n0_16179_9954 1.074286e+00
R30403 n0_16179_9954 n0_17116_9954 5.354286e+00
R30404 n0_17116_9954 n0_17304_9954 1.074286e+00
R30405 n0_17304_9954 n0_18241_9954 5.354286e+00
R30406 n0_18241_9954 n0_18429_9954 1.074286e+00
R30407 n0_18429_9954 n0_19366_9954 5.354286e+00
R30408 n0_19366_9954 n0_19554_9954 1.074286e+00
R30409 n0_241_10137 n0_429_10137 1.074286e+00
R30410 n0_429_10137 n0_1366_10137 5.354286e+00
R30411 n0_1366_10137 n0_1554_10137 1.074286e+00
R30412 n0_1554_10137 n0_2491_10137 5.354286e+00
R30413 n0_2491_10137 n0_2679_10137 1.074286e+00
R30414 n0_2679_10137 n0_3616_10137 5.354286e+00
R30415 n0_3616_10137 n0_3804_10137 1.074286e+00
R30416 n0_3804_10137 n0_4741_10137 5.354286e+00
R30417 n0_4741_10137 n0_4929_10137 1.074286e+00
R30418 n0_4929_10137 n0_5866_10137 5.354286e+00
R30419 n0_5866_10137 n0_6054_10137 1.074286e+00
R30420 n0_6054_10137 n0_6991_10137 5.354286e+00
R30421 n0_6991_10137 n0_7179_10137 1.074286e+00
R30422 n0_7179_10137 n0_8116_10137 5.354286e+00
R30423 n0_8116_10137 n0_8304_10137 1.074286e+00
R30424 n0_8304_10137 n0_9241_10137 5.354286e+00
R30425 n0_9241_10137 n0_9429_10137 1.074286e+00
R30426 n0_9429_10137 n0_10366_10137 5.354286e+00
R30427 n0_10366_10137 n0_10458_10137 5.257143e-01
R30428 n0_10458_10137 n0_10554_10137 5.485714e-01
R30429 n0_10554_10137 n0_10646_10137 5.257143e-01
R30430 n0_10646_10137 n0_11491_10137 4.828571e+00
R30431 n0_11491_10137 n0_11679_10137 1.074286e+00
R30432 n0_11679_10137 n0_12616_10137 5.354286e+00
R30433 n0_12616_10137 n0_12804_10137 1.074286e+00
R30434 n0_12804_10137 n0_13741_10137 5.354286e+00
R30435 n0_13741_10137 n0_13929_10137 1.074286e+00
R30436 n0_13929_10137 n0_14866_10137 5.354286e+00
R30437 n0_14866_10137 n0_15054_10137 1.074286e+00
R30438 n0_15054_10137 n0_15991_10137 5.354286e+00
R30439 n0_15991_10137 n0_16179_10137 1.074286e+00
R30440 n0_16179_10137 n0_17116_10137 5.354286e+00
R30441 n0_17116_10137 n0_17304_10137 1.074286e+00
R30442 n0_17304_10137 n0_18241_10137 5.354286e+00
R30443 n0_18241_10137 n0_18429_10137 1.074286e+00
R30444 n0_18429_10137 n0_19366_10137 5.354286e+00
R30445 n0_19366_10137 n0_19554_10137 1.074286e+00
R30446 n0_241_10170 n0_429_10170 1.074286e+00
R30447 n0_429_10170 n0_1366_10170 5.354286e+00
R30448 n0_1366_10170 n0_1554_10170 1.074286e+00
R30449 n0_1554_10170 n0_2491_10170 5.354286e+00
R30450 n0_2491_10170 n0_2679_10170 1.074286e+00
R30451 n0_2679_10170 n0_3616_10170 5.354286e+00
R30452 n0_3616_10170 n0_3804_10170 1.074286e+00
R30453 n0_3804_10170 n0_4741_10170 5.354286e+00
R30454 n0_4741_10170 n0_4929_10170 1.074286e+00
R30455 n0_4929_10170 n0_5866_10170 5.354286e+00
R30456 n0_5866_10170 n0_6054_10170 1.074286e+00
R30457 n0_6054_10170 n0_6991_10170 5.354286e+00
R30458 n0_6991_10170 n0_7179_10170 1.074286e+00
R30459 n0_7179_10170 n0_8116_10170 5.354286e+00
R30460 n0_8116_10170 n0_8304_10170 1.074286e+00
R30461 n0_8304_10170 n0_9241_10170 5.354286e+00
R30462 n0_9241_10170 n0_9429_10170 1.074286e+00
R30463 n0_9429_10170 n0_10366_10170 5.354286e+00
R30464 n0_10366_10170 n0_10458_10170 5.257143e-01
R30465 n0_10458_10170 n0_10554_10170 5.485714e-01
R30466 n0_10554_10170 n0_10646_10170 5.257143e-01
R30467 n0_10646_10170 n0_11491_10170 4.828571e+00
R30468 n0_11491_10170 n0_11679_10170 1.074286e+00
R30469 n0_11679_10170 n0_12616_10170 5.354286e+00
R30470 n0_12616_10170 n0_12804_10170 1.074286e+00
R30471 n0_12804_10170 n0_13741_10170 5.354286e+00
R30472 n0_13741_10170 n0_13929_10170 1.074286e+00
R30473 n0_13929_10170 n0_14866_10170 5.354286e+00
R30474 n0_14866_10170 n0_15054_10170 1.074286e+00
R30475 n0_15054_10170 n0_15991_10170 5.354286e+00
R30476 n0_15991_10170 n0_16179_10170 1.074286e+00
R30477 n0_16179_10170 n0_17116_10170 5.354286e+00
R30478 n0_17116_10170 n0_17304_10170 1.074286e+00
R30479 n0_17304_10170 n0_18241_10170 5.354286e+00
R30480 n0_18241_10170 n0_18429_10170 1.074286e+00
R30481 n0_18429_10170 n0_19366_10170 5.354286e+00
R30482 n0_19366_10170 n0_19554_10170 1.074286e+00
R30483 n0_241_10353 n0_429_10353 1.074286e+00
R30484 n0_429_10353 n0_1366_10353 5.354286e+00
R30485 n0_1366_10353 n0_1554_10353 1.074286e+00
R30486 n0_1554_10353 n0_2491_10353 5.354286e+00
R30487 n0_2491_10353 n0_2679_10353 1.074286e+00
R30488 n0_2679_10353 n0_3616_10353 5.354286e+00
R30489 n0_3616_10353 n0_3804_10353 1.074286e+00
R30490 n0_3804_10353 n0_4741_10353 5.354286e+00
R30491 n0_4741_10353 n0_4929_10353 1.074286e+00
R30492 n0_4929_10353 n0_5866_10353 5.354286e+00
R30493 n0_5866_10353 n0_6054_10353 1.074286e+00
R30494 n0_6054_10353 n0_6991_10353 5.354286e+00
R30495 n0_6991_10353 n0_7179_10353 1.074286e+00
R30496 n0_7179_10353 n0_8116_10353 5.354286e+00
R30497 n0_8116_10353 n0_8304_10353 1.074286e+00
R30498 n0_8304_10353 n0_9241_10353 5.354286e+00
R30499 n0_9241_10353 n0_9429_10353 1.074286e+00
R30500 n0_9429_10353 n0_10366_10353 5.354286e+00
R30501 n0_10366_10353 n0_10458_10353 5.257143e-01
R30502 n0_10458_10353 n0_10554_10353 5.485714e-01
R30503 n0_10554_10353 n0_10646_10353 5.257143e-01
R30504 n0_10646_10353 n0_11491_10353 4.828571e+00
R30505 n0_11491_10353 n0_11679_10353 1.074286e+00
R30506 n0_11679_10353 n0_12616_10353 5.354286e+00
R30507 n0_12616_10353 n0_12804_10353 1.074286e+00
R30508 n0_12804_10353 n0_13741_10353 5.354286e+00
R30509 n0_13741_10353 n0_13929_10353 1.074286e+00
R30510 n0_13929_10353 n0_14866_10353 5.354286e+00
R30511 n0_14866_10353 n0_15054_10353 1.074286e+00
R30512 n0_15054_10353 n0_15991_10353 5.354286e+00
R30513 n0_15991_10353 n0_16179_10353 1.074286e+00
R30514 n0_16179_10353 n0_17116_10353 5.354286e+00
R30515 n0_17116_10353 n0_17304_10353 1.074286e+00
R30516 n0_17304_10353 n0_18241_10353 5.354286e+00
R30517 n0_18241_10353 n0_18429_10353 1.074286e+00
R30518 n0_18429_10353 n0_19366_10353 5.354286e+00
R30519 n0_19366_10353 n0_19554_10353 1.074286e+00
R30520 n0_241_10386 n0_429_10386 1.074286e+00
R30521 n0_429_10386 n0_1366_10386 5.354286e+00
R30522 n0_1366_10386 n0_1554_10386 1.074286e+00
R30523 n0_1554_10386 n0_2491_10386 5.354286e+00
R30524 n0_2491_10386 n0_2679_10386 1.074286e+00
R30525 n0_2679_10386 n0_3616_10386 5.354286e+00
R30526 n0_3616_10386 n0_3804_10386 1.074286e+00
R30527 n0_3804_10386 n0_4741_10386 5.354286e+00
R30528 n0_4741_10386 n0_4929_10386 1.074286e+00
R30529 n0_4929_10386 n0_5866_10386 5.354286e+00
R30530 n0_5866_10386 n0_6054_10386 1.074286e+00
R30531 n0_6054_10386 n0_6991_10386 5.354286e+00
R30532 n0_6991_10386 n0_7179_10386 1.074286e+00
R30533 n0_7179_10386 n0_8116_10386 5.354286e+00
R30534 n0_8116_10386 n0_8304_10386 1.074286e+00
R30535 n0_8304_10386 n0_9241_10386 5.354286e+00
R30536 n0_9241_10386 n0_9429_10386 1.074286e+00
R30537 n0_9429_10386 n0_10366_10386 5.354286e+00
R30538 n0_10366_10386 n0_10458_10386 5.257143e-01
R30539 n0_10458_10386 n0_10554_10386 5.485714e-01
R30540 n0_10554_10386 n0_10646_10386 5.257143e-01
R30541 n0_10646_10386 n0_11491_10386 4.828571e+00
R30542 n0_11491_10386 n0_11679_10386 1.074286e+00
R30543 n0_11679_10386 n0_12616_10386 5.354286e+00
R30544 n0_12616_10386 n0_12804_10386 1.074286e+00
R30545 n0_12804_10386 n0_13741_10386 5.354286e+00
R30546 n0_13741_10386 n0_13929_10386 1.074286e+00
R30547 n0_13929_10386 n0_14866_10386 5.354286e+00
R30548 n0_14866_10386 n0_15054_10386 1.074286e+00
R30549 n0_15054_10386 n0_15991_10386 5.354286e+00
R30550 n0_15991_10386 n0_16179_10386 1.074286e+00
R30551 n0_16179_10386 n0_17116_10386 5.354286e+00
R30552 n0_17116_10386 n0_17304_10386 1.074286e+00
R30553 n0_17304_10386 n0_18241_10386 5.354286e+00
R30554 n0_18241_10386 n0_18429_10386 1.074286e+00
R30555 n0_18429_10386 n0_19366_10386 5.354286e+00
R30556 n0_19366_10386 n0_19554_10386 1.074286e+00
R30557 n0_241_10569 n0_380_10569 7.942857e-01
R30558 n0_380_10569 n0_429_10569 2.800000e-01
R30559 n0_429_10569 n0_1366_10569 5.354286e+00
R30560 n0_1366_10569 n0_1505_10569 7.942857e-01
R30561 n0_1505_10569 n0_1554_10569 2.800000e-01
R30562 n0_1554_10569 n0_2491_10569 5.354286e+00
R30563 n0_2491_10569 n0_2630_10569 7.942857e-01
R30564 n0_2630_10569 n0_2679_10569 2.800000e-01
R30565 n0_2679_10569 n0_3616_10569 5.354286e+00
R30566 n0_3616_10569 n0_3755_10569 7.942857e-01
R30567 n0_3755_10569 n0_3804_10569 2.800000e-01
R30568 n0_3804_10569 n0_4741_10569 5.354286e+00
R30569 n0_4741_10569 n0_4880_10569 7.942857e-01
R30570 n0_4880_10569 n0_4929_10569 2.800000e-01
R30571 n0_4929_10569 n0_5866_10569 5.354286e+00
R30572 n0_5866_10569 n0_6005_10569 7.942857e-01
R30573 n0_6005_10569 n0_6054_10569 2.800000e-01
R30574 n0_6054_10569 n0_6991_10569 5.354286e+00
R30575 n0_6991_10569 n0_7130_10569 7.942857e-01
R30576 n0_7130_10569 n0_7179_10569 2.800000e-01
R30577 n0_7179_10569 n0_8116_10569 5.354286e+00
R30578 n0_8116_10569 n0_8255_10569 7.942857e-01
R30579 n0_8255_10569 n0_8304_10569 2.800000e-01
R30580 n0_8304_10569 n0_9241_10569 5.354286e+00
R30581 n0_9241_10569 n0_9380_10569 7.942857e-01
R30582 n0_9380_10569 n0_9429_10569 2.800000e-01
R30583 n0_9429_10569 n0_10366_10569 5.354286e+00
R30584 n0_10366_10569 n0_10458_10569 5.257143e-01
R30585 n0_10458_10569 n0_10505_10569 2.685714e-01
R30586 n0_10505_10569 n0_10554_10569 2.800000e-01
R30587 n0_10554_10569 n0_10646_10569 5.257143e-01
R30588 n0_10646_10569 n0_11491_10569 4.828571e+00
R30589 n0_11491_10569 n0_11630_10569 7.942857e-01
R30590 n0_11630_10569 n0_11679_10569 2.800000e-01
R30591 n0_11679_10569 n0_12616_10569 5.354286e+00
R30592 n0_12616_10569 n0_12755_10569 7.942857e-01
R30593 n0_12755_10569 n0_12804_10569 2.800000e-01
R30594 n0_12804_10569 n0_13741_10569 5.354286e+00
R30595 n0_13741_10569 n0_13880_10569 7.942857e-01
R30596 n0_13880_10569 n0_13929_10569 2.800000e-01
R30597 n0_13929_10569 n0_14866_10569 5.354286e+00
R30598 n0_14866_10569 n0_15005_10569 7.942857e-01
R30599 n0_15005_10569 n0_15054_10569 2.800000e-01
R30600 n0_15054_10569 n0_15991_10569 5.354286e+00
R30601 n0_15991_10569 n0_16130_10569 7.942857e-01
R30602 n0_16130_10569 n0_16179_10569 2.800000e-01
R30603 n0_16179_10569 n0_17116_10569 5.354286e+00
R30604 n0_17116_10569 n0_17255_10569 7.942857e-01
R30605 n0_17255_10569 n0_17304_10569 2.800000e-01
R30606 n0_17304_10569 n0_18241_10569 5.354286e+00
R30607 n0_18241_10569 n0_18380_10569 7.942857e-01
R30608 n0_18380_10569 n0_18429_10569 2.800000e-01
R30609 n0_18429_10569 n0_19366_10569 5.354286e+00
R30610 n0_19366_10569 n0_19505_10569 7.942857e-01
R30611 n0_19505_10569 n0_19554_10569 2.800000e-01
R30612 n0_380_10602 n0_429_10602 2.800000e-01
R30613 n0_429_10602 n0_1505_10602 6.148571e+00
R30614 n0_1505_10602 n0_1554_10602 2.800000e-01
R30615 n0_1554_10602 n0_2630_10602 6.148571e+00
R30616 n0_2630_10602 n0_2679_10602 2.800000e-01
R30617 n0_2679_10602 n0_3755_10602 6.148571e+00
R30618 n0_3755_10602 n0_3804_10602 2.800000e-01
R30619 n0_3804_10602 n0_4880_10602 6.148571e+00
R30620 n0_4880_10602 n0_4929_10602 2.800000e-01
R30621 n0_4929_10602 n0_6005_10602 6.148571e+00
R30622 n0_6005_10602 n0_6054_10602 2.800000e-01
R30623 n0_6054_10602 n0_7130_10602 6.148571e+00
R30624 n0_7130_10602 n0_7179_10602 2.800000e-01
R30625 n0_7179_10602 n0_8255_10602 6.148571e+00
R30626 n0_8255_10602 n0_8304_10602 2.800000e-01
R30627 n0_8304_10602 n0_9380_10602 6.148571e+00
R30628 n0_9380_10602 n0_9429_10602 2.800000e-01
R30629 n0_9429_10602 n0_10458_10602 5.880000e+00
R30630 n0_10458_10602 n0_10505_10602 2.685714e-01
R30631 n0_10505_10602 n0_10554_10602 2.800000e-01
R30632 n0_10554_10602 n0_11630_10602 6.148571e+00
R30633 n0_11630_10602 n0_11679_10602 2.800000e-01
R30634 n0_11679_10602 n0_12755_10602 6.148571e+00
R30635 n0_12755_10602 n0_12804_10602 2.800000e-01
R30636 n0_12804_10602 n0_13880_10602 6.148571e+00
R30637 n0_13880_10602 n0_13929_10602 2.800000e-01
R30638 n0_13929_10602 n0_15005_10602 6.148571e+00
R30639 n0_15005_10602 n0_15054_10602 2.800000e-01
R30640 n0_15054_10602 n0_16130_10602 6.148571e+00
R30641 n0_16130_10602 n0_16179_10602 2.800000e-01
R30642 n0_16179_10602 n0_17255_10602 6.148571e+00
R30643 n0_17255_10602 n0_17304_10602 2.800000e-01
R30644 n0_17304_10602 n0_18380_10602 6.148571e+00
R30645 n0_18380_10602 n0_18429_10602 2.800000e-01
R30646 n0_18429_10602 n0_19505_10602 6.148571e+00
R30647 n0_19505_10602 n0_19554_10602 2.800000e-01
R30648 n0_241_10785 n0_429_10785 1.074286e+00
R30649 n0_429_10785 n0_1366_10785 5.354286e+00
R30650 n0_1366_10785 n0_1554_10785 1.074286e+00
R30651 n0_1554_10785 n0_2491_10785 5.354286e+00
R30652 n0_2491_10785 n0_2679_10785 1.074286e+00
R30653 n0_2679_10785 n0_3616_10785 5.354286e+00
R30654 n0_3616_10785 n0_3804_10785 1.074286e+00
R30655 n0_3804_10785 n0_4741_10785 5.354286e+00
R30656 n0_4741_10785 n0_4929_10785 1.074286e+00
R30657 n0_4929_10785 n0_5866_10785 5.354286e+00
R30658 n0_5866_10785 n0_6054_10785 1.074286e+00
R30659 n0_6054_10785 n0_6991_10785 5.354286e+00
R30660 n0_6991_10785 n0_7179_10785 1.074286e+00
R30661 n0_7179_10785 n0_8116_10785 5.354286e+00
R30662 n0_8116_10785 n0_8304_10785 1.074286e+00
R30663 n0_8304_10785 n0_9241_10785 5.354286e+00
R30664 n0_9241_10785 n0_9429_10785 1.074286e+00
R30665 n0_9429_10785 n0_10366_10785 5.354286e+00
R30666 n0_10366_10785 n0_10458_10785 5.257143e-01
R30667 n0_10458_10785 n0_10554_10785 5.485714e-01
R30668 n0_10554_10785 n0_10646_10785 5.257143e-01
R30669 n0_10646_10785 n0_11491_10785 4.828571e+00
R30670 n0_11491_10785 n0_11679_10785 1.074286e+00
R30671 n0_11679_10785 n0_12616_10785 5.354286e+00
R30672 n0_12616_10785 n0_12804_10785 1.074286e+00
R30673 n0_12804_10785 n0_13741_10785 5.354286e+00
R30674 n0_13741_10785 n0_13929_10785 1.074286e+00
R30675 n0_13929_10785 n0_14866_10785 5.354286e+00
R30676 n0_14866_10785 n0_15054_10785 1.074286e+00
R30677 n0_15054_10785 n0_15991_10785 5.354286e+00
R30678 n0_15991_10785 n0_16179_10785 1.074286e+00
R30679 n0_16179_10785 n0_17116_10785 5.354286e+00
R30680 n0_17116_10785 n0_17304_10785 1.074286e+00
R30681 n0_17304_10785 n0_18241_10785 5.354286e+00
R30682 n0_18241_10785 n0_18429_10785 1.074286e+00
R30683 n0_18429_10785 n0_19366_10785 5.354286e+00
R30684 n0_19366_10785 n0_19554_10785 1.074286e+00
R30685 n0_241_10818 n0_429_10818 1.074286e+00
R30686 n0_429_10818 n0_1366_10818 5.354286e+00
R30687 n0_1366_10818 n0_1554_10818 1.074286e+00
R30688 n0_1554_10818 n0_2491_10818 5.354286e+00
R30689 n0_2491_10818 n0_2679_10818 1.074286e+00
R30690 n0_2679_10818 n0_3616_10818 5.354286e+00
R30691 n0_3616_10818 n0_3804_10818 1.074286e+00
R30692 n0_3804_10818 n0_4741_10818 5.354286e+00
R30693 n0_4741_10818 n0_4929_10818 1.074286e+00
R30694 n0_4929_10818 n0_5866_10818 5.354286e+00
R30695 n0_5866_10818 n0_6054_10818 1.074286e+00
R30696 n0_6054_10818 n0_6991_10818 5.354286e+00
R30697 n0_6991_10818 n0_7179_10818 1.074286e+00
R30698 n0_7179_10818 n0_8116_10818 5.354286e+00
R30699 n0_8116_10818 n0_8304_10818 1.074286e+00
R30700 n0_8304_10818 n0_9241_10818 5.354286e+00
R30701 n0_9241_10818 n0_9429_10818 1.074286e+00
R30702 n0_9429_10818 n0_10366_10818 5.354286e+00
R30703 n0_10366_10818 n0_10458_10818 5.257143e-01
R30704 n0_10458_10818 n0_10554_10818 5.485714e-01
R30705 n0_10554_10818 n0_10646_10818 5.257143e-01
R30706 n0_10646_10818 n0_11491_10818 4.828571e+00
R30707 n0_11491_10818 n0_11679_10818 1.074286e+00
R30708 n0_11679_10818 n0_12616_10818 5.354286e+00
R30709 n0_12616_10818 n0_12804_10818 1.074286e+00
R30710 n0_12804_10818 n0_13741_10818 5.354286e+00
R30711 n0_13741_10818 n0_13929_10818 1.074286e+00
R30712 n0_13929_10818 n0_14866_10818 5.354286e+00
R30713 n0_14866_10818 n0_15054_10818 1.074286e+00
R30714 n0_15054_10818 n0_15991_10818 5.354286e+00
R30715 n0_15991_10818 n0_16179_10818 1.074286e+00
R30716 n0_16179_10818 n0_17116_10818 5.354286e+00
R30717 n0_17116_10818 n0_17304_10818 1.074286e+00
R30718 n0_17304_10818 n0_18241_10818 5.354286e+00
R30719 n0_18241_10818 n0_18429_10818 1.074286e+00
R30720 n0_18429_10818 n0_19366_10818 5.354286e+00
R30721 n0_19366_10818 n0_19554_10818 1.074286e+00
R30722 n0_241_11001 n0_429_11001 1.074286e+00
R30723 n0_429_11001 n0_1366_11001 5.354286e+00
R30724 n0_1366_11001 n0_1554_11001 1.074286e+00
R30725 n0_1554_11001 n0_2491_11001 5.354286e+00
R30726 n0_2491_11001 n0_2679_11001 1.074286e+00
R30727 n0_2679_11001 n0_3616_11001 5.354286e+00
R30728 n0_3616_11001 n0_3804_11001 1.074286e+00
R30729 n0_3804_11001 n0_4741_11001 5.354286e+00
R30730 n0_4741_11001 n0_4929_11001 1.074286e+00
R30731 n0_4929_11001 n0_5866_11001 5.354286e+00
R30732 n0_5866_11001 n0_6054_11001 1.074286e+00
R30733 n0_6054_11001 n0_6991_11001 5.354286e+00
R30734 n0_6991_11001 n0_7179_11001 1.074286e+00
R30735 n0_7179_11001 n0_8116_11001 5.354286e+00
R30736 n0_8116_11001 n0_8304_11001 1.074286e+00
R30737 n0_8304_11001 n0_9241_11001 5.354286e+00
R30738 n0_9241_11001 n0_9429_11001 1.074286e+00
R30739 n0_9429_11001 n0_10366_11001 5.354286e+00
R30740 n0_10366_11001 n0_10458_11001 5.257143e-01
R30741 n0_10458_11001 n0_10554_11001 5.485714e-01
R30742 n0_10554_11001 n0_10646_11001 5.257143e-01
R30743 n0_10646_11001 n0_11491_11001 4.828571e+00
R30744 n0_11491_11001 n0_11679_11001 1.074286e+00
R30745 n0_11679_11001 n0_12616_11001 5.354286e+00
R30746 n0_12616_11001 n0_12804_11001 1.074286e+00
R30747 n0_12804_11001 n0_13741_11001 5.354286e+00
R30748 n0_13741_11001 n0_13929_11001 1.074286e+00
R30749 n0_13929_11001 n0_14866_11001 5.354286e+00
R30750 n0_14866_11001 n0_15054_11001 1.074286e+00
R30751 n0_15054_11001 n0_15991_11001 5.354286e+00
R30752 n0_15991_11001 n0_16179_11001 1.074286e+00
R30753 n0_16179_11001 n0_17116_11001 5.354286e+00
R30754 n0_17116_11001 n0_17304_11001 1.074286e+00
R30755 n0_17304_11001 n0_18241_11001 5.354286e+00
R30756 n0_18241_11001 n0_18429_11001 1.074286e+00
R30757 n0_18429_11001 n0_19366_11001 5.354286e+00
R30758 n0_19366_11001 n0_19554_11001 1.074286e+00
R30759 n0_241_11034 n0_429_11034 1.074286e+00
R30760 n0_429_11034 n0_1366_11034 5.354286e+00
R30761 n0_1366_11034 n0_1554_11034 1.074286e+00
R30762 n0_1554_11034 n0_2491_11034 5.354286e+00
R30763 n0_2491_11034 n0_2679_11034 1.074286e+00
R30764 n0_2679_11034 n0_3616_11034 5.354286e+00
R30765 n0_3616_11034 n0_3804_11034 1.074286e+00
R30766 n0_3804_11034 n0_4741_11034 5.354286e+00
R30767 n0_4741_11034 n0_4929_11034 1.074286e+00
R30768 n0_4929_11034 n0_5866_11034 5.354286e+00
R30769 n0_5866_11034 n0_6054_11034 1.074286e+00
R30770 n0_6054_11034 n0_6991_11034 5.354286e+00
R30771 n0_6991_11034 n0_7179_11034 1.074286e+00
R30772 n0_7179_11034 n0_8116_11034 5.354286e+00
R30773 n0_8116_11034 n0_8304_11034 1.074286e+00
R30774 n0_8304_11034 n0_9241_11034 5.354286e+00
R30775 n0_9241_11034 n0_9429_11034 1.074286e+00
R30776 n0_9429_11034 n0_10366_11034 5.354286e+00
R30777 n0_10366_11034 n0_10458_11034 5.257143e-01
R30778 n0_10458_11034 n0_10554_11034 5.485714e-01
R30779 n0_10554_11034 n0_10646_11034 5.257143e-01
R30780 n0_10646_11034 n0_11491_11034 4.828571e+00
R30781 n0_11491_11034 n0_11679_11034 1.074286e+00
R30782 n0_11679_11034 n0_12616_11034 5.354286e+00
R30783 n0_12616_11034 n0_12804_11034 1.074286e+00
R30784 n0_12804_11034 n0_13741_11034 5.354286e+00
R30785 n0_13741_11034 n0_13929_11034 1.074286e+00
R30786 n0_13929_11034 n0_14866_11034 5.354286e+00
R30787 n0_14866_11034 n0_15054_11034 1.074286e+00
R30788 n0_15054_11034 n0_15991_11034 5.354286e+00
R30789 n0_15991_11034 n0_16179_11034 1.074286e+00
R30790 n0_16179_11034 n0_17116_11034 5.354286e+00
R30791 n0_17116_11034 n0_17304_11034 1.074286e+00
R30792 n0_17304_11034 n0_18241_11034 5.354286e+00
R30793 n0_18241_11034 n0_18429_11034 1.074286e+00
R30794 n0_18429_11034 n0_19366_11034 5.354286e+00
R30795 n0_19366_11034 n0_19554_11034 1.074286e+00
R30796 n0_241_11217 n0_429_11217 1.074286e+00
R30797 n0_429_11217 n0_1366_11217 5.354286e+00
R30798 n0_1366_11217 n0_1554_11217 1.074286e+00
R30799 n0_1554_11217 n0_2491_11217 5.354286e+00
R30800 n0_2491_11217 n0_2679_11217 1.074286e+00
R30801 n0_2679_11217 n0_3616_11217 5.354286e+00
R30802 n0_3616_11217 n0_3804_11217 1.074286e+00
R30803 n0_3804_11217 n0_4741_11217 5.354286e+00
R30804 n0_4741_11217 n0_4929_11217 1.074286e+00
R30805 n0_4929_11217 n0_5866_11217 5.354286e+00
R30806 n0_5866_11217 n0_6054_11217 1.074286e+00
R30807 n0_6054_11217 n0_6991_11217 5.354286e+00
R30808 n0_6991_11217 n0_7179_11217 1.074286e+00
R30809 n0_7179_11217 n0_8116_11217 5.354286e+00
R30810 n0_8116_11217 n0_8304_11217 1.074286e+00
R30811 n0_8304_11217 n0_9241_11217 5.354286e+00
R30812 n0_9241_11217 n0_9429_11217 1.074286e+00
R30813 n0_9429_11217 n0_10366_11217 5.354286e+00
R30814 n0_10366_11217 n0_10458_11217 5.257143e-01
R30815 n0_10458_11217 n0_10554_11217 5.485714e-01
R30816 n0_10554_11217 n0_10646_11217 5.257143e-01
R30817 n0_10646_11217 n0_11491_11217 4.828571e+00
R30818 n0_11491_11217 n0_11679_11217 1.074286e+00
R30819 n0_11679_11217 n0_12616_11217 5.354286e+00
R30820 n0_12616_11217 n0_12804_11217 1.074286e+00
R30821 n0_12804_11217 n0_13741_11217 5.354286e+00
R30822 n0_13741_11217 n0_13929_11217 1.074286e+00
R30823 n0_13929_11217 n0_14866_11217 5.354286e+00
R30824 n0_14866_11217 n0_15054_11217 1.074286e+00
R30825 n0_15054_11217 n0_15991_11217 5.354286e+00
R30826 n0_15991_11217 n0_16179_11217 1.074286e+00
R30827 n0_16179_11217 n0_17116_11217 5.354286e+00
R30828 n0_17116_11217 n0_17304_11217 1.074286e+00
R30829 n0_17304_11217 n0_18241_11217 5.354286e+00
R30830 n0_18241_11217 n0_18429_11217 1.074286e+00
R30831 n0_18429_11217 n0_19366_11217 5.354286e+00
R30832 n0_19366_11217 n0_19554_11217 1.074286e+00
R30833 n0_241_11250 n0_429_11250 1.074286e+00
R30834 n0_429_11250 n0_1366_11250 5.354286e+00
R30835 n0_1366_11250 n0_1554_11250 1.074286e+00
R30836 n0_1554_11250 n0_2491_11250 5.354286e+00
R30837 n0_2491_11250 n0_2679_11250 1.074286e+00
R30838 n0_2679_11250 n0_3616_11250 5.354286e+00
R30839 n0_3616_11250 n0_3804_11250 1.074286e+00
R30840 n0_3804_11250 n0_4741_11250 5.354286e+00
R30841 n0_4741_11250 n0_4929_11250 1.074286e+00
R30842 n0_4929_11250 n0_5866_11250 5.354286e+00
R30843 n0_5866_11250 n0_6054_11250 1.074286e+00
R30844 n0_6054_11250 n0_6991_11250 5.354286e+00
R30845 n0_6991_11250 n0_7179_11250 1.074286e+00
R30846 n0_7179_11250 n0_8116_11250 5.354286e+00
R30847 n0_8116_11250 n0_8304_11250 1.074286e+00
R30848 n0_8304_11250 n0_9241_11250 5.354286e+00
R30849 n0_9241_11250 n0_9429_11250 1.074286e+00
R30850 n0_9429_11250 n0_10366_11250 5.354286e+00
R30851 n0_10366_11250 n0_10458_11250 5.257143e-01
R30852 n0_10458_11250 n0_10554_11250 5.485714e-01
R30853 n0_10554_11250 n0_10646_11250 5.257143e-01
R30854 n0_10646_11250 n0_11491_11250 4.828571e+00
R30855 n0_11491_11250 n0_11679_11250 1.074286e+00
R30856 n0_11679_11250 n0_12616_11250 5.354286e+00
R30857 n0_12616_11250 n0_12804_11250 1.074286e+00
R30858 n0_12804_11250 n0_13741_11250 5.354286e+00
R30859 n0_13741_11250 n0_13929_11250 1.074286e+00
R30860 n0_13929_11250 n0_14866_11250 5.354286e+00
R30861 n0_14866_11250 n0_15054_11250 1.074286e+00
R30862 n0_15054_11250 n0_15991_11250 5.354286e+00
R30863 n0_15991_11250 n0_16179_11250 1.074286e+00
R30864 n0_16179_11250 n0_17116_11250 5.354286e+00
R30865 n0_17116_11250 n0_17304_11250 1.074286e+00
R30866 n0_17304_11250 n0_18241_11250 5.354286e+00
R30867 n0_18241_11250 n0_18429_11250 1.074286e+00
R30868 n0_18429_11250 n0_19366_11250 5.354286e+00
R30869 n0_19366_11250 n0_19554_11250 1.074286e+00
R30870 n0_241_11433 n0_429_11433 1.074286e+00
R30871 n0_429_11433 n0_1366_11433 5.354286e+00
R30872 n0_1366_11433 n0_1554_11433 1.074286e+00
R30873 n0_1554_11433 n0_2491_11433 5.354286e+00
R30874 n0_2491_11433 n0_2679_11433 1.074286e+00
R30875 n0_2679_11433 n0_3616_11433 5.354286e+00
R30876 n0_3616_11433 n0_3804_11433 1.074286e+00
R30877 n0_3804_11433 n0_4741_11433 5.354286e+00
R30878 n0_4741_11433 n0_4929_11433 1.074286e+00
R30879 n0_4929_11433 n0_5866_11433 5.354286e+00
R30880 n0_5866_11433 n0_6054_11433 1.074286e+00
R30881 n0_6054_11433 n0_6991_11433 5.354286e+00
R30882 n0_6991_11433 n0_7179_11433 1.074286e+00
R30883 n0_7179_11433 n0_8116_11433 5.354286e+00
R30884 n0_8116_11433 n0_8304_11433 1.074286e+00
R30885 n0_8304_11433 n0_9241_11433 5.354286e+00
R30886 n0_9241_11433 n0_9429_11433 1.074286e+00
R30887 n0_9429_11433 n0_10366_11433 5.354286e+00
R30888 n0_10366_11433 n0_10458_11433 5.257143e-01
R30889 n0_10458_11433 n0_10554_11433 5.485714e-01
R30890 n0_10554_11433 n0_10646_11433 5.257143e-01
R30891 n0_10646_11433 n0_11491_11433 4.828571e+00
R30892 n0_11491_11433 n0_11679_11433 1.074286e+00
R30893 n0_11679_11433 n0_12616_11433 5.354286e+00
R30894 n0_12616_11433 n0_12804_11433 1.074286e+00
R30895 n0_12804_11433 n0_13741_11433 5.354286e+00
R30896 n0_13741_11433 n0_13929_11433 1.074286e+00
R30897 n0_13929_11433 n0_14866_11433 5.354286e+00
R30898 n0_14866_11433 n0_15054_11433 1.074286e+00
R30899 n0_15054_11433 n0_15991_11433 5.354286e+00
R30900 n0_15991_11433 n0_16179_11433 1.074286e+00
R30901 n0_16179_11433 n0_17116_11433 5.354286e+00
R30902 n0_17116_11433 n0_17304_11433 1.074286e+00
R30903 n0_17304_11433 n0_18241_11433 5.354286e+00
R30904 n0_18241_11433 n0_18429_11433 1.074286e+00
R30905 n0_18429_11433 n0_19366_11433 5.354286e+00
R30906 n0_19366_11433 n0_19554_11433 1.074286e+00
R30907 n0_241_11466 n0_429_11466 1.074286e+00
R30908 n0_429_11466 n0_1366_11466 5.354286e+00
R30909 n0_1366_11466 n0_1554_11466 1.074286e+00
R30910 n0_1554_11466 n0_2491_11466 5.354286e+00
R30911 n0_2491_11466 n0_2679_11466 1.074286e+00
R30912 n0_2679_11466 n0_3616_11466 5.354286e+00
R30913 n0_3616_11466 n0_3804_11466 1.074286e+00
R30914 n0_3804_11466 n0_4741_11466 5.354286e+00
R30915 n0_4741_11466 n0_4929_11466 1.074286e+00
R30916 n0_4929_11466 n0_5866_11466 5.354286e+00
R30917 n0_5866_11466 n0_6054_11466 1.074286e+00
R30918 n0_6054_11466 n0_6991_11466 5.354286e+00
R30919 n0_6991_11466 n0_7179_11466 1.074286e+00
R30920 n0_7179_11466 n0_8116_11466 5.354286e+00
R30921 n0_8116_11466 n0_8304_11466 1.074286e+00
R30922 n0_8304_11466 n0_9241_11466 5.354286e+00
R30923 n0_9241_11466 n0_9429_11466 1.074286e+00
R30924 n0_9429_11466 n0_10366_11466 5.354286e+00
R30925 n0_10366_11466 n0_10458_11466 5.257143e-01
R30926 n0_10458_11466 n0_10554_11466 5.485714e-01
R30927 n0_10554_11466 n0_10646_11466 5.257143e-01
R30928 n0_10646_11466 n0_11491_11466 4.828571e+00
R30929 n0_11491_11466 n0_11679_11466 1.074286e+00
R30930 n0_11679_11466 n0_12616_11466 5.354286e+00
R30931 n0_12616_11466 n0_12804_11466 1.074286e+00
R30932 n0_12804_11466 n0_13741_11466 5.354286e+00
R30933 n0_13741_11466 n0_13929_11466 1.074286e+00
R30934 n0_13929_11466 n0_14866_11466 5.354286e+00
R30935 n0_14866_11466 n0_15054_11466 1.074286e+00
R30936 n0_15054_11466 n0_15991_11466 5.354286e+00
R30937 n0_15991_11466 n0_16179_11466 1.074286e+00
R30938 n0_16179_11466 n0_17116_11466 5.354286e+00
R30939 n0_17116_11466 n0_17304_11466 1.074286e+00
R30940 n0_17304_11466 n0_18241_11466 5.354286e+00
R30941 n0_18241_11466 n0_18429_11466 1.074286e+00
R30942 n0_18429_11466 n0_19366_11466 5.354286e+00
R30943 n0_19366_11466 n0_19554_11466 1.074286e+00
R30944 n0_241_11649 n0_1366_11649 6.428571e+00
R30945 n0_1366_11649 n0_2491_11649 6.428571e+00
R30946 n0_2491_11649 n0_3616_11649 6.428571e+00
R30947 n0_3616_11649 n0_4741_11649 6.428571e+00
R30948 n0_4741_11649 n0_5866_11649 6.428571e+00
R30949 n0_5866_11649 n0_6991_11649 6.428571e+00
R30950 n0_6991_11649 n0_8116_11649 6.428571e+00
R30951 n0_8116_11649 n0_9241_11649 6.428571e+00
R30952 n0_9241_11649 n0_10366_11649 6.428571e+00
R30953 n0_10366_11649 n0_10458_11649 5.257143e-01
R30954 n0_10458_11649 n0_10505_11649 2.685714e-01
R30955 n0_10505_11649 n0_10554_11649 2.800000e-01
R30956 n0_10554_11649 n0_10646_11649 5.257143e-01
R30957 n0_10646_11649 n0_11491_11649 4.828571e+00
R30958 n0_11491_11649 n0_12616_11649 6.428571e+00
R30959 n0_12616_11649 n0_13741_11649 6.428571e+00
R30960 n0_13741_11649 n0_14866_11649 6.428571e+00
R30961 n0_14866_11649 n0_15991_11649 6.428571e+00
R30962 n0_15991_11649 n0_17116_11649 6.428571e+00
R30963 n0_17116_11649 n0_18241_11649 6.428571e+00
R30964 n0_18241_11649 n0_19366_11649 6.428571e+00
R30965 n0_241_11682 n0_1366_11682 6.428571e+00
R30966 n0_1366_11682 n0_2491_11682 6.428571e+00
R30967 n0_2491_11682 n0_3616_11682 6.428571e+00
R30968 n0_3616_11682 n0_4741_11682 6.428571e+00
R30969 n0_4741_11682 n0_5866_11682 6.428571e+00
R30970 n0_5866_11682 n0_6991_11682 6.428571e+00
R30971 n0_6991_11682 n0_8116_11682 6.428571e+00
R30972 n0_8116_11682 n0_9241_11682 6.428571e+00
R30973 n0_9241_11682 n0_10366_11682 6.428571e+00
R30974 n0_10366_11682 n0_10458_11682 5.257143e-01
R30975 n0_10458_11682 n0_10505_11682 2.685714e-01
R30976 n0_10505_11682 n0_10554_11682 2.800000e-01
R30977 n0_10554_11682 n0_10646_11682 5.257143e-01
R30978 n0_10646_11682 n0_11491_11682 4.828571e+00
R30979 n0_11491_11682 n0_12616_11682 6.428571e+00
R30980 n0_12616_11682 n0_13741_11682 6.428571e+00
R30981 n0_13741_11682 n0_14866_11682 6.428571e+00
R30982 n0_14866_11682 n0_15991_11682 6.428571e+00
R30983 n0_15991_11682 n0_17116_11682 6.428571e+00
R30984 n0_17116_11682 n0_18241_11682 6.428571e+00
R30985 n0_18241_11682 n0_19366_11682 6.428571e+00
R30986 n0_241_11865 n0_429_11865 1.074286e+00
R30987 n0_429_11865 n0_1366_11865 5.354286e+00
R30988 n0_1366_11865 n0_1554_11865 1.074286e+00
R30989 n0_1554_11865 n0_2491_11865 5.354286e+00
R30990 n0_2491_11865 n0_2679_11865 1.074286e+00
R30991 n0_2679_11865 n0_3616_11865 5.354286e+00
R30992 n0_3616_11865 n0_3804_11865 1.074286e+00
R30993 n0_3804_11865 n0_4741_11865 5.354286e+00
R30994 n0_4741_11865 n0_4929_11865 1.074286e+00
R30995 n0_4929_11865 n0_5866_11865 5.354286e+00
R30996 n0_5866_11865 n0_6054_11865 1.074286e+00
R30997 n0_6054_11865 n0_6991_11865 5.354286e+00
R30998 n0_6991_11865 n0_7179_11865 1.074286e+00
R30999 n0_7179_11865 n0_8116_11865 5.354286e+00
R31000 n0_8116_11865 n0_8304_11865 1.074286e+00
R31001 n0_8304_11865 n0_10366_11865 1.178286e+01
R31002 n0_10366_11865 n0_10458_11865 5.257143e-01
R31003 n0_10458_11865 n0_10554_11865 5.485714e-01
R31004 n0_10554_11865 n0_10646_11865 5.257143e-01
R31005 n0_10646_11865 n0_12616_11865 1.125714e+01
R31006 n0_12616_11865 n0_12804_11865 1.074286e+00
R31007 n0_12804_11865 n0_13741_11865 5.354286e+00
R31008 n0_13741_11865 n0_13929_11865 1.074286e+00
R31009 n0_13929_11865 n0_14866_11865 5.354286e+00
R31010 n0_14866_11865 n0_15054_11865 1.074286e+00
R31011 n0_15054_11865 n0_15991_11865 5.354286e+00
R31012 n0_15991_11865 n0_16179_11865 1.074286e+00
R31013 n0_16179_11865 n0_17116_11865 5.354286e+00
R31014 n0_17116_11865 n0_17304_11865 1.074286e+00
R31015 n0_17304_11865 n0_18241_11865 5.354286e+00
R31016 n0_18241_11865 n0_18429_11865 1.074286e+00
R31017 n0_18429_11865 n0_19366_11865 5.354286e+00
R31018 n0_19366_11865 n0_19554_11865 1.074286e+00
R31019 n0_241_11898 n0_429_11898 1.074286e+00
R31020 n0_429_11898 n0_1366_11898 5.354286e+00
R31021 n0_1366_11898 n0_1554_11898 1.074286e+00
R31022 n0_1554_11898 n0_2491_11898 5.354286e+00
R31023 n0_2491_11898 n0_2679_11898 1.074286e+00
R31024 n0_2679_11898 n0_3616_11898 5.354286e+00
R31025 n0_3616_11898 n0_3804_11898 1.074286e+00
R31026 n0_3804_11898 n0_4741_11898 5.354286e+00
R31027 n0_4741_11898 n0_4929_11898 1.074286e+00
R31028 n0_4929_11898 n0_5866_11898 5.354286e+00
R31029 n0_5866_11898 n0_6054_11898 1.074286e+00
R31030 n0_6054_11898 n0_6991_11898 5.354286e+00
R31031 n0_6991_11898 n0_7179_11898 1.074286e+00
R31032 n0_7179_11898 n0_8116_11898 5.354286e+00
R31033 n0_8116_11898 n0_8304_11898 1.074286e+00
R31034 n0_8304_11898 n0_10366_11898 1.178286e+01
R31035 n0_10366_11898 n0_10458_11898 5.257143e-01
R31036 n0_10458_11898 n0_10554_11898 5.485714e-01
R31037 n0_10554_11898 n0_10646_11898 5.257143e-01
R31038 n0_10646_11898 n0_12616_11898 1.125714e+01
R31039 n0_12616_11898 n0_12804_11898 1.074286e+00
R31040 n0_12804_11898 n0_13741_11898 5.354286e+00
R31041 n0_13741_11898 n0_13929_11898 1.074286e+00
R31042 n0_13929_11898 n0_14866_11898 5.354286e+00
R31043 n0_14866_11898 n0_15054_11898 1.074286e+00
R31044 n0_15054_11898 n0_15991_11898 5.354286e+00
R31045 n0_15991_11898 n0_16179_11898 1.074286e+00
R31046 n0_16179_11898 n0_17116_11898 5.354286e+00
R31047 n0_17116_11898 n0_17304_11898 1.074286e+00
R31048 n0_17304_11898 n0_18241_11898 5.354286e+00
R31049 n0_18241_11898 n0_18429_11898 1.074286e+00
R31050 n0_18429_11898 n0_19366_11898 5.354286e+00
R31051 n0_19366_11898 n0_19554_11898 1.074286e+00
R31052 n0_241_1098 n0_429_1098 1.074286e+00
R31053 n0_429_1098 n0_1366_1098 5.354286e+00
R31054 n0_1366_1098 n0_1458_1098 5.257143e-01
R31055 n0_1458_1098 n0_1554_1098 5.485714e-01
R31056 n0_1554_1098 n0_1646_1098 5.257143e-01
R31057 n0_1646_1098 n0_3616_1098 1.125714e+01
R31058 n0_3616_1098 n0_3708_1098 5.257143e-01
R31059 n0_3708_1098 n0_3804_1098 5.485714e-01
R31060 n0_3804_1098 n0_3896_1098 5.257143e-01
R31061 n0_3896_1098 n0_5866_1098 1.125714e+01
R31062 n0_5866_1098 n0_5958_1098 5.257143e-01
R31063 n0_5958_1098 n0_6054_1098 5.485714e-01
R31064 n0_6054_1098 n0_6146_1098 5.257143e-01
R31065 n0_6146_1098 n0_8116_1098 1.125714e+01
R31066 n0_8116_1098 n0_8208_1098 5.257143e-01
R31067 n0_8208_1098 n0_8304_1098 5.485714e-01
R31068 n0_8304_1098 n0_8396_1098 5.257143e-01
R31069 n0_8396_1098 n0_10366_1098 1.125714e+01
R31070 n0_10366_1098 n0_10458_1098 5.257143e-01
R31071 n0_10458_1098 n0_10554_1098 5.485714e-01
R31072 n0_10554_1098 n0_10646_1098 5.257143e-01
R31073 n0_10646_1098 n0_12616_1098 1.125714e+01
R31074 n0_12616_1098 n0_12708_1098 5.257143e-01
R31075 n0_12708_1098 n0_12804_1098 5.485714e-01
R31076 n0_12804_1098 n0_12896_1098 5.257143e-01
R31077 n0_12896_1098 n0_14866_1098 1.125714e+01
R31078 n0_14866_1098 n0_14958_1098 5.257143e-01
R31079 n0_14958_1098 n0_15054_1098 5.485714e-01
R31080 n0_15054_1098 n0_15146_1098 5.257143e-01
R31081 n0_15146_1098 n0_17116_1098 1.125714e+01
R31082 n0_17116_1098 n0_17208_1098 5.257143e-01
R31083 n0_17208_1098 n0_17304_1098 5.485714e-01
R31084 n0_17304_1098 n0_17396_1098 5.257143e-01
R31085 n0_17396_1098 n0_19366_1098 1.125714e+01
R31086 n0_19366_1098 n0_19458_1098 5.257143e-01
R31087 n0_19458_1098 n0_19554_1098 5.485714e-01
R31088 n0_19554_1098 n0_19646_1098 5.257143e-01
R31089 n0_19646_1098 n0_20491_1098 4.828571e+00
R31090 n0_20491_1098 n0_20679_1098 1.074286e+00
R31091 n0_241_1281 n0_429_1281 1.074286e+00
R31092 n0_429_1281 n0_1366_1281 5.354286e+00
R31093 n0_1366_1281 n0_1458_1281 5.257143e-01
R31094 n0_1458_1281 n0_1554_1281 5.485714e-01
R31095 n0_1554_1281 n0_1646_1281 5.257143e-01
R31096 n0_1646_1281 n0_3616_1281 1.125714e+01
R31097 n0_3616_1281 n0_3708_1281 5.257143e-01
R31098 n0_3708_1281 n0_3804_1281 5.485714e-01
R31099 n0_3804_1281 n0_3896_1281 5.257143e-01
R31100 n0_3896_1281 n0_5866_1281 1.125714e+01
R31101 n0_5866_1281 n0_5958_1281 5.257143e-01
R31102 n0_5958_1281 n0_6054_1281 5.485714e-01
R31103 n0_6054_1281 n0_6146_1281 5.257143e-01
R31104 n0_6146_1281 n0_8116_1281 1.125714e+01
R31105 n0_8116_1281 n0_8208_1281 5.257143e-01
R31106 n0_8208_1281 n0_8304_1281 5.485714e-01
R31107 n0_8304_1281 n0_8396_1281 5.257143e-01
R31108 n0_8396_1281 n0_10366_1281 1.125714e+01
R31109 n0_10366_1281 n0_10458_1281 5.257143e-01
R31110 n0_10458_1281 n0_10554_1281 5.485714e-01
R31111 n0_10554_1281 n0_10646_1281 5.257143e-01
R31112 n0_10646_1281 n0_12616_1281 1.125714e+01
R31113 n0_12616_1281 n0_12708_1281 5.257143e-01
R31114 n0_12708_1281 n0_12804_1281 5.485714e-01
R31115 n0_12804_1281 n0_12896_1281 5.257143e-01
R31116 n0_12896_1281 n0_14866_1281 1.125714e+01
R31117 n0_14866_1281 n0_14958_1281 5.257143e-01
R31118 n0_14958_1281 n0_15054_1281 5.485714e-01
R31119 n0_15054_1281 n0_15146_1281 5.257143e-01
R31120 n0_15146_1281 n0_17116_1281 1.125714e+01
R31121 n0_17116_1281 n0_17208_1281 5.257143e-01
R31122 n0_17208_1281 n0_17304_1281 5.485714e-01
R31123 n0_17304_1281 n0_17396_1281 5.257143e-01
R31124 n0_17396_1281 n0_19366_1281 1.125714e+01
R31125 n0_19366_1281 n0_19458_1281 5.257143e-01
R31126 n0_19458_1281 n0_19554_1281 5.485714e-01
R31127 n0_19554_1281 n0_19646_1281 5.257143e-01
R31128 n0_19646_1281 n0_20491_1281 4.828571e+00
R31129 n0_20491_1281 n0_20679_1281 1.074286e+00
R31130 n0_241_1314 n0_429_1314 1.074286e+00
R31131 n0_429_1314 n0_1366_1314 5.354286e+00
R31132 n0_1366_1314 n0_1458_1314 5.257143e-01
R31133 n0_1458_1314 n0_1554_1314 5.485714e-01
R31134 n0_1554_1314 n0_1646_1314 5.257143e-01
R31135 n0_1646_1314 n0_3616_1314 1.125714e+01
R31136 n0_3616_1314 n0_3708_1314 5.257143e-01
R31137 n0_3708_1314 n0_3804_1314 5.485714e-01
R31138 n0_3804_1314 n0_3896_1314 5.257143e-01
R31139 n0_3896_1314 n0_5866_1314 1.125714e+01
R31140 n0_5866_1314 n0_5958_1314 5.257143e-01
R31141 n0_5958_1314 n0_6054_1314 5.485714e-01
R31142 n0_6054_1314 n0_6146_1314 5.257143e-01
R31143 n0_6146_1314 n0_8116_1314 1.125714e+01
R31144 n0_8116_1314 n0_8208_1314 5.257143e-01
R31145 n0_8208_1314 n0_8304_1314 5.485714e-01
R31146 n0_8304_1314 n0_8396_1314 5.257143e-01
R31147 n0_8396_1314 n0_10366_1314 1.125714e+01
R31148 n0_10366_1314 n0_10458_1314 5.257143e-01
R31149 n0_10458_1314 n0_10554_1314 5.485714e-01
R31150 n0_10554_1314 n0_10646_1314 5.257143e-01
R31151 n0_10646_1314 n0_12616_1314 1.125714e+01
R31152 n0_12616_1314 n0_12708_1314 5.257143e-01
R31153 n0_12708_1314 n0_12804_1314 5.485714e-01
R31154 n0_12804_1314 n0_12896_1314 5.257143e-01
R31155 n0_12896_1314 n0_14866_1314 1.125714e+01
R31156 n0_14866_1314 n0_14958_1314 5.257143e-01
R31157 n0_14958_1314 n0_15054_1314 5.485714e-01
R31158 n0_15054_1314 n0_15146_1314 5.257143e-01
R31159 n0_15146_1314 n0_17116_1314 1.125714e+01
R31160 n0_17116_1314 n0_17208_1314 5.257143e-01
R31161 n0_17208_1314 n0_17304_1314 5.485714e-01
R31162 n0_17304_1314 n0_17396_1314 5.257143e-01
R31163 n0_17396_1314 n0_19366_1314 1.125714e+01
R31164 n0_19366_1314 n0_19458_1314 5.257143e-01
R31165 n0_19458_1314 n0_19554_1314 5.485714e-01
R31166 n0_19554_1314 n0_19646_1314 5.257143e-01
R31167 n0_19646_1314 n0_20491_1314 4.828571e+00
R31168 n0_20491_1314 n0_20679_1314 1.074286e+00
R31169 n0_241_1497 n0_429_1497 1.074286e+00
R31170 n0_429_1497 n0_1366_1497 5.354286e+00
R31171 n0_1366_1497 n0_1458_1497 5.257143e-01
R31172 n0_1458_1497 n0_1554_1497 5.485714e-01
R31173 n0_1554_1497 n0_1646_1497 5.257143e-01
R31174 n0_1646_1497 n0_3616_1497 1.125714e+01
R31175 n0_3616_1497 n0_3708_1497 5.257143e-01
R31176 n0_3708_1497 n0_3804_1497 5.485714e-01
R31177 n0_3804_1497 n0_3896_1497 5.257143e-01
R31178 n0_3896_1497 n0_5866_1497 1.125714e+01
R31179 n0_5866_1497 n0_5958_1497 5.257143e-01
R31180 n0_5958_1497 n0_6054_1497 5.485714e-01
R31181 n0_6054_1497 n0_6146_1497 5.257143e-01
R31182 n0_6146_1497 n0_8116_1497 1.125714e+01
R31183 n0_8116_1497 n0_8208_1497 5.257143e-01
R31184 n0_8208_1497 n0_8304_1497 5.485714e-01
R31185 n0_8304_1497 n0_8396_1497 5.257143e-01
R31186 n0_8396_1497 n0_10366_1497 1.125714e+01
R31187 n0_10366_1497 n0_10458_1497 5.257143e-01
R31188 n0_10458_1497 n0_10554_1497 5.485714e-01
R31189 n0_10554_1497 n0_10646_1497 5.257143e-01
R31190 n0_10646_1497 n0_12616_1497 1.125714e+01
R31191 n0_12616_1497 n0_12708_1497 5.257143e-01
R31192 n0_12708_1497 n0_12804_1497 5.485714e-01
R31193 n0_12804_1497 n0_12896_1497 5.257143e-01
R31194 n0_12896_1497 n0_14866_1497 1.125714e+01
R31195 n0_14866_1497 n0_14958_1497 5.257143e-01
R31196 n0_14958_1497 n0_15054_1497 5.485714e-01
R31197 n0_15054_1497 n0_15146_1497 5.257143e-01
R31198 n0_15146_1497 n0_17116_1497 1.125714e+01
R31199 n0_17116_1497 n0_17208_1497 5.257143e-01
R31200 n0_17208_1497 n0_17304_1497 5.485714e-01
R31201 n0_17304_1497 n0_17396_1497 5.257143e-01
R31202 n0_17396_1497 n0_19366_1497 1.125714e+01
R31203 n0_19366_1497 n0_19458_1497 5.257143e-01
R31204 n0_19458_1497 n0_19554_1497 5.485714e-01
R31205 n0_19554_1497 n0_19646_1497 5.257143e-01
R31206 n0_19646_1497 n0_20491_1497 4.828571e+00
R31207 n0_20491_1497 n0_20679_1497 1.074286e+00
R31208 n0_241_1530 n0_380_1530 7.942857e-01
R31209 n0_380_1530 n0_429_1530 2.800000e-01
R31210 n0_429_1530 n0_1366_1530 5.354286e+00
R31211 n0_1366_1530 n0_1646_1530 1.600000e+00
R31212 n0_1646_1530 n0_3616_1530 1.125714e+01
R31213 n0_3616_1530 n0_3708_1530 5.257143e-01
R31214 n0_3708_1530 n0_3755_1530 2.685714e-01
R31215 n0_3755_1530 n0_3804_1530 2.800000e-01
R31216 n0_3804_1530 n0_3896_1530 5.257143e-01
R31217 n0_3896_1530 n0_5866_1530 1.125714e+01
R31218 n0_5866_1530 n0_5958_1530 5.257143e-01
R31219 n0_5958_1530 n0_6005_1530 2.685714e-01
R31220 n0_6005_1530 n0_6054_1530 2.800000e-01
R31221 n0_6054_1530 n0_6146_1530 5.257143e-01
R31222 n0_6146_1530 n0_8116_1530 1.125714e+01
R31223 n0_8116_1530 n0_8208_1530 5.257143e-01
R31224 n0_8208_1530 n0_8255_1530 2.685714e-01
R31225 n0_8255_1530 n0_8304_1530 2.800000e-01
R31226 n0_8304_1530 n0_8396_1530 5.257143e-01
R31227 n0_8396_1530 n0_10366_1530 1.125714e+01
R31228 n0_10366_1530 n0_10458_1530 5.257143e-01
R31229 n0_10458_1530 n0_10505_1530 2.685714e-01
R31230 n0_10505_1530 n0_10554_1530 2.800000e-01
R31231 n0_10554_1530 n0_10646_1530 5.257143e-01
R31232 n0_10646_1530 n0_12616_1530 1.125714e+01
R31233 n0_12616_1530 n0_12708_1530 5.257143e-01
R31234 n0_12708_1530 n0_12755_1530 2.685714e-01
R31235 n0_12755_1530 n0_12804_1530 2.800000e-01
R31236 n0_12804_1530 n0_12896_1530 5.257143e-01
R31237 n0_12896_1530 n0_14866_1530 1.125714e+01
R31238 n0_14866_1530 n0_14958_1530 5.257143e-01
R31239 n0_14958_1530 n0_15005_1530 2.685714e-01
R31240 n0_15005_1530 n0_15054_1530 2.800000e-01
R31241 n0_15054_1530 n0_15146_1530 5.257143e-01
R31242 n0_15146_1530 n0_17116_1530 1.125714e+01
R31243 n0_17116_1530 n0_17208_1530 5.257143e-01
R31244 n0_17208_1530 n0_17255_1530 2.685714e-01
R31245 n0_17255_1530 n0_17304_1530 2.800000e-01
R31246 n0_17304_1530 n0_17396_1530 5.257143e-01
R31247 n0_17396_1530 n0_19366_1530 1.125714e+01
R31248 n0_19366_1530 n0_19646_1530 1.600000e+00
R31249 n0_19646_1530 n0_20491_1530 4.828571e+00
R31250 n0_20491_1530 n0_20630_1530 7.942857e-01
R31251 n0_20630_1530 n0_20679_1530 2.800000e-01
R31252 n0_241_1713 n0_429_1713 1.074286e+00
R31253 n0_429_1713 n0_1366_1713 5.354286e+00
R31254 n0_1366_1713 n0_1554_1713 1.074286e+00
R31255 n0_1554_1713 n0_3616_1713 1.178286e+01
R31256 n0_3616_1713 n0_3708_1713 5.257143e-01
R31257 n0_3708_1713 n0_3804_1713 5.485714e-01
R31258 n0_3804_1713 n0_3896_1713 5.257143e-01
R31259 n0_3896_1713 n0_5866_1713 1.125714e+01
R31260 n0_5866_1713 n0_5958_1713 5.257143e-01
R31261 n0_5958_1713 n0_6054_1713 5.485714e-01
R31262 n0_6054_1713 n0_6146_1713 5.257143e-01
R31263 n0_6146_1713 n0_8116_1713 1.125714e+01
R31264 n0_8116_1713 n0_8208_1713 5.257143e-01
R31265 n0_8208_1713 n0_8304_1713 5.485714e-01
R31266 n0_8304_1713 n0_8396_1713 5.257143e-01
R31267 n0_8396_1713 n0_10366_1713 1.125714e+01
R31268 n0_10366_1713 n0_10458_1713 5.257143e-01
R31269 n0_10458_1713 n0_10554_1713 5.485714e-01
R31270 n0_10554_1713 n0_10646_1713 5.257143e-01
R31271 n0_10646_1713 n0_12616_1713 1.125714e+01
R31272 n0_12616_1713 n0_12708_1713 5.257143e-01
R31273 n0_12708_1713 n0_12804_1713 5.485714e-01
R31274 n0_12804_1713 n0_12896_1713 5.257143e-01
R31275 n0_12896_1713 n0_14866_1713 1.125714e+01
R31276 n0_14866_1713 n0_14958_1713 5.257143e-01
R31277 n0_14958_1713 n0_15054_1713 5.485714e-01
R31278 n0_15054_1713 n0_15146_1713 5.257143e-01
R31279 n0_15146_1713 n0_17116_1713 1.125714e+01
R31280 n0_17116_1713 n0_17208_1713 5.257143e-01
R31281 n0_17208_1713 n0_17304_1713 5.485714e-01
R31282 n0_17304_1713 n0_17396_1713 5.257143e-01
R31283 n0_17396_1713 n0_19366_1713 1.125714e+01
R31284 n0_19366_1713 n0_19554_1713 1.074286e+00
R31285 n0_19554_1713 n0_20491_1713 5.354286e+00
R31286 n0_20491_1713 n0_20679_1713 1.074286e+00
R31287 n0_241_1746 n0_429_1746 1.074286e+00
R31288 n0_429_1746 n0_1366_1746 5.354286e+00
R31289 n0_1366_1746 n0_1554_1746 1.074286e+00
R31290 n0_1554_1746 n0_3616_1746 1.178286e+01
R31291 n0_3616_1746 n0_3708_1746 5.257143e-01
R31292 n0_3708_1746 n0_3804_1746 5.485714e-01
R31293 n0_3804_1746 n0_3896_1746 5.257143e-01
R31294 n0_3896_1746 n0_5866_1746 1.125714e+01
R31295 n0_5866_1746 n0_5958_1746 5.257143e-01
R31296 n0_5958_1746 n0_6054_1746 5.485714e-01
R31297 n0_6054_1746 n0_6146_1746 5.257143e-01
R31298 n0_6146_1746 n0_8116_1746 1.125714e+01
R31299 n0_8116_1746 n0_8208_1746 5.257143e-01
R31300 n0_8208_1746 n0_8304_1746 5.485714e-01
R31301 n0_8304_1746 n0_8396_1746 5.257143e-01
R31302 n0_8396_1746 n0_10366_1746 1.125714e+01
R31303 n0_10366_1746 n0_10458_1746 5.257143e-01
R31304 n0_10458_1746 n0_10554_1746 5.485714e-01
R31305 n0_10554_1746 n0_10646_1746 5.257143e-01
R31306 n0_10646_1746 n0_12616_1746 1.125714e+01
R31307 n0_12616_1746 n0_12708_1746 5.257143e-01
R31308 n0_12708_1746 n0_12804_1746 5.485714e-01
R31309 n0_12804_1746 n0_12896_1746 5.257143e-01
R31310 n0_12896_1746 n0_14866_1746 1.125714e+01
R31311 n0_14866_1746 n0_14958_1746 5.257143e-01
R31312 n0_14958_1746 n0_15054_1746 5.485714e-01
R31313 n0_15054_1746 n0_15146_1746 5.257143e-01
R31314 n0_15146_1746 n0_17116_1746 1.125714e+01
R31315 n0_17116_1746 n0_17208_1746 5.257143e-01
R31316 n0_17208_1746 n0_17304_1746 5.485714e-01
R31317 n0_17304_1746 n0_17396_1746 5.257143e-01
R31318 n0_17396_1746 n0_19366_1746 1.125714e+01
R31319 n0_19366_1746 n0_19554_1746 1.074286e+00
R31320 n0_19554_1746 n0_20491_1746 5.354286e+00
R31321 n0_20491_1746 n0_20679_1746 1.074286e+00
R31322 n0_241_1929 n0_429_1929 1.074286e+00
R31323 n0_429_1929 n0_1366_1929 5.354286e+00
R31324 n0_1366_1929 n0_1554_1929 1.074286e+00
R31325 n0_1554_1929 n0_3616_1929 1.178286e+01
R31326 n0_3616_1929 n0_3708_1929 5.257143e-01
R31327 n0_3708_1929 n0_3804_1929 5.485714e-01
R31328 n0_3804_1929 n0_3896_1929 5.257143e-01
R31329 n0_3896_1929 n0_5866_1929 1.125714e+01
R31330 n0_5866_1929 n0_5958_1929 5.257143e-01
R31331 n0_5958_1929 n0_6054_1929 5.485714e-01
R31332 n0_6054_1929 n0_6146_1929 5.257143e-01
R31333 n0_6146_1929 n0_8116_1929 1.125714e+01
R31334 n0_8116_1929 n0_8208_1929 5.257143e-01
R31335 n0_8208_1929 n0_8304_1929 5.485714e-01
R31336 n0_8304_1929 n0_8396_1929 5.257143e-01
R31337 n0_8396_1929 n0_10366_1929 1.125714e+01
R31338 n0_10366_1929 n0_10458_1929 5.257143e-01
R31339 n0_10458_1929 n0_10554_1929 5.485714e-01
R31340 n0_10554_1929 n0_10646_1929 5.257143e-01
R31341 n0_10646_1929 n0_12616_1929 1.125714e+01
R31342 n0_12616_1929 n0_12708_1929 5.257143e-01
R31343 n0_12708_1929 n0_12804_1929 5.485714e-01
R31344 n0_12804_1929 n0_12896_1929 5.257143e-01
R31345 n0_12896_1929 n0_14866_1929 1.125714e+01
R31346 n0_14866_1929 n0_14958_1929 5.257143e-01
R31347 n0_14958_1929 n0_15054_1929 5.485714e-01
R31348 n0_15054_1929 n0_15146_1929 5.257143e-01
R31349 n0_15146_1929 n0_17116_1929 1.125714e+01
R31350 n0_17116_1929 n0_17208_1929 5.257143e-01
R31351 n0_17208_1929 n0_17304_1929 5.485714e-01
R31352 n0_17304_1929 n0_17396_1929 5.257143e-01
R31353 n0_17396_1929 n0_19366_1929 1.125714e+01
R31354 n0_19366_1929 n0_19554_1929 1.074286e+00
R31355 n0_19554_1929 n0_20491_1929 5.354286e+00
R31356 n0_20491_1929 n0_20679_1929 1.074286e+00
R31357 n0_241_1962 n0_429_1962 1.074286e+00
R31358 n0_429_1962 n0_1366_1962 5.354286e+00
R31359 n0_1366_1962 n0_1554_1962 1.074286e+00
R31360 n0_1554_1962 n0_3616_1962 1.178286e+01
R31361 n0_3616_1962 n0_3708_1962 5.257143e-01
R31362 n0_3708_1962 n0_3804_1962 5.485714e-01
R31363 n0_3804_1962 n0_3896_1962 5.257143e-01
R31364 n0_3896_1962 n0_5866_1962 1.125714e+01
R31365 n0_5866_1962 n0_5958_1962 5.257143e-01
R31366 n0_5958_1962 n0_6054_1962 5.485714e-01
R31367 n0_6054_1962 n0_6146_1962 5.257143e-01
R31368 n0_6146_1962 n0_8116_1962 1.125714e+01
R31369 n0_8116_1962 n0_8208_1962 5.257143e-01
R31370 n0_8208_1962 n0_8304_1962 5.485714e-01
R31371 n0_8304_1962 n0_8396_1962 5.257143e-01
R31372 n0_8396_1962 n0_10366_1962 1.125714e+01
R31373 n0_10366_1962 n0_10458_1962 5.257143e-01
R31374 n0_10458_1962 n0_10554_1962 5.485714e-01
R31375 n0_10554_1962 n0_10646_1962 5.257143e-01
R31376 n0_10646_1962 n0_12616_1962 1.125714e+01
R31377 n0_12616_1962 n0_12708_1962 5.257143e-01
R31378 n0_12708_1962 n0_12804_1962 5.485714e-01
R31379 n0_12804_1962 n0_12896_1962 5.257143e-01
R31380 n0_12896_1962 n0_14866_1962 1.125714e+01
R31381 n0_14866_1962 n0_14958_1962 5.257143e-01
R31382 n0_14958_1962 n0_15054_1962 5.485714e-01
R31383 n0_15054_1962 n0_15146_1962 5.257143e-01
R31384 n0_15146_1962 n0_17116_1962 1.125714e+01
R31385 n0_17116_1962 n0_17208_1962 5.257143e-01
R31386 n0_17208_1962 n0_17304_1962 5.485714e-01
R31387 n0_17304_1962 n0_17396_1962 5.257143e-01
R31388 n0_17396_1962 n0_19366_1962 1.125714e+01
R31389 n0_19366_1962 n0_19554_1962 1.074286e+00
R31390 n0_19554_1962 n0_20491_1962 5.354286e+00
R31391 n0_20491_1962 n0_20679_1962 1.074286e+00
R31392 n0_241_2145 n0_429_2145 1.074286e+00
R31393 n0_429_2145 n0_1366_2145 5.354286e+00
R31394 n0_1366_2145 n0_1554_2145 1.074286e+00
R31395 n0_1554_2145 n0_3616_2145 1.178286e+01
R31396 n0_3616_2145 n0_3708_2145 5.257143e-01
R31397 n0_3708_2145 n0_3804_2145 5.485714e-01
R31398 n0_3804_2145 n0_3896_2145 5.257143e-01
R31399 n0_3896_2145 n0_5866_2145 1.125714e+01
R31400 n0_5866_2145 n0_5958_2145 5.257143e-01
R31401 n0_5958_2145 n0_6054_2145 5.485714e-01
R31402 n0_6054_2145 n0_6146_2145 5.257143e-01
R31403 n0_6146_2145 n0_8116_2145 1.125714e+01
R31404 n0_8116_2145 n0_8208_2145 5.257143e-01
R31405 n0_8208_2145 n0_8304_2145 5.485714e-01
R31406 n0_8304_2145 n0_8396_2145 5.257143e-01
R31407 n0_8396_2145 n0_10366_2145 1.125714e+01
R31408 n0_10366_2145 n0_10458_2145 5.257143e-01
R31409 n0_10458_2145 n0_10554_2145 5.485714e-01
R31410 n0_10554_2145 n0_10646_2145 5.257143e-01
R31411 n0_10646_2145 n0_12616_2145 1.125714e+01
R31412 n0_12616_2145 n0_12708_2145 5.257143e-01
R31413 n0_12708_2145 n0_12804_2145 5.485714e-01
R31414 n0_12804_2145 n0_12896_2145 5.257143e-01
R31415 n0_12896_2145 n0_14866_2145 1.125714e+01
R31416 n0_14866_2145 n0_14958_2145 5.257143e-01
R31417 n0_14958_2145 n0_15054_2145 5.485714e-01
R31418 n0_15054_2145 n0_15146_2145 5.257143e-01
R31419 n0_15146_2145 n0_17116_2145 1.125714e+01
R31420 n0_17116_2145 n0_17208_2145 5.257143e-01
R31421 n0_17208_2145 n0_17304_2145 5.485714e-01
R31422 n0_17304_2145 n0_17396_2145 5.257143e-01
R31423 n0_17396_2145 n0_19366_2145 1.125714e+01
R31424 n0_19366_2145 n0_19554_2145 1.074286e+00
R31425 n0_19554_2145 n0_20491_2145 5.354286e+00
R31426 n0_20491_2145 n0_20679_2145 1.074286e+00
R31427 n0_241_2178 n0_429_2178 1.074286e+00
R31428 n0_429_2178 n0_1366_2178 5.354286e+00
R31429 n0_1366_2178 n0_1554_2178 1.074286e+00
R31430 n0_1554_2178 n0_3616_2178 1.178286e+01
R31431 n0_3616_2178 n0_3708_2178 5.257143e-01
R31432 n0_3708_2178 n0_3804_2178 5.485714e-01
R31433 n0_3804_2178 n0_3896_2178 5.257143e-01
R31434 n0_3896_2178 n0_5866_2178 1.125714e+01
R31435 n0_5866_2178 n0_5958_2178 5.257143e-01
R31436 n0_5958_2178 n0_6054_2178 5.485714e-01
R31437 n0_6054_2178 n0_6146_2178 5.257143e-01
R31438 n0_6146_2178 n0_8116_2178 1.125714e+01
R31439 n0_8116_2178 n0_8208_2178 5.257143e-01
R31440 n0_8208_2178 n0_8304_2178 5.485714e-01
R31441 n0_8304_2178 n0_8396_2178 5.257143e-01
R31442 n0_8396_2178 n0_10366_2178 1.125714e+01
R31443 n0_10366_2178 n0_10458_2178 5.257143e-01
R31444 n0_10458_2178 n0_10554_2178 5.485714e-01
R31445 n0_10554_2178 n0_10646_2178 5.257143e-01
R31446 n0_10646_2178 n0_12616_2178 1.125714e+01
R31447 n0_12616_2178 n0_12708_2178 5.257143e-01
R31448 n0_12708_2178 n0_12804_2178 5.485714e-01
R31449 n0_12804_2178 n0_12896_2178 5.257143e-01
R31450 n0_12896_2178 n0_14866_2178 1.125714e+01
R31451 n0_14866_2178 n0_14958_2178 5.257143e-01
R31452 n0_14958_2178 n0_15054_2178 5.485714e-01
R31453 n0_15054_2178 n0_15146_2178 5.257143e-01
R31454 n0_15146_2178 n0_17116_2178 1.125714e+01
R31455 n0_17116_2178 n0_17208_2178 5.257143e-01
R31456 n0_17208_2178 n0_17304_2178 5.485714e-01
R31457 n0_17304_2178 n0_17396_2178 5.257143e-01
R31458 n0_17396_2178 n0_19366_2178 1.125714e+01
R31459 n0_19366_2178 n0_19554_2178 1.074286e+00
R31460 n0_19554_2178 n0_20491_2178 5.354286e+00
R31461 n0_20491_2178 n0_20679_2178 1.074286e+00
R31462 n0_241_2361 n0_429_2361 1.074286e+00
R31463 n0_429_2361 n0_1366_2361 5.354286e+00
R31464 n0_1366_2361 n0_1554_2361 1.074286e+00
R31465 n0_1554_2361 n0_3616_2361 1.178286e+01
R31466 n0_3616_2361 n0_3708_2361 5.257143e-01
R31467 n0_3708_2361 n0_3804_2361 5.485714e-01
R31468 n0_3804_2361 n0_3896_2361 5.257143e-01
R31469 n0_3896_2361 n0_5866_2361 1.125714e+01
R31470 n0_5866_2361 n0_5958_2361 5.257143e-01
R31471 n0_5958_2361 n0_6054_2361 5.485714e-01
R31472 n0_6054_2361 n0_6146_2361 5.257143e-01
R31473 n0_6146_2361 n0_8116_2361 1.125714e+01
R31474 n0_8116_2361 n0_8208_2361 5.257143e-01
R31475 n0_8208_2361 n0_8304_2361 5.485714e-01
R31476 n0_8304_2361 n0_8396_2361 5.257143e-01
R31477 n0_8396_2361 n0_10366_2361 1.125714e+01
R31478 n0_10366_2361 n0_10458_2361 5.257143e-01
R31479 n0_10458_2361 n0_10554_2361 5.485714e-01
R31480 n0_10554_2361 n0_10646_2361 5.257143e-01
R31481 n0_10646_2361 n0_12616_2361 1.125714e+01
R31482 n0_12616_2361 n0_12708_2361 5.257143e-01
R31483 n0_12708_2361 n0_12804_2361 5.485714e-01
R31484 n0_12804_2361 n0_12896_2361 5.257143e-01
R31485 n0_12896_2361 n0_14866_2361 1.125714e+01
R31486 n0_14866_2361 n0_14958_2361 5.257143e-01
R31487 n0_14958_2361 n0_15054_2361 5.485714e-01
R31488 n0_15054_2361 n0_15146_2361 5.257143e-01
R31489 n0_15146_2361 n0_17116_2361 1.125714e+01
R31490 n0_17116_2361 n0_17208_2361 5.257143e-01
R31491 n0_17208_2361 n0_17304_2361 5.485714e-01
R31492 n0_17304_2361 n0_17396_2361 5.257143e-01
R31493 n0_17396_2361 n0_19366_2361 1.125714e+01
R31494 n0_19366_2361 n0_19554_2361 1.074286e+00
R31495 n0_19554_2361 n0_20491_2361 5.354286e+00
R31496 n0_20491_2361 n0_20679_2361 1.074286e+00
R31497 n0_241_2394 n0_429_2394 1.074286e+00
R31498 n0_429_2394 n0_1366_2394 5.354286e+00
R31499 n0_1366_2394 n0_1554_2394 1.074286e+00
R31500 n0_1554_2394 n0_3616_2394 1.178286e+01
R31501 n0_3616_2394 n0_3708_2394 5.257143e-01
R31502 n0_3708_2394 n0_3804_2394 5.485714e-01
R31503 n0_3804_2394 n0_3896_2394 5.257143e-01
R31504 n0_3896_2394 n0_5866_2394 1.125714e+01
R31505 n0_5866_2394 n0_5958_2394 5.257143e-01
R31506 n0_5958_2394 n0_6054_2394 5.485714e-01
R31507 n0_6054_2394 n0_6146_2394 5.257143e-01
R31508 n0_6146_2394 n0_8116_2394 1.125714e+01
R31509 n0_8116_2394 n0_8208_2394 5.257143e-01
R31510 n0_8208_2394 n0_8304_2394 5.485714e-01
R31511 n0_8304_2394 n0_8396_2394 5.257143e-01
R31512 n0_8396_2394 n0_10366_2394 1.125714e+01
R31513 n0_10366_2394 n0_10458_2394 5.257143e-01
R31514 n0_10458_2394 n0_10554_2394 5.485714e-01
R31515 n0_10554_2394 n0_10646_2394 5.257143e-01
R31516 n0_10646_2394 n0_12616_2394 1.125714e+01
R31517 n0_12616_2394 n0_12708_2394 5.257143e-01
R31518 n0_12708_2394 n0_12804_2394 5.485714e-01
R31519 n0_12804_2394 n0_12896_2394 5.257143e-01
R31520 n0_12896_2394 n0_14866_2394 1.125714e+01
R31521 n0_14866_2394 n0_14958_2394 5.257143e-01
R31522 n0_14958_2394 n0_15054_2394 5.485714e-01
R31523 n0_15054_2394 n0_15146_2394 5.257143e-01
R31524 n0_15146_2394 n0_17116_2394 1.125714e+01
R31525 n0_17116_2394 n0_17208_2394 5.257143e-01
R31526 n0_17208_2394 n0_17304_2394 5.485714e-01
R31527 n0_17304_2394 n0_17396_2394 5.257143e-01
R31528 n0_17396_2394 n0_19366_2394 1.125714e+01
R31529 n0_19366_2394 n0_19554_2394 1.074286e+00
R31530 n0_19554_2394 n0_20491_2394 5.354286e+00
R31531 n0_20491_2394 n0_20679_2394 1.074286e+00
R31532 n0_241_2577 n0_429_2577 1.074286e+00
R31533 n0_429_2577 n0_1366_2577 5.354286e+00
R31534 n0_1366_2577 n0_1554_2577 1.074286e+00
R31535 n0_1554_2577 n0_3616_2577 1.178286e+01
R31536 n0_3616_2577 n0_3708_2577 5.257143e-01
R31537 n0_3708_2577 n0_3804_2577 5.485714e-01
R31538 n0_3804_2577 n0_3896_2577 5.257143e-01
R31539 n0_3896_2577 n0_5866_2577 1.125714e+01
R31540 n0_5866_2577 n0_5958_2577 5.257143e-01
R31541 n0_5958_2577 n0_6054_2577 5.485714e-01
R31542 n0_6054_2577 n0_6146_2577 5.257143e-01
R31543 n0_6146_2577 n0_8116_2577 1.125714e+01
R31544 n0_8116_2577 n0_8208_2577 5.257143e-01
R31545 n0_8208_2577 n0_8304_2577 5.485714e-01
R31546 n0_8304_2577 n0_8396_2577 5.257143e-01
R31547 n0_8396_2577 n0_10366_2577 1.125714e+01
R31548 n0_10366_2577 n0_10458_2577 5.257143e-01
R31549 n0_10458_2577 n0_10554_2577 5.485714e-01
R31550 n0_10554_2577 n0_10646_2577 5.257143e-01
R31551 n0_10646_2577 n0_12616_2577 1.125714e+01
R31552 n0_12616_2577 n0_12708_2577 5.257143e-01
R31553 n0_12708_2577 n0_12804_2577 5.485714e-01
R31554 n0_12804_2577 n0_12896_2577 5.257143e-01
R31555 n0_12896_2577 n0_14866_2577 1.125714e+01
R31556 n0_14866_2577 n0_14958_2577 5.257143e-01
R31557 n0_14958_2577 n0_15054_2577 5.485714e-01
R31558 n0_15054_2577 n0_15146_2577 5.257143e-01
R31559 n0_15146_2577 n0_17116_2577 1.125714e+01
R31560 n0_17116_2577 n0_17208_2577 5.257143e-01
R31561 n0_17208_2577 n0_17304_2577 5.485714e-01
R31562 n0_17304_2577 n0_17396_2577 5.257143e-01
R31563 n0_17396_2577 n0_19366_2577 1.125714e+01
R31564 n0_19366_2577 n0_19554_2577 1.074286e+00
R31565 n0_19554_2577 n0_20491_2577 5.354286e+00
R31566 n0_20491_2577 n0_20679_2577 1.074286e+00
R31567 n0_241_2610 n0_429_2610 1.074286e+00
R31568 n0_429_2610 n0_1366_2610 5.354286e+00
R31569 n0_1366_2610 n0_1554_2610 1.074286e+00
R31570 n0_1554_2610 n0_3616_2610 1.178286e+01
R31571 n0_3616_2610 n0_3708_2610 5.257143e-01
R31572 n0_3708_2610 n0_3804_2610 5.485714e-01
R31573 n0_3804_2610 n0_3896_2610 5.257143e-01
R31574 n0_3896_2610 n0_5866_2610 1.125714e+01
R31575 n0_5866_2610 n0_5958_2610 5.257143e-01
R31576 n0_5958_2610 n0_6054_2610 5.485714e-01
R31577 n0_6054_2610 n0_6146_2610 5.257143e-01
R31578 n0_6146_2610 n0_8116_2610 1.125714e+01
R31579 n0_8116_2610 n0_8208_2610 5.257143e-01
R31580 n0_8208_2610 n0_8304_2610 5.485714e-01
R31581 n0_8304_2610 n0_8396_2610 5.257143e-01
R31582 n0_8396_2610 n0_10366_2610 1.125714e+01
R31583 n0_10366_2610 n0_10458_2610 5.257143e-01
R31584 n0_10458_2610 n0_10554_2610 5.485714e-01
R31585 n0_10554_2610 n0_10646_2610 5.257143e-01
R31586 n0_10646_2610 n0_12616_2610 1.125714e+01
R31587 n0_12616_2610 n0_12708_2610 5.257143e-01
R31588 n0_12708_2610 n0_12804_2610 5.485714e-01
R31589 n0_12804_2610 n0_12896_2610 5.257143e-01
R31590 n0_12896_2610 n0_14866_2610 1.125714e+01
R31591 n0_14866_2610 n0_14958_2610 5.257143e-01
R31592 n0_14958_2610 n0_15054_2610 5.485714e-01
R31593 n0_15054_2610 n0_15146_2610 5.257143e-01
R31594 n0_15146_2610 n0_17116_2610 1.125714e+01
R31595 n0_17116_2610 n0_17208_2610 5.257143e-01
R31596 n0_17208_2610 n0_17304_2610 5.485714e-01
R31597 n0_17304_2610 n0_17396_2610 5.257143e-01
R31598 n0_17396_2610 n0_19366_2610 1.125714e+01
R31599 n0_19366_2610 n0_19554_2610 1.074286e+00
R31600 n0_19554_2610 n0_20491_2610 5.354286e+00
R31601 n0_20491_2610 n0_20679_2610 1.074286e+00
R31602 n0_241_2793 n0_1366_2793 6.428571e+00
R31603 n0_1366_2793 n0_2491_2793 6.428571e+00
R31604 n0_2491_2793 n0_3616_2793 6.428571e+00
R31605 n0_3616_2793 n0_3708_2793 5.257143e-01
R31606 n0_3708_2793 n0_3755_2793 2.685714e-01
R31607 n0_3755_2793 n0_3804_2793 2.800000e-01
R31608 n0_3804_2793 n0_3896_2793 5.257143e-01
R31609 n0_3896_2793 n0_5866_2793 1.125714e+01
R31610 n0_5866_2793 n0_5958_2793 5.257143e-01
R31611 n0_5958_2793 n0_6005_2793 2.685714e-01
R31612 n0_6005_2793 n0_6054_2793 2.800000e-01
R31613 n0_6054_2793 n0_6146_2793 5.257143e-01
R31614 n0_6146_2793 n0_8116_2793 1.125714e+01
R31615 n0_8116_2793 n0_8208_2793 5.257143e-01
R31616 n0_8208_2793 n0_8255_2793 2.685714e-01
R31617 n0_8255_2793 n0_8304_2793 2.800000e-01
R31618 n0_8304_2793 n0_8396_2793 5.257143e-01
R31619 n0_8396_2793 n0_10366_2793 1.125714e+01
R31620 n0_10366_2793 n0_10458_2793 5.257143e-01
R31621 n0_10458_2793 n0_10505_2793 2.685714e-01
R31622 n0_10505_2793 n0_10554_2793 2.800000e-01
R31623 n0_10554_2793 n0_10646_2793 5.257143e-01
R31624 n0_10646_2793 n0_12616_2793 1.125714e+01
R31625 n0_12616_2793 n0_12708_2793 5.257143e-01
R31626 n0_12708_2793 n0_12755_2793 2.685714e-01
R31627 n0_12755_2793 n0_12804_2793 2.800000e-01
R31628 n0_12804_2793 n0_12896_2793 5.257143e-01
R31629 n0_12896_2793 n0_14866_2793 1.125714e+01
R31630 n0_14866_2793 n0_14958_2793 5.257143e-01
R31631 n0_14958_2793 n0_15005_2793 2.685714e-01
R31632 n0_15005_2793 n0_15054_2793 2.800000e-01
R31633 n0_15054_2793 n0_15146_2793 5.257143e-01
R31634 n0_15146_2793 n0_17116_2793 1.125714e+01
R31635 n0_17116_2793 n0_17208_2793 5.257143e-01
R31636 n0_17208_2793 n0_17255_2793 2.685714e-01
R31637 n0_17255_2793 n0_17304_2793 2.800000e-01
R31638 n0_17304_2793 n0_17396_2793 5.257143e-01
R31639 n0_17396_2793 n0_18241_2793 4.828571e+00
R31640 n0_18241_2793 n0_19366_2793 6.428571e+00
R31641 n0_19366_2793 n0_20491_2793 6.428571e+00
R31642 n0_241_2826 n0_429_2826 1.074286e+00
R31643 n0_429_2826 n0_1366_2826 5.354286e+00
R31644 n0_1366_2826 n0_1554_2826 1.074286e+00
R31645 n0_1554_2826 n0_2491_2826 5.354286e+00
R31646 n0_2491_2826 n0_2679_2826 1.074286e+00
R31647 n0_2679_2826 n0_3616_2826 5.354286e+00
R31648 n0_3616_2826 n0_3708_2826 5.257143e-01
R31649 n0_3708_2826 n0_3804_2826 5.485714e-01
R31650 n0_3804_2826 n0_3896_2826 5.257143e-01
R31651 n0_3896_2826 n0_5866_2826 1.125714e+01
R31652 n0_5866_2826 n0_5958_2826 5.257143e-01
R31653 n0_5958_2826 n0_6054_2826 5.485714e-01
R31654 n0_6054_2826 n0_6146_2826 5.257143e-01
R31655 n0_6146_2826 n0_8116_2826 1.125714e+01
R31656 n0_8116_2826 n0_8208_2826 5.257143e-01
R31657 n0_8208_2826 n0_8304_2826 5.485714e-01
R31658 n0_8304_2826 n0_8396_2826 5.257143e-01
R31659 n0_8396_2826 n0_10366_2826 1.125714e+01
R31660 n0_10366_2826 n0_10458_2826 5.257143e-01
R31661 n0_10458_2826 n0_10554_2826 5.485714e-01
R31662 n0_10554_2826 n0_10646_2826 5.257143e-01
R31663 n0_10646_2826 n0_12616_2826 1.125714e+01
R31664 n0_12616_2826 n0_12708_2826 5.257143e-01
R31665 n0_12708_2826 n0_12804_2826 5.485714e-01
R31666 n0_12804_2826 n0_12896_2826 5.257143e-01
R31667 n0_12896_2826 n0_14866_2826 1.125714e+01
R31668 n0_14866_2826 n0_14958_2826 5.257143e-01
R31669 n0_14958_2826 n0_15054_2826 5.485714e-01
R31670 n0_15054_2826 n0_15146_2826 5.257143e-01
R31671 n0_15146_2826 n0_17116_2826 1.125714e+01
R31672 n0_17116_2826 n0_17208_2826 5.257143e-01
R31673 n0_17208_2826 n0_17304_2826 5.485714e-01
R31674 n0_17304_2826 n0_17396_2826 5.257143e-01
R31675 n0_17396_2826 n0_18241_2826 4.828571e+00
R31676 n0_18241_2826 n0_18429_2826 1.074286e+00
R31677 n0_18429_2826 n0_19366_2826 5.354286e+00
R31678 n0_19366_2826 n0_19554_2826 1.074286e+00
R31679 n0_19554_2826 n0_20491_2826 5.354286e+00
R31680 n0_20491_2826 n0_20679_2826 1.074286e+00
R31681 n0_241_3009 n0_429_3009 1.074286e+00
R31682 n0_429_3009 n0_1366_3009 5.354286e+00
R31683 n0_1366_3009 n0_1554_3009 1.074286e+00
R31684 n0_1554_3009 n0_2491_3009 5.354286e+00
R31685 n0_2491_3009 n0_2679_3009 1.074286e+00
R31686 n0_2679_3009 n0_3616_3009 5.354286e+00
R31687 n0_3616_3009 n0_3708_3009 5.257143e-01
R31688 n0_3708_3009 n0_3804_3009 5.485714e-01
R31689 n0_3804_3009 n0_3896_3009 5.257143e-01
R31690 n0_3896_3009 n0_5866_3009 1.125714e+01
R31691 n0_5866_3009 n0_5958_3009 5.257143e-01
R31692 n0_5958_3009 n0_6054_3009 5.485714e-01
R31693 n0_6054_3009 n0_6146_3009 5.257143e-01
R31694 n0_6146_3009 n0_8116_3009 1.125714e+01
R31695 n0_8116_3009 n0_8208_3009 5.257143e-01
R31696 n0_8208_3009 n0_8304_3009 5.485714e-01
R31697 n0_8304_3009 n0_8396_3009 5.257143e-01
R31698 n0_8396_3009 n0_10366_3009 1.125714e+01
R31699 n0_10366_3009 n0_10458_3009 5.257143e-01
R31700 n0_10458_3009 n0_10554_3009 5.485714e-01
R31701 n0_10554_3009 n0_10646_3009 5.257143e-01
R31702 n0_10646_3009 n0_12616_3009 1.125714e+01
R31703 n0_12616_3009 n0_12708_3009 5.257143e-01
R31704 n0_12708_3009 n0_12804_3009 5.485714e-01
R31705 n0_12804_3009 n0_12896_3009 5.257143e-01
R31706 n0_12896_3009 n0_14866_3009 1.125714e+01
R31707 n0_14866_3009 n0_14958_3009 5.257143e-01
R31708 n0_14958_3009 n0_15054_3009 5.485714e-01
R31709 n0_15054_3009 n0_15146_3009 5.257143e-01
R31710 n0_15146_3009 n0_17116_3009 1.125714e+01
R31711 n0_17116_3009 n0_17208_3009 5.257143e-01
R31712 n0_17208_3009 n0_17304_3009 5.485714e-01
R31713 n0_17304_3009 n0_17396_3009 5.257143e-01
R31714 n0_17396_3009 n0_18241_3009 4.828571e+00
R31715 n0_18241_3009 n0_18429_3009 1.074286e+00
R31716 n0_18429_3009 n0_19366_3009 5.354286e+00
R31717 n0_19366_3009 n0_19554_3009 1.074286e+00
R31718 n0_19554_3009 n0_20491_3009 5.354286e+00
R31719 n0_20491_3009 n0_20679_3009 1.074286e+00
R31720 n0_241_3042 n0_429_3042 1.074286e+00
R31721 n0_429_3042 n0_1366_3042 5.354286e+00
R31722 n0_1366_3042 n0_1554_3042 1.074286e+00
R31723 n0_1554_3042 n0_2491_3042 5.354286e+00
R31724 n0_2491_3042 n0_2679_3042 1.074286e+00
R31725 n0_2679_3042 n0_3616_3042 5.354286e+00
R31726 n0_3616_3042 n0_3708_3042 5.257143e-01
R31727 n0_3708_3042 n0_3804_3042 5.485714e-01
R31728 n0_3804_3042 n0_3896_3042 5.257143e-01
R31729 n0_3896_3042 n0_5866_3042 1.125714e+01
R31730 n0_5866_3042 n0_5958_3042 5.257143e-01
R31731 n0_5958_3042 n0_6054_3042 5.485714e-01
R31732 n0_6054_3042 n0_6146_3042 5.257143e-01
R31733 n0_6146_3042 n0_8116_3042 1.125714e+01
R31734 n0_8116_3042 n0_8208_3042 5.257143e-01
R31735 n0_8208_3042 n0_8304_3042 5.485714e-01
R31736 n0_8304_3042 n0_8396_3042 5.257143e-01
R31737 n0_8396_3042 n0_10366_3042 1.125714e+01
R31738 n0_10366_3042 n0_10458_3042 5.257143e-01
R31739 n0_10458_3042 n0_10554_3042 5.485714e-01
R31740 n0_10554_3042 n0_10646_3042 5.257143e-01
R31741 n0_10646_3042 n0_12616_3042 1.125714e+01
R31742 n0_12616_3042 n0_12708_3042 5.257143e-01
R31743 n0_12708_3042 n0_12804_3042 5.485714e-01
R31744 n0_12804_3042 n0_12896_3042 5.257143e-01
R31745 n0_12896_3042 n0_14866_3042 1.125714e+01
R31746 n0_14866_3042 n0_14958_3042 5.257143e-01
R31747 n0_14958_3042 n0_15054_3042 5.485714e-01
R31748 n0_15054_3042 n0_15146_3042 5.257143e-01
R31749 n0_15146_3042 n0_17116_3042 1.125714e+01
R31750 n0_17116_3042 n0_17208_3042 5.257143e-01
R31751 n0_17208_3042 n0_17304_3042 5.485714e-01
R31752 n0_17304_3042 n0_17396_3042 5.257143e-01
R31753 n0_17396_3042 n0_18241_3042 4.828571e+00
R31754 n0_18241_3042 n0_18429_3042 1.074286e+00
R31755 n0_18429_3042 n0_19366_3042 5.354286e+00
R31756 n0_19366_3042 n0_19554_3042 1.074286e+00
R31757 n0_19554_3042 n0_20491_3042 5.354286e+00
R31758 n0_20491_3042 n0_20679_3042 1.074286e+00
R31759 n0_241_3225 n0_429_3225 1.074286e+00
R31760 n0_429_3225 n0_1366_3225 5.354286e+00
R31761 n0_1366_3225 n0_1554_3225 1.074286e+00
R31762 n0_1554_3225 n0_2491_3225 5.354286e+00
R31763 n0_2491_3225 n0_2679_3225 1.074286e+00
R31764 n0_2679_3225 n0_3616_3225 5.354286e+00
R31765 n0_3616_3225 n0_3708_3225 5.257143e-01
R31766 n0_3708_3225 n0_3804_3225 5.485714e-01
R31767 n0_3804_3225 n0_3896_3225 5.257143e-01
R31768 n0_3896_3225 n0_5866_3225 1.125714e+01
R31769 n0_5866_3225 n0_5958_3225 5.257143e-01
R31770 n0_5958_3225 n0_6054_3225 5.485714e-01
R31771 n0_6054_3225 n0_6146_3225 5.257143e-01
R31772 n0_6146_3225 n0_8116_3225 1.125714e+01
R31773 n0_8116_3225 n0_8208_3225 5.257143e-01
R31774 n0_8208_3225 n0_8304_3225 5.485714e-01
R31775 n0_8304_3225 n0_8396_3225 5.257143e-01
R31776 n0_8396_3225 n0_10366_3225 1.125714e+01
R31777 n0_10366_3225 n0_10458_3225 5.257143e-01
R31778 n0_10458_3225 n0_10554_3225 5.485714e-01
R31779 n0_10554_3225 n0_10646_3225 5.257143e-01
R31780 n0_10646_3225 n0_12616_3225 1.125714e+01
R31781 n0_12616_3225 n0_12708_3225 5.257143e-01
R31782 n0_12708_3225 n0_12804_3225 5.485714e-01
R31783 n0_12804_3225 n0_12896_3225 5.257143e-01
R31784 n0_12896_3225 n0_14866_3225 1.125714e+01
R31785 n0_14866_3225 n0_14958_3225 5.257143e-01
R31786 n0_14958_3225 n0_15054_3225 5.485714e-01
R31787 n0_15054_3225 n0_15146_3225 5.257143e-01
R31788 n0_15146_3225 n0_17116_3225 1.125714e+01
R31789 n0_17116_3225 n0_17208_3225 5.257143e-01
R31790 n0_17208_3225 n0_17304_3225 5.485714e-01
R31791 n0_17304_3225 n0_17396_3225 5.257143e-01
R31792 n0_17396_3225 n0_18241_3225 4.828571e+00
R31793 n0_18241_3225 n0_18429_3225 1.074286e+00
R31794 n0_18429_3225 n0_19366_3225 5.354286e+00
R31795 n0_19366_3225 n0_19554_3225 1.074286e+00
R31796 n0_19554_3225 n0_20491_3225 5.354286e+00
R31797 n0_20491_3225 n0_20679_3225 1.074286e+00
R31798 n0_241_3258 n0_429_3258 1.074286e+00
R31799 n0_429_3258 n0_1366_3258 5.354286e+00
R31800 n0_1366_3258 n0_1554_3258 1.074286e+00
R31801 n0_1554_3258 n0_2491_3258 5.354286e+00
R31802 n0_2491_3258 n0_2679_3258 1.074286e+00
R31803 n0_2679_3258 n0_3616_3258 5.354286e+00
R31804 n0_3616_3258 n0_3708_3258 5.257143e-01
R31805 n0_3708_3258 n0_3804_3258 5.485714e-01
R31806 n0_3804_3258 n0_3896_3258 5.257143e-01
R31807 n0_3896_3258 n0_5866_3258 1.125714e+01
R31808 n0_5866_3258 n0_5958_3258 5.257143e-01
R31809 n0_5958_3258 n0_6054_3258 5.485714e-01
R31810 n0_6054_3258 n0_6146_3258 5.257143e-01
R31811 n0_6146_3258 n0_8116_3258 1.125714e+01
R31812 n0_8116_3258 n0_8208_3258 5.257143e-01
R31813 n0_8208_3258 n0_8304_3258 5.485714e-01
R31814 n0_8304_3258 n0_8396_3258 5.257143e-01
R31815 n0_8396_3258 n0_10366_3258 1.125714e+01
R31816 n0_10366_3258 n0_10458_3258 5.257143e-01
R31817 n0_10458_3258 n0_10554_3258 5.485714e-01
R31818 n0_10554_3258 n0_10646_3258 5.257143e-01
R31819 n0_10646_3258 n0_12616_3258 1.125714e+01
R31820 n0_12616_3258 n0_12708_3258 5.257143e-01
R31821 n0_12708_3258 n0_12804_3258 5.485714e-01
R31822 n0_12804_3258 n0_12896_3258 5.257143e-01
R31823 n0_12896_3258 n0_14866_3258 1.125714e+01
R31824 n0_14866_3258 n0_14958_3258 5.257143e-01
R31825 n0_14958_3258 n0_15054_3258 5.485714e-01
R31826 n0_15054_3258 n0_15146_3258 5.257143e-01
R31827 n0_15146_3258 n0_17116_3258 1.125714e+01
R31828 n0_17116_3258 n0_17208_3258 5.257143e-01
R31829 n0_17208_3258 n0_17304_3258 5.485714e-01
R31830 n0_17304_3258 n0_17396_3258 5.257143e-01
R31831 n0_17396_3258 n0_18241_3258 4.828571e+00
R31832 n0_18241_3258 n0_18429_3258 1.074286e+00
R31833 n0_18429_3258 n0_19366_3258 5.354286e+00
R31834 n0_19366_3258 n0_19554_3258 1.074286e+00
R31835 n0_19554_3258 n0_20491_3258 5.354286e+00
R31836 n0_20491_3258 n0_20679_3258 1.074286e+00
R31837 n0_241_3441 n0_429_3441 1.074286e+00
R31838 n0_429_3441 n0_1366_3441 5.354286e+00
R31839 n0_1366_3441 n0_1554_3441 1.074286e+00
R31840 n0_1554_3441 n0_2491_3441 5.354286e+00
R31841 n0_2491_3441 n0_2679_3441 1.074286e+00
R31842 n0_2679_3441 n0_3616_3441 5.354286e+00
R31843 n0_3616_3441 n0_3708_3441 5.257143e-01
R31844 n0_3708_3441 n0_3804_3441 5.485714e-01
R31845 n0_3804_3441 n0_3896_3441 5.257143e-01
R31846 n0_3896_3441 n0_5866_3441 1.125714e+01
R31847 n0_5866_3441 n0_5958_3441 5.257143e-01
R31848 n0_5958_3441 n0_6054_3441 5.485714e-01
R31849 n0_6054_3441 n0_6146_3441 5.257143e-01
R31850 n0_6146_3441 n0_8116_3441 1.125714e+01
R31851 n0_8116_3441 n0_8208_3441 5.257143e-01
R31852 n0_8208_3441 n0_8304_3441 5.485714e-01
R31853 n0_8304_3441 n0_8396_3441 5.257143e-01
R31854 n0_8396_3441 n0_10366_3441 1.125714e+01
R31855 n0_10366_3441 n0_10458_3441 5.257143e-01
R31856 n0_10458_3441 n0_10554_3441 5.485714e-01
R31857 n0_10554_3441 n0_10646_3441 5.257143e-01
R31858 n0_10646_3441 n0_12616_3441 1.125714e+01
R31859 n0_12616_3441 n0_12708_3441 5.257143e-01
R31860 n0_12708_3441 n0_12804_3441 5.485714e-01
R31861 n0_12804_3441 n0_12896_3441 5.257143e-01
R31862 n0_12896_3441 n0_14866_3441 1.125714e+01
R31863 n0_14866_3441 n0_14958_3441 5.257143e-01
R31864 n0_14958_3441 n0_15054_3441 5.485714e-01
R31865 n0_15054_3441 n0_15146_3441 5.257143e-01
R31866 n0_15146_3441 n0_17116_3441 1.125714e+01
R31867 n0_17116_3441 n0_17208_3441 5.257143e-01
R31868 n0_17208_3441 n0_17304_3441 5.485714e-01
R31869 n0_17304_3441 n0_17396_3441 5.257143e-01
R31870 n0_17396_3441 n0_18241_3441 4.828571e+00
R31871 n0_18241_3441 n0_18429_3441 1.074286e+00
R31872 n0_18429_3441 n0_19366_3441 5.354286e+00
R31873 n0_19366_3441 n0_19554_3441 1.074286e+00
R31874 n0_19554_3441 n0_20491_3441 5.354286e+00
R31875 n0_20491_3441 n0_20679_3441 1.074286e+00
R31876 n0_241_3474 n0_429_3474 1.074286e+00
R31877 n0_429_3474 n0_1366_3474 5.354286e+00
R31878 n0_1366_3474 n0_1554_3474 1.074286e+00
R31879 n0_1554_3474 n0_2491_3474 5.354286e+00
R31880 n0_2491_3474 n0_2679_3474 1.074286e+00
R31881 n0_2679_3474 n0_3616_3474 5.354286e+00
R31882 n0_3616_3474 n0_3708_3474 5.257143e-01
R31883 n0_3708_3474 n0_3804_3474 5.485714e-01
R31884 n0_3804_3474 n0_3896_3474 5.257143e-01
R31885 n0_3896_3474 n0_5866_3474 1.125714e+01
R31886 n0_5866_3474 n0_5958_3474 5.257143e-01
R31887 n0_5958_3474 n0_6054_3474 5.485714e-01
R31888 n0_6054_3474 n0_6146_3474 5.257143e-01
R31889 n0_6146_3474 n0_8116_3474 1.125714e+01
R31890 n0_8116_3474 n0_8208_3474 5.257143e-01
R31891 n0_8208_3474 n0_8304_3474 5.485714e-01
R31892 n0_8304_3474 n0_8396_3474 5.257143e-01
R31893 n0_8396_3474 n0_10366_3474 1.125714e+01
R31894 n0_10366_3474 n0_10458_3474 5.257143e-01
R31895 n0_10458_3474 n0_10554_3474 5.485714e-01
R31896 n0_10554_3474 n0_10646_3474 5.257143e-01
R31897 n0_10646_3474 n0_12616_3474 1.125714e+01
R31898 n0_12616_3474 n0_12708_3474 5.257143e-01
R31899 n0_12708_3474 n0_12804_3474 5.485714e-01
R31900 n0_12804_3474 n0_12896_3474 5.257143e-01
R31901 n0_12896_3474 n0_14866_3474 1.125714e+01
R31902 n0_14866_3474 n0_14958_3474 5.257143e-01
R31903 n0_14958_3474 n0_15054_3474 5.485714e-01
R31904 n0_15054_3474 n0_15146_3474 5.257143e-01
R31905 n0_15146_3474 n0_17116_3474 1.125714e+01
R31906 n0_17116_3474 n0_17208_3474 5.257143e-01
R31907 n0_17208_3474 n0_17304_3474 5.485714e-01
R31908 n0_17304_3474 n0_17396_3474 5.257143e-01
R31909 n0_17396_3474 n0_18241_3474 4.828571e+00
R31910 n0_18241_3474 n0_18429_3474 1.074286e+00
R31911 n0_18429_3474 n0_19366_3474 5.354286e+00
R31912 n0_19366_3474 n0_19554_3474 1.074286e+00
R31913 n0_19554_3474 n0_20491_3474 5.354286e+00
R31914 n0_20491_3474 n0_20679_3474 1.074286e+00
R31915 n0_241_3657 n0_429_3657 1.074286e+00
R31916 n0_429_3657 n0_1366_3657 5.354286e+00
R31917 n0_1366_3657 n0_1554_3657 1.074286e+00
R31918 n0_1554_3657 n0_2491_3657 5.354286e+00
R31919 n0_2491_3657 n0_2679_3657 1.074286e+00
R31920 n0_2679_3657 n0_3616_3657 5.354286e+00
R31921 n0_3616_3657 n0_3708_3657 5.257143e-01
R31922 n0_3708_3657 n0_3804_3657 5.485714e-01
R31923 n0_3804_3657 n0_3896_3657 5.257143e-01
R31924 n0_3896_3657 n0_5866_3657 1.125714e+01
R31925 n0_5866_3657 n0_5958_3657 5.257143e-01
R31926 n0_5958_3657 n0_6054_3657 5.485714e-01
R31927 n0_6054_3657 n0_6146_3657 5.257143e-01
R31928 n0_6146_3657 n0_8116_3657 1.125714e+01
R31929 n0_8116_3657 n0_8208_3657 5.257143e-01
R31930 n0_8208_3657 n0_8304_3657 5.485714e-01
R31931 n0_8304_3657 n0_8396_3657 5.257143e-01
R31932 n0_8396_3657 n0_10366_3657 1.125714e+01
R31933 n0_10366_3657 n0_10458_3657 5.257143e-01
R31934 n0_10458_3657 n0_10554_3657 5.485714e-01
R31935 n0_10554_3657 n0_10646_3657 5.257143e-01
R31936 n0_10646_3657 n0_12616_3657 1.125714e+01
R31937 n0_12616_3657 n0_12708_3657 5.257143e-01
R31938 n0_12708_3657 n0_12804_3657 5.485714e-01
R31939 n0_12804_3657 n0_12896_3657 5.257143e-01
R31940 n0_12896_3657 n0_14866_3657 1.125714e+01
R31941 n0_14866_3657 n0_14958_3657 5.257143e-01
R31942 n0_14958_3657 n0_15054_3657 5.485714e-01
R31943 n0_15054_3657 n0_15146_3657 5.257143e-01
R31944 n0_15146_3657 n0_17116_3657 1.125714e+01
R31945 n0_17116_3657 n0_17208_3657 5.257143e-01
R31946 n0_17208_3657 n0_17304_3657 5.485714e-01
R31947 n0_17304_3657 n0_17396_3657 5.257143e-01
R31948 n0_17396_3657 n0_18241_3657 4.828571e+00
R31949 n0_18241_3657 n0_18429_3657 1.074286e+00
R31950 n0_18429_3657 n0_19366_3657 5.354286e+00
R31951 n0_19366_3657 n0_19554_3657 1.074286e+00
R31952 n0_19554_3657 n0_20491_3657 5.354286e+00
R31953 n0_20491_3657 n0_20679_3657 1.074286e+00
R31954 n0_241_3690 n0_429_3690 1.074286e+00
R31955 n0_429_3690 n0_1366_3690 5.354286e+00
R31956 n0_1366_3690 n0_1554_3690 1.074286e+00
R31957 n0_1554_3690 n0_2491_3690 5.354286e+00
R31958 n0_2491_3690 n0_2679_3690 1.074286e+00
R31959 n0_2679_3690 n0_3616_3690 5.354286e+00
R31960 n0_3616_3690 n0_3708_3690 5.257143e-01
R31961 n0_3708_3690 n0_3804_3690 5.485714e-01
R31962 n0_3804_3690 n0_3896_3690 5.257143e-01
R31963 n0_3896_3690 n0_5866_3690 1.125714e+01
R31964 n0_5866_3690 n0_5958_3690 5.257143e-01
R31965 n0_5958_3690 n0_6054_3690 5.485714e-01
R31966 n0_6054_3690 n0_6146_3690 5.257143e-01
R31967 n0_6146_3690 n0_8116_3690 1.125714e+01
R31968 n0_8116_3690 n0_8208_3690 5.257143e-01
R31969 n0_8208_3690 n0_8304_3690 5.485714e-01
R31970 n0_8304_3690 n0_8396_3690 5.257143e-01
R31971 n0_8396_3690 n0_10366_3690 1.125714e+01
R31972 n0_10366_3690 n0_10458_3690 5.257143e-01
R31973 n0_10458_3690 n0_10554_3690 5.485714e-01
R31974 n0_10554_3690 n0_10646_3690 5.257143e-01
R31975 n0_10646_3690 n0_12616_3690 1.125714e+01
R31976 n0_12616_3690 n0_12708_3690 5.257143e-01
R31977 n0_12708_3690 n0_12804_3690 5.485714e-01
R31978 n0_12804_3690 n0_12896_3690 5.257143e-01
R31979 n0_12896_3690 n0_14866_3690 1.125714e+01
R31980 n0_14866_3690 n0_14958_3690 5.257143e-01
R31981 n0_14958_3690 n0_15054_3690 5.485714e-01
R31982 n0_15054_3690 n0_15146_3690 5.257143e-01
R31983 n0_15146_3690 n0_17116_3690 1.125714e+01
R31984 n0_17116_3690 n0_17208_3690 5.257143e-01
R31985 n0_17208_3690 n0_17304_3690 5.485714e-01
R31986 n0_17304_3690 n0_17396_3690 5.257143e-01
R31987 n0_17396_3690 n0_18241_3690 4.828571e+00
R31988 n0_18241_3690 n0_18429_3690 1.074286e+00
R31989 n0_18429_3690 n0_19366_3690 5.354286e+00
R31990 n0_19366_3690 n0_19554_3690 1.074286e+00
R31991 n0_19554_3690 n0_20491_3690 5.354286e+00
R31992 n0_20491_3690 n0_20679_3690 1.074286e+00
R31993 n0_241_3873 n0_380_3873 7.942857e-01
R31994 n0_380_3873 n0_429_3873 2.800000e-01
R31995 n0_429_3873 n0_1366_3873 5.354286e+00
R31996 n0_1366_3873 n0_1505_3873 7.942857e-01
R31997 n0_1505_3873 n0_1554_3873 2.800000e-01
R31998 n0_1554_3873 n0_2491_3873 5.354286e+00
R31999 n0_2491_3873 n0_2630_3873 7.942857e-01
R32000 n0_2630_3873 n0_2679_3873 2.800000e-01
R32001 n0_2679_3873 n0_3616_3873 5.354286e+00
R32002 n0_3616_3873 n0_3708_3873 5.257143e-01
R32003 n0_3708_3873 n0_3755_3873 2.685714e-01
R32004 n0_3755_3873 n0_3804_3873 2.800000e-01
R32005 n0_3804_3873 n0_5866_3873 1.178286e+01
R32006 n0_5866_3873 n0_5958_3873 5.257143e-01
R32007 n0_5958_3873 n0_6005_3873 2.685714e-01
R32008 n0_6005_3873 n0_6054_3873 2.800000e-01
R32009 n0_6054_3873 n0_6146_3873 5.257143e-01
R32010 n0_6146_3873 n0_8116_3873 1.125714e+01
R32011 n0_8116_3873 n0_8208_3873 5.257143e-01
R32012 n0_8208_3873 n0_8255_3873 2.685714e-01
R32013 n0_8255_3873 n0_8304_3873 2.800000e-01
R32014 n0_8304_3873 n0_8396_3873 5.257143e-01
R32015 n0_8396_3873 n0_10366_3873 1.125714e+01
R32016 n0_10366_3873 n0_10458_3873 5.257143e-01
R32017 n0_10458_3873 n0_10505_3873 2.685714e-01
R32018 n0_10505_3873 n0_10554_3873 2.800000e-01
R32019 n0_10554_3873 n0_10646_3873 5.257143e-01
R32020 n0_10646_3873 n0_12616_3873 1.125714e+01
R32021 n0_12616_3873 n0_12708_3873 5.257143e-01
R32022 n0_12708_3873 n0_12755_3873 2.685714e-01
R32023 n0_12755_3873 n0_12804_3873 2.800000e-01
R32024 n0_12804_3873 n0_12896_3873 5.257143e-01
R32025 n0_12896_3873 n0_14866_3873 1.125714e+01
R32026 n0_14866_3873 n0_14958_3873 5.257143e-01
R32027 n0_14958_3873 n0_15005_3873 2.685714e-01
R32028 n0_15005_3873 n0_15054_3873 2.800000e-01
R32029 n0_15054_3873 n0_15146_3873 5.257143e-01
R32030 n0_15146_3873 n0_17116_3873 1.125714e+01
R32031 n0_17116_3873 n0_17208_3873 5.257143e-01
R32032 n0_17208_3873 n0_17255_3873 2.685714e-01
R32033 n0_17255_3873 n0_17304_3873 2.800000e-01
R32034 n0_17304_3873 n0_18241_3873 5.354286e+00
R32035 n0_18241_3873 n0_18380_3873 7.942857e-01
R32036 n0_18380_3873 n0_18429_3873 2.800000e-01
R32037 n0_18429_3873 n0_19366_3873 5.354286e+00
R32038 n0_19366_3873 n0_19505_3873 7.942857e-01
R32039 n0_19505_3873 n0_19554_3873 2.800000e-01
R32040 n0_19554_3873 n0_20491_3873 5.354286e+00
R32041 n0_20491_3873 n0_20630_3873 7.942857e-01
R32042 n0_20630_3873 n0_20679_3873 2.800000e-01
R32043 n0_241_3906 n0_380_3906 7.942857e-01
R32044 n0_380_3906 n0_429_3906 2.800000e-01
R32045 n0_429_3906 n0_1366_3906 5.354286e+00
R32046 n0_1366_3906 n0_1505_3906 7.942857e-01
R32047 n0_1505_3906 n0_1554_3906 2.800000e-01
R32048 n0_1554_3906 n0_2491_3906 5.354286e+00
R32049 n0_2491_3906 n0_2630_3906 7.942857e-01
R32050 n0_2630_3906 n0_2679_3906 2.800000e-01
R32051 n0_2679_3906 n0_3616_3906 5.354286e+00
R32052 n0_3616_3906 n0_3708_3906 5.257143e-01
R32053 n0_3708_3906 n0_3755_3906 2.685714e-01
R32054 n0_3755_3906 n0_3804_3906 2.800000e-01
R32055 n0_3804_3906 n0_5866_3906 1.178286e+01
R32056 n0_5866_3906 n0_5958_3906 5.257143e-01
R32057 n0_5958_3906 n0_6005_3906 2.685714e-01
R32058 n0_6005_3906 n0_6054_3906 2.800000e-01
R32059 n0_6054_3906 n0_6146_3906 5.257143e-01
R32060 n0_6146_3906 n0_8116_3906 1.125714e+01
R32061 n0_8116_3906 n0_8208_3906 5.257143e-01
R32062 n0_8208_3906 n0_8255_3906 2.685714e-01
R32063 n0_8255_3906 n0_8304_3906 2.800000e-01
R32064 n0_8304_3906 n0_8396_3906 5.257143e-01
R32065 n0_8396_3906 n0_10366_3906 1.125714e+01
R32066 n0_10366_3906 n0_10458_3906 5.257143e-01
R32067 n0_10458_3906 n0_10505_3906 2.685714e-01
R32068 n0_10505_3906 n0_10554_3906 2.800000e-01
R32069 n0_10554_3906 n0_10646_3906 5.257143e-01
R32070 n0_10646_3906 n0_12616_3906 1.125714e+01
R32071 n0_12616_3906 n0_12708_3906 5.257143e-01
R32072 n0_12708_3906 n0_12755_3906 2.685714e-01
R32073 n0_12755_3906 n0_12804_3906 2.800000e-01
R32074 n0_12804_3906 n0_12896_3906 5.257143e-01
R32075 n0_12896_3906 n0_14866_3906 1.125714e+01
R32076 n0_14866_3906 n0_14958_3906 5.257143e-01
R32077 n0_14958_3906 n0_15005_3906 2.685714e-01
R32078 n0_15005_3906 n0_15054_3906 2.800000e-01
R32079 n0_15054_3906 n0_15146_3906 5.257143e-01
R32080 n0_15146_3906 n0_17116_3906 1.125714e+01
R32081 n0_17116_3906 n0_17208_3906 5.257143e-01
R32082 n0_17208_3906 n0_17255_3906 2.685714e-01
R32083 n0_17255_3906 n0_17304_3906 2.800000e-01
R32084 n0_17304_3906 n0_18241_3906 5.354286e+00
R32085 n0_18241_3906 n0_18380_3906 7.942857e-01
R32086 n0_18380_3906 n0_18429_3906 2.800000e-01
R32087 n0_18429_3906 n0_19366_3906 5.354286e+00
R32088 n0_19366_3906 n0_19505_3906 7.942857e-01
R32089 n0_19505_3906 n0_19554_3906 2.800000e-01
R32090 n0_19554_3906 n0_20491_3906 5.354286e+00
R32091 n0_20491_3906 n0_20630_3906 7.942857e-01
R32092 n0_20630_3906 n0_20679_3906 2.800000e-01
R32093 n0_241_4089 n0_429_4089 1.074286e+00
R32094 n0_429_4089 n0_1366_4089 5.354286e+00
R32095 n0_1366_4089 n0_1554_4089 1.074286e+00
R32096 n0_1554_4089 n0_2491_4089 5.354286e+00
R32097 n0_2491_4089 n0_2679_4089 1.074286e+00
R32098 n0_2679_4089 n0_3616_4089 5.354286e+00
R32099 n0_3616_4089 n0_3804_4089 1.074286e+00
R32100 n0_3804_4089 n0_5866_4089 1.178286e+01
R32101 n0_5866_4089 n0_5958_4089 5.257143e-01
R32102 n0_5958_4089 n0_6054_4089 5.485714e-01
R32103 n0_6054_4089 n0_6146_4089 5.257143e-01
R32104 n0_6146_4089 n0_8116_4089 1.125714e+01
R32105 n0_8116_4089 n0_8208_4089 5.257143e-01
R32106 n0_8208_4089 n0_8304_4089 5.485714e-01
R32107 n0_8304_4089 n0_8396_4089 5.257143e-01
R32108 n0_8396_4089 n0_10366_4089 1.125714e+01
R32109 n0_10366_4089 n0_10458_4089 5.257143e-01
R32110 n0_10458_4089 n0_10554_4089 5.485714e-01
R32111 n0_10554_4089 n0_10646_4089 5.257143e-01
R32112 n0_10646_4089 n0_12616_4089 1.125714e+01
R32113 n0_12616_4089 n0_12708_4089 5.257143e-01
R32114 n0_12708_4089 n0_12804_4089 5.485714e-01
R32115 n0_12804_4089 n0_12896_4089 5.257143e-01
R32116 n0_12896_4089 n0_14866_4089 1.125714e+01
R32117 n0_14866_4089 n0_14958_4089 5.257143e-01
R32118 n0_14958_4089 n0_15054_4089 5.485714e-01
R32119 n0_15054_4089 n0_15146_4089 5.257143e-01
R32120 n0_15146_4089 n0_17116_4089 1.125714e+01
R32121 n0_17116_4089 n0_17304_4089 1.074286e+00
R32122 n0_17304_4089 n0_18241_4089 5.354286e+00
R32123 n0_18241_4089 n0_18429_4089 1.074286e+00
R32124 n0_18429_4089 n0_19366_4089 5.354286e+00
R32125 n0_19366_4089 n0_19554_4089 1.074286e+00
R32126 n0_19554_4089 n0_20491_4089 5.354286e+00
R32127 n0_20491_4089 n0_20679_4089 1.074286e+00
R32128 n0_241_4122 n0_429_4122 1.074286e+00
R32129 n0_429_4122 n0_1366_4122 5.354286e+00
R32130 n0_1366_4122 n0_1554_4122 1.074286e+00
R32131 n0_1554_4122 n0_2491_4122 5.354286e+00
R32132 n0_2491_4122 n0_2679_4122 1.074286e+00
R32133 n0_2679_4122 n0_3616_4122 5.354286e+00
R32134 n0_3616_4122 n0_3804_4122 1.074286e+00
R32135 n0_3804_4122 n0_5866_4122 1.178286e+01
R32136 n0_5866_4122 n0_5958_4122 5.257143e-01
R32137 n0_5958_4122 n0_6054_4122 5.485714e-01
R32138 n0_6054_4122 n0_6146_4122 5.257143e-01
R32139 n0_6146_4122 n0_8116_4122 1.125714e+01
R32140 n0_8116_4122 n0_8208_4122 5.257143e-01
R32141 n0_8208_4122 n0_8304_4122 5.485714e-01
R32142 n0_8304_4122 n0_8396_4122 5.257143e-01
R32143 n0_8396_4122 n0_10366_4122 1.125714e+01
R32144 n0_10366_4122 n0_10458_4122 5.257143e-01
R32145 n0_10458_4122 n0_10554_4122 5.485714e-01
R32146 n0_10554_4122 n0_10646_4122 5.257143e-01
R32147 n0_10646_4122 n0_12616_4122 1.125714e+01
R32148 n0_12616_4122 n0_12708_4122 5.257143e-01
R32149 n0_12708_4122 n0_12804_4122 5.485714e-01
R32150 n0_12804_4122 n0_12896_4122 5.257143e-01
R32151 n0_12896_4122 n0_14866_4122 1.125714e+01
R32152 n0_14866_4122 n0_14958_4122 5.257143e-01
R32153 n0_14958_4122 n0_15054_4122 5.485714e-01
R32154 n0_15054_4122 n0_15146_4122 5.257143e-01
R32155 n0_15146_4122 n0_17116_4122 1.125714e+01
R32156 n0_17116_4122 n0_17304_4122 1.074286e+00
R32157 n0_17304_4122 n0_18241_4122 5.354286e+00
R32158 n0_18241_4122 n0_18429_4122 1.074286e+00
R32159 n0_18429_4122 n0_19366_4122 5.354286e+00
R32160 n0_19366_4122 n0_19554_4122 1.074286e+00
R32161 n0_19554_4122 n0_20491_4122 5.354286e+00
R32162 n0_20491_4122 n0_20679_4122 1.074286e+00
R32163 n0_241_4305 n0_429_4305 1.074286e+00
R32164 n0_429_4305 n0_1366_4305 5.354286e+00
R32165 n0_1366_4305 n0_1554_4305 1.074286e+00
R32166 n0_1554_4305 n0_2491_4305 5.354286e+00
R32167 n0_2491_4305 n0_2679_4305 1.074286e+00
R32168 n0_2679_4305 n0_3616_4305 5.354286e+00
R32169 n0_3616_4305 n0_3804_4305 1.074286e+00
R32170 n0_3804_4305 n0_5866_4305 1.178286e+01
R32171 n0_5866_4305 n0_5958_4305 5.257143e-01
R32172 n0_5958_4305 n0_6054_4305 5.485714e-01
R32173 n0_6054_4305 n0_6146_4305 5.257143e-01
R32174 n0_6146_4305 n0_8116_4305 1.125714e+01
R32175 n0_8116_4305 n0_8208_4305 5.257143e-01
R32176 n0_8208_4305 n0_8304_4305 5.485714e-01
R32177 n0_8304_4305 n0_8396_4305 5.257143e-01
R32178 n0_8396_4305 n0_10366_4305 1.125714e+01
R32179 n0_10366_4305 n0_10458_4305 5.257143e-01
R32180 n0_10458_4305 n0_10554_4305 5.485714e-01
R32181 n0_10554_4305 n0_10646_4305 5.257143e-01
R32182 n0_10646_4305 n0_12616_4305 1.125714e+01
R32183 n0_12616_4305 n0_12708_4305 5.257143e-01
R32184 n0_12708_4305 n0_12804_4305 5.485714e-01
R32185 n0_12804_4305 n0_12896_4305 5.257143e-01
R32186 n0_12896_4305 n0_14866_4305 1.125714e+01
R32187 n0_14866_4305 n0_14958_4305 5.257143e-01
R32188 n0_14958_4305 n0_15054_4305 5.485714e-01
R32189 n0_15054_4305 n0_15146_4305 5.257143e-01
R32190 n0_15146_4305 n0_17116_4305 1.125714e+01
R32191 n0_17116_4305 n0_17304_4305 1.074286e+00
R32192 n0_17304_4305 n0_18241_4305 5.354286e+00
R32193 n0_18241_4305 n0_18429_4305 1.074286e+00
R32194 n0_18429_4305 n0_19366_4305 5.354286e+00
R32195 n0_19366_4305 n0_19554_4305 1.074286e+00
R32196 n0_19554_4305 n0_20491_4305 5.354286e+00
R32197 n0_20491_4305 n0_20679_4305 1.074286e+00
R32198 n0_241_4338 n0_429_4338 1.074286e+00
R32199 n0_429_4338 n0_1366_4338 5.354286e+00
R32200 n0_1366_4338 n0_1554_4338 1.074286e+00
R32201 n0_1554_4338 n0_2491_4338 5.354286e+00
R32202 n0_2491_4338 n0_2679_4338 1.074286e+00
R32203 n0_2679_4338 n0_3616_4338 5.354286e+00
R32204 n0_3616_4338 n0_3804_4338 1.074286e+00
R32205 n0_3804_4338 n0_5866_4338 1.178286e+01
R32206 n0_5866_4338 n0_5958_4338 5.257143e-01
R32207 n0_5958_4338 n0_6054_4338 5.485714e-01
R32208 n0_6054_4338 n0_6146_4338 5.257143e-01
R32209 n0_6146_4338 n0_8116_4338 1.125714e+01
R32210 n0_8116_4338 n0_8208_4338 5.257143e-01
R32211 n0_8208_4338 n0_8304_4338 5.485714e-01
R32212 n0_8304_4338 n0_8396_4338 5.257143e-01
R32213 n0_8396_4338 n0_10366_4338 1.125714e+01
R32214 n0_10366_4338 n0_10458_4338 5.257143e-01
R32215 n0_10458_4338 n0_10554_4338 5.485714e-01
R32216 n0_10554_4338 n0_10646_4338 5.257143e-01
R32217 n0_10646_4338 n0_12616_4338 1.125714e+01
R32218 n0_12616_4338 n0_12708_4338 5.257143e-01
R32219 n0_12708_4338 n0_12804_4338 5.485714e-01
R32220 n0_12804_4338 n0_12896_4338 5.257143e-01
R32221 n0_12896_4338 n0_14866_4338 1.125714e+01
R32222 n0_14866_4338 n0_14958_4338 5.257143e-01
R32223 n0_14958_4338 n0_15054_4338 5.485714e-01
R32224 n0_15054_4338 n0_15146_4338 5.257143e-01
R32225 n0_15146_4338 n0_17116_4338 1.125714e+01
R32226 n0_17116_4338 n0_17304_4338 1.074286e+00
R32227 n0_17304_4338 n0_18241_4338 5.354286e+00
R32228 n0_18241_4338 n0_18429_4338 1.074286e+00
R32229 n0_18429_4338 n0_19366_4338 5.354286e+00
R32230 n0_19366_4338 n0_19554_4338 1.074286e+00
R32231 n0_19554_4338 n0_20491_4338 5.354286e+00
R32232 n0_20491_4338 n0_20679_4338 1.074286e+00
R32233 n0_241_4521 n0_429_4521 1.074286e+00
R32234 n0_429_4521 n0_1366_4521 5.354286e+00
R32235 n0_1366_4521 n0_1554_4521 1.074286e+00
R32236 n0_1554_4521 n0_2491_4521 5.354286e+00
R32237 n0_2491_4521 n0_2679_4521 1.074286e+00
R32238 n0_2679_4521 n0_3616_4521 5.354286e+00
R32239 n0_3616_4521 n0_3804_4521 1.074286e+00
R32240 n0_3804_4521 n0_5866_4521 1.178286e+01
R32241 n0_5866_4521 n0_5958_4521 5.257143e-01
R32242 n0_5958_4521 n0_6054_4521 5.485714e-01
R32243 n0_6054_4521 n0_6146_4521 5.257143e-01
R32244 n0_6146_4521 n0_8116_4521 1.125714e+01
R32245 n0_8116_4521 n0_8208_4521 5.257143e-01
R32246 n0_8208_4521 n0_8304_4521 5.485714e-01
R32247 n0_8304_4521 n0_8396_4521 5.257143e-01
R32248 n0_8396_4521 n0_10366_4521 1.125714e+01
R32249 n0_10366_4521 n0_10458_4521 5.257143e-01
R32250 n0_10458_4521 n0_10554_4521 5.485714e-01
R32251 n0_10554_4521 n0_10646_4521 5.257143e-01
R32252 n0_10646_4521 n0_12616_4521 1.125714e+01
R32253 n0_12616_4521 n0_12708_4521 5.257143e-01
R32254 n0_12708_4521 n0_12804_4521 5.485714e-01
R32255 n0_12804_4521 n0_12896_4521 5.257143e-01
R32256 n0_12896_4521 n0_14866_4521 1.125714e+01
R32257 n0_14866_4521 n0_14958_4521 5.257143e-01
R32258 n0_14958_4521 n0_15054_4521 5.485714e-01
R32259 n0_15054_4521 n0_15146_4521 5.257143e-01
R32260 n0_15146_4521 n0_17116_4521 1.125714e+01
R32261 n0_17116_4521 n0_17304_4521 1.074286e+00
R32262 n0_17304_4521 n0_18241_4521 5.354286e+00
R32263 n0_18241_4521 n0_18429_4521 1.074286e+00
R32264 n0_18429_4521 n0_19366_4521 5.354286e+00
R32265 n0_19366_4521 n0_19554_4521 1.074286e+00
R32266 n0_19554_4521 n0_20491_4521 5.354286e+00
R32267 n0_20491_4521 n0_20679_4521 1.074286e+00
R32268 n0_241_4554 n0_429_4554 1.074286e+00
R32269 n0_429_4554 n0_1366_4554 5.354286e+00
R32270 n0_1366_4554 n0_1554_4554 1.074286e+00
R32271 n0_1554_4554 n0_2491_4554 5.354286e+00
R32272 n0_2491_4554 n0_2679_4554 1.074286e+00
R32273 n0_2679_4554 n0_3616_4554 5.354286e+00
R32274 n0_3616_4554 n0_3804_4554 1.074286e+00
R32275 n0_3804_4554 n0_5866_4554 1.178286e+01
R32276 n0_5866_4554 n0_5958_4554 5.257143e-01
R32277 n0_5958_4554 n0_6054_4554 5.485714e-01
R32278 n0_6054_4554 n0_6146_4554 5.257143e-01
R32279 n0_6146_4554 n0_8116_4554 1.125714e+01
R32280 n0_8116_4554 n0_8208_4554 5.257143e-01
R32281 n0_8208_4554 n0_8304_4554 5.485714e-01
R32282 n0_8304_4554 n0_8396_4554 5.257143e-01
R32283 n0_8396_4554 n0_10366_4554 1.125714e+01
R32284 n0_10366_4554 n0_10458_4554 5.257143e-01
R32285 n0_10458_4554 n0_10554_4554 5.485714e-01
R32286 n0_10554_4554 n0_10646_4554 5.257143e-01
R32287 n0_10646_4554 n0_12616_4554 1.125714e+01
R32288 n0_12616_4554 n0_12708_4554 5.257143e-01
R32289 n0_12708_4554 n0_12804_4554 5.485714e-01
R32290 n0_12804_4554 n0_12896_4554 5.257143e-01
R32291 n0_12896_4554 n0_14866_4554 1.125714e+01
R32292 n0_14866_4554 n0_14958_4554 5.257143e-01
R32293 n0_14958_4554 n0_15054_4554 5.485714e-01
R32294 n0_15054_4554 n0_15146_4554 5.257143e-01
R32295 n0_15146_4554 n0_17116_4554 1.125714e+01
R32296 n0_17116_4554 n0_17304_4554 1.074286e+00
R32297 n0_17304_4554 n0_18241_4554 5.354286e+00
R32298 n0_18241_4554 n0_18429_4554 1.074286e+00
R32299 n0_18429_4554 n0_19366_4554 5.354286e+00
R32300 n0_19366_4554 n0_19554_4554 1.074286e+00
R32301 n0_19554_4554 n0_20491_4554 5.354286e+00
R32302 n0_20491_4554 n0_20679_4554 1.074286e+00
R32303 n0_241_4737 n0_429_4737 1.074286e+00
R32304 n0_429_4737 n0_1366_4737 5.354286e+00
R32305 n0_1366_4737 n0_1554_4737 1.074286e+00
R32306 n0_1554_4737 n0_2491_4737 5.354286e+00
R32307 n0_2491_4737 n0_2679_4737 1.074286e+00
R32308 n0_2679_4737 n0_3616_4737 5.354286e+00
R32309 n0_3616_4737 n0_3804_4737 1.074286e+00
R32310 n0_3804_4737 n0_5866_4737 1.178286e+01
R32311 n0_5866_4737 n0_5958_4737 5.257143e-01
R32312 n0_5958_4737 n0_6054_4737 5.485714e-01
R32313 n0_6054_4737 n0_6146_4737 5.257143e-01
R32314 n0_6146_4737 n0_8116_4737 1.125714e+01
R32315 n0_8116_4737 n0_8208_4737 5.257143e-01
R32316 n0_8208_4737 n0_8304_4737 5.485714e-01
R32317 n0_8304_4737 n0_8396_4737 5.257143e-01
R32318 n0_8396_4737 n0_10366_4737 1.125714e+01
R32319 n0_10366_4737 n0_10458_4737 5.257143e-01
R32320 n0_10458_4737 n0_10554_4737 5.485714e-01
R32321 n0_10554_4737 n0_10646_4737 5.257143e-01
R32322 n0_10646_4737 n0_12616_4737 1.125714e+01
R32323 n0_12616_4737 n0_12708_4737 5.257143e-01
R32324 n0_12708_4737 n0_12804_4737 5.485714e-01
R32325 n0_12804_4737 n0_12896_4737 5.257143e-01
R32326 n0_12896_4737 n0_14866_4737 1.125714e+01
R32327 n0_14866_4737 n0_14958_4737 5.257143e-01
R32328 n0_14958_4737 n0_15054_4737 5.485714e-01
R32329 n0_15054_4737 n0_15146_4737 5.257143e-01
R32330 n0_15146_4737 n0_17116_4737 1.125714e+01
R32331 n0_17116_4737 n0_17304_4737 1.074286e+00
R32332 n0_17304_4737 n0_18241_4737 5.354286e+00
R32333 n0_18241_4737 n0_18429_4737 1.074286e+00
R32334 n0_18429_4737 n0_19366_4737 5.354286e+00
R32335 n0_19366_4737 n0_19554_4737 1.074286e+00
R32336 n0_19554_4737 n0_20491_4737 5.354286e+00
R32337 n0_20491_4737 n0_20679_4737 1.074286e+00
R32338 n0_241_4770 n0_429_4770 1.074286e+00
R32339 n0_429_4770 n0_1366_4770 5.354286e+00
R32340 n0_1366_4770 n0_1554_4770 1.074286e+00
R32341 n0_1554_4770 n0_2491_4770 5.354286e+00
R32342 n0_2491_4770 n0_2679_4770 1.074286e+00
R32343 n0_2679_4770 n0_3616_4770 5.354286e+00
R32344 n0_3616_4770 n0_3804_4770 1.074286e+00
R32345 n0_3804_4770 n0_5866_4770 1.178286e+01
R32346 n0_5866_4770 n0_5958_4770 5.257143e-01
R32347 n0_5958_4770 n0_6054_4770 5.485714e-01
R32348 n0_6054_4770 n0_6146_4770 5.257143e-01
R32349 n0_6146_4770 n0_8116_4770 1.125714e+01
R32350 n0_8116_4770 n0_8208_4770 5.257143e-01
R32351 n0_8208_4770 n0_8304_4770 5.485714e-01
R32352 n0_8304_4770 n0_8396_4770 5.257143e-01
R32353 n0_8396_4770 n0_10366_4770 1.125714e+01
R32354 n0_10366_4770 n0_10458_4770 5.257143e-01
R32355 n0_10458_4770 n0_10554_4770 5.485714e-01
R32356 n0_10554_4770 n0_10646_4770 5.257143e-01
R32357 n0_10646_4770 n0_12616_4770 1.125714e+01
R32358 n0_12616_4770 n0_12708_4770 5.257143e-01
R32359 n0_12708_4770 n0_12804_4770 5.485714e-01
R32360 n0_12804_4770 n0_12896_4770 5.257143e-01
R32361 n0_12896_4770 n0_14866_4770 1.125714e+01
R32362 n0_14866_4770 n0_14958_4770 5.257143e-01
R32363 n0_14958_4770 n0_15054_4770 5.485714e-01
R32364 n0_15054_4770 n0_15146_4770 5.257143e-01
R32365 n0_15146_4770 n0_17116_4770 1.125714e+01
R32366 n0_17116_4770 n0_17304_4770 1.074286e+00
R32367 n0_17304_4770 n0_18241_4770 5.354286e+00
R32368 n0_18241_4770 n0_18429_4770 1.074286e+00
R32369 n0_18429_4770 n0_19366_4770 5.354286e+00
R32370 n0_19366_4770 n0_19554_4770 1.074286e+00
R32371 n0_19554_4770 n0_20491_4770 5.354286e+00
R32372 n0_20491_4770 n0_20679_4770 1.074286e+00
R32373 n0_241_4953 n0_1366_4953 6.428571e+00
R32374 n0_1366_4953 n0_2491_4953 6.428571e+00
R32375 n0_2491_4953 n0_3616_4953 6.428571e+00
R32376 n0_3616_4953 n0_5866_4953 1.285714e+01
R32377 n0_5866_4953 n0_5958_4953 5.257143e-01
R32378 n0_5958_4953 n0_6005_4953 2.685714e-01
R32379 n0_6005_4953 n0_6054_4953 2.800000e-01
R32380 n0_6054_4953 n0_6146_4953 5.257143e-01
R32381 n0_6146_4953 n0_8116_4953 1.125714e+01
R32382 n0_8116_4953 n0_8208_4953 5.257143e-01
R32383 n0_8208_4953 n0_8255_4953 2.685714e-01
R32384 n0_8255_4953 n0_8304_4953 2.800000e-01
R32385 n0_8304_4953 n0_8396_4953 5.257143e-01
R32386 n0_8396_4953 n0_10366_4953 1.125714e+01
R32387 n0_10366_4953 n0_10458_4953 5.257143e-01
R32388 n0_10458_4953 n0_10505_4953 2.685714e-01
R32389 n0_10505_4953 n0_10554_4953 2.800000e-01
R32390 n0_10554_4953 n0_10646_4953 5.257143e-01
R32391 n0_10646_4953 n0_12616_4953 1.125714e+01
R32392 n0_12616_4953 n0_12708_4953 5.257143e-01
R32393 n0_12708_4953 n0_12755_4953 2.685714e-01
R32394 n0_12755_4953 n0_12804_4953 2.800000e-01
R32395 n0_12804_4953 n0_12896_4953 5.257143e-01
R32396 n0_12896_4953 n0_14866_4953 1.125714e+01
R32397 n0_14866_4953 n0_14958_4953 5.257143e-01
R32398 n0_14958_4953 n0_15005_4953 2.685714e-01
R32399 n0_15005_4953 n0_15054_4953 2.800000e-01
R32400 n0_15054_4953 n0_15146_4953 5.257143e-01
R32401 n0_15146_4953 n0_17116_4953 1.125714e+01
R32402 n0_17116_4953 n0_18241_4953 6.428571e+00
R32403 n0_18241_4953 n0_19366_4953 6.428571e+00
R32404 n0_19366_4953 n0_20491_4953 6.428571e+00
R32405 n0_241_4986 n0_1366_4986 6.428571e+00
R32406 n0_1366_4986 n0_2491_4986 6.428571e+00
R32407 n0_2491_4986 n0_3616_4986 6.428571e+00
R32408 n0_3616_4986 n0_5958_4986 1.338286e+01
R32409 n0_5958_4986 n0_6005_4986 2.685714e-01
R32410 n0_6005_4986 n0_6054_4986 2.800000e-01
R32411 n0_6054_4986 n0_8208_4986 1.230857e+01
R32412 n0_8208_4986 n0_8255_4986 2.685714e-01
R32413 n0_8255_4986 n0_8304_4986 2.800000e-01
R32414 n0_8304_4986 n0_10458_4986 1.230857e+01
R32415 n0_10458_4986 n0_10505_4986 2.685714e-01
R32416 n0_10505_4986 n0_10554_4986 2.800000e-01
R32417 n0_10554_4986 n0_12708_4986 1.230857e+01
R32418 n0_12708_4986 n0_12755_4986 2.685714e-01
R32419 n0_12755_4986 n0_12804_4986 2.800000e-01
R32420 n0_12804_4986 n0_14958_4986 1.230857e+01
R32421 n0_14958_4986 n0_15005_4986 2.685714e-01
R32422 n0_15005_4986 n0_15054_4986 2.800000e-01
R32423 n0_15054_4986 n0_17116_4986 1.178286e+01
R32424 n0_17116_4986 n0_18241_4986 6.428571e+00
R32425 n0_18241_4986 n0_19366_4986 6.428571e+00
R32426 n0_19366_4986 n0_20491_4986 6.428571e+00
R32427 n0_241_5169 n0_429_5169 1.074286e+00
R32428 n0_429_5169 n0_1366_5169 5.354286e+00
R32429 n0_1366_5169 n0_1554_5169 1.074286e+00
R32430 n0_1554_5169 n0_2491_5169 5.354286e+00
R32431 n0_2491_5169 n0_2679_5169 1.074286e+00
R32432 n0_2679_5169 n0_3616_5169 5.354286e+00
R32433 n0_3616_5169 n0_3804_5169 1.074286e+00
R32434 n0_3804_5169 n0_4741_5169 5.354286e+00
R32435 n0_4741_5169 n0_4929_5169 1.074286e+00
R32436 n0_4929_5169 n0_5866_5169 5.354286e+00
R32437 n0_5866_5169 n0_5958_5169 5.257143e-01
R32438 n0_5958_5169 n0_6054_5169 5.485714e-01
R32439 n0_6054_5169 n0_6146_5169 5.257143e-01
R32440 n0_6146_5169 n0_8116_5169 1.125714e+01
R32441 n0_8116_5169 n0_8208_5169 5.257143e-01
R32442 n0_8208_5169 n0_8304_5169 5.485714e-01
R32443 n0_8304_5169 n0_8396_5169 5.257143e-01
R32444 n0_8396_5169 n0_10366_5169 1.125714e+01
R32445 n0_10366_5169 n0_10458_5169 5.257143e-01
R32446 n0_10458_5169 n0_10554_5169 5.485714e-01
R32447 n0_10554_5169 n0_10646_5169 5.257143e-01
R32448 n0_10646_5169 n0_12616_5169 1.125714e+01
R32449 n0_12616_5169 n0_12708_5169 5.257143e-01
R32450 n0_12708_5169 n0_12804_5169 5.485714e-01
R32451 n0_12804_5169 n0_12896_5169 5.257143e-01
R32452 n0_12896_5169 n0_14866_5169 1.125714e+01
R32453 n0_14866_5169 n0_14958_5169 5.257143e-01
R32454 n0_14958_5169 n0_15054_5169 5.485714e-01
R32455 n0_15054_5169 n0_15146_5169 5.257143e-01
R32456 n0_15146_5169 n0_15991_5169 4.828571e+00
R32457 n0_15991_5169 n0_16179_5169 1.074286e+00
R32458 n0_16179_5169 n0_17116_5169 5.354286e+00
R32459 n0_17116_5169 n0_17304_5169 1.074286e+00
R32460 n0_17304_5169 n0_18241_5169 5.354286e+00
R32461 n0_18241_5169 n0_18429_5169 1.074286e+00
R32462 n0_18429_5169 n0_19366_5169 5.354286e+00
R32463 n0_19366_5169 n0_19554_5169 1.074286e+00
R32464 n0_19554_5169 n0_20491_5169 5.354286e+00
R32465 n0_20491_5169 n0_20679_5169 1.074286e+00
R32466 n0_241_5202 n0_429_5202 1.074286e+00
R32467 n0_429_5202 n0_1366_5202 5.354286e+00
R32468 n0_1366_5202 n0_1554_5202 1.074286e+00
R32469 n0_1554_5202 n0_2491_5202 5.354286e+00
R32470 n0_2491_5202 n0_2679_5202 1.074286e+00
R32471 n0_2679_5202 n0_3616_5202 5.354286e+00
R32472 n0_3616_5202 n0_3804_5202 1.074286e+00
R32473 n0_3804_5202 n0_4741_5202 5.354286e+00
R32474 n0_4741_5202 n0_4929_5202 1.074286e+00
R32475 n0_4929_5202 n0_5866_5202 5.354286e+00
R32476 n0_5866_5202 n0_5958_5202 5.257143e-01
R32477 n0_5958_5202 n0_6054_5202 5.485714e-01
R32478 n0_6054_5202 n0_6146_5202 5.257143e-01
R32479 n0_6146_5202 n0_8116_5202 1.125714e+01
R32480 n0_8116_5202 n0_8208_5202 5.257143e-01
R32481 n0_8208_5202 n0_8304_5202 5.485714e-01
R32482 n0_8304_5202 n0_8396_5202 5.257143e-01
R32483 n0_8396_5202 n0_10366_5202 1.125714e+01
R32484 n0_10366_5202 n0_10458_5202 5.257143e-01
R32485 n0_10458_5202 n0_10554_5202 5.485714e-01
R32486 n0_10554_5202 n0_10646_5202 5.257143e-01
R32487 n0_10646_5202 n0_12616_5202 1.125714e+01
R32488 n0_12616_5202 n0_12708_5202 5.257143e-01
R32489 n0_12708_5202 n0_12804_5202 5.485714e-01
R32490 n0_12804_5202 n0_12896_5202 5.257143e-01
R32491 n0_12896_5202 n0_14866_5202 1.125714e+01
R32492 n0_14866_5202 n0_14958_5202 5.257143e-01
R32493 n0_14958_5202 n0_15054_5202 5.485714e-01
R32494 n0_15054_5202 n0_15146_5202 5.257143e-01
R32495 n0_15146_5202 n0_15991_5202 4.828571e+00
R32496 n0_15991_5202 n0_16179_5202 1.074286e+00
R32497 n0_16179_5202 n0_17116_5202 5.354286e+00
R32498 n0_17116_5202 n0_17304_5202 1.074286e+00
R32499 n0_17304_5202 n0_18241_5202 5.354286e+00
R32500 n0_18241_5202 n0_18429_5202 1.074286e+00
R32501 n0_18429_5202 n0_19366_5202 5.354286e+00
R32502 n0_19366_5202 n0_19554_5202 1.074286e+00
R32503 n0_19554_5202 n0_20491_5202 5.354286e+00
R32504 n0_20491_5202 n0_20679_5202 1.074286e+00
R32505 n0_241_5385 n0_429_5385 1.074286e+00
R32506 n0_429_5385 n0_1366_5385 5.354286e+00
R32507 n0_1366_5385 n0_1554_5385 1.074286e+00
R32508 n0_1554_5385 n0_2491_5385 5.354286e+00
R32509 n0_2491_5385 n0_2679_5385 1.074286e+00
R32510 n0_2679_5385 n0_3616_5385 5.354286e+00
R32511 n0_3616_5385 n0_3804_5385 1.074286e+00
R32512 n0_3804_5385 n0_4741_5385 5.354286e+00
R32513 n0_4741_5385 n0_4929_5385 1.074286e+00
R32514 n0_4929_5385 n0_5866_5385 5.354286e+00
R32515 n0_5866_5385 n0_5958_5385 5.257143e-01
R32516 n0_5958_5385 n0_6054_5385 5.485714e-01
R32517 n0_6054_5385 n0_6146_5385 5.257143e-01
R32518 n0_6146_5385 n0_8116_5385 1.125714e+01
R32519 n0_8116_5385 n0_8208_5385 5.257143e-01
R32520 n0_8208_5385 n0_8304_5385 5.485714e-01
R32521 n0_8304_5385 n0_8396_5385 5.257143e-01
R32522 n0_8396_5385 n0_10366_5385 1.125714e+01
R32523 n0_10366_5385 n0_10458_5385 5.257143e-01
R32524 n0_10458_5385 n0_10554_5385 5.485714e-01
R32525 n0_10554_5385 n0_10646_5385 5.257143e-01
R32526 n0_10646_5385 n0_12616_5385 1.125714e+01
R32527 n0_12616_5385 n0_12708_5385 5.257143e-01
R32528 n0_12708_5385 n0_12804_5385 5.485714e-01
R32529 n0_12804_5385 n0_12896_5385 5.257143e-01
R32530 n0_12896_5385 n0_14866_5385 1.125714e+01
R32531 n0_14866_5385 n0_14958_5385 5.257143e-01
R32532 n0_14958_5385 n0_15054_5385 5.485714e-01
R32533 n0_15054_5385 n0_15146_5385 5.257143e-01
R32534 n0_15146_5385 n0_15991_5385 4.828571e+00
R32535 n0_15991_5385 n0_16179_5385 1.074286e+00
R32536 n0_16179_5385 n0_17116_5385 5.354286e+00
R32537 n0_17116_5385 n0_17304_5385 1.074286e+00
R32538 n0_17304_5385 n0_18241_5385 5.354286e+00
R32539 n0_18241_5385 n0_18429_5385 1.074286e+00
R32540 n0_18429_5385 n0_19366_5385 5.354286e+00
R32541 n0_19366_5385 n0_19554_5385 1.074286e+00
R32542 n0_19554_5385 n0_20491_5385 5.354286e+00
R32543 n0_20491_5385 n0_20679_5385 1.074286e+00
R32544 n0_241_5418 n0_429_5418 1.074286e+00
R32545 n0_429_5418 n0_1366_5418 5.354286e+00
R32546 n0_1366_5418 n0_1554_5418 1.074286e+00
R32547 n0_1554_5418 n0_2491_5418 5.354286e+00
R32548 n0_2491_5418 n0_2679_5418 1.074286e+00
R32549 n0_2679_5418 n0_3616_5418 5.354286e+00
R32550 n0_3616_5418 n0_3804_5418 1.074286e+00
R32551 n0_3804_5418 n0_4741_5418 5.354286e+00
R32552 n0_4741_5418 n0_4929_5418 1.074286e+00
R32553 n0_4929_5418 n0_5866_5418 5.354286e+00
R32554 n0_5866_5418 n0_5958_5418 5.257143e-01
R32555 n0_5958_5418 n0_6054_5418 5.485714e-01
R32556 n0_6054_5418 n0_6146_5418 5.257143e-01
R32557 n0_6146_5418 n0_8116_5418 1.125714e+01
R32558 n0_8116_5418 n0_8208_5418 5.257143e-01
R32559 n0_8208_5418 n0_8304_5418 5.485714e-01
R32560 n0_8304_5418 n0_8396_5418 5.257143e-01
R32561 n0_8396_5418 n0_10366_5418 1.125714e+01
R32562 n0_10366_5418 n0_10458_5418 5.257143e-01
R32563 n0_10458_5418 n0_10554_5418 5.485714e-01
R32564 n0_10554_5418 n0_10646_5418 5.257143e-01
R32565 n0_10646_5418 n0_12616_5418 1.125714e+01
R32566 n0_12616_5418 n0_12708_5418 5.257143e-01
R32567 n0_12708_5418 n0_12804_5418 5.485714e-01
R32568 n0_12804_5418 n0_12896_5418 5.257143e-01
R32569 n0_12896_5418 n0_14866_5418 1.125714e+01
R32570 n0_14866_5418 n0_14958_5418 5.257143e-01
R32571 n0_14958_5418 n0_15054_5418 5.485714e-01
R32572 n0_15054_5418 n0_15146_5418 5.257143e-01
R32573 n0_15146_5418 n0_15991_5418 4.828571e+00
R32574 n0_15991_5418 n0_16179_5418 1.074286e+00
R32575 n0_16179_5418 n0_17116_5418 5.354286e+00
R32576 n0_17116_5418 n0_17304_5418 1.074286e+00
R32577 n0_17304_5418 n0_18241_5418 5.354286e+00
R32578 n0_18241_5418 n0_18429_5418 1.074286e+00
R32579 n0_18429_5418 n0_19366_5418 5.354286e+00
R32580 n0_19366_5418 n0_19554_5418 1.074286e+00
R32581 n0_19554_5418 n0_20491_5418 5.354286e+00
R32582 n0_20491_5418 n0_20679_5418 1.074286e+00
R32583 n0_241_5601 n0_429_5601 1.074286e+00
R32584 n0_429_5601 n0_1366_5601 5.354286e+00
R32585 n0_1366_5601 n0_1554_5601 1.074286e+00
R32586 n0_1554_5601 n0_2491_5601 5.354286e+00
R32587 n0_2491_5601 n0_2679_5601 1.074286e+00
R32588 n0_2679_5601 n0_3616_5601 5.354286e+00
R32589 n0_3616_5601 n0_3804_5601 1.074286e+00
R32590 n0_3804_5601 n0_4741_5601 5.354286e+00
R32591 n0_4741_5601 n0_4929_5601 1.074286e+00
R32592 n0_4929_5601 n0_5866_5601 5.354286e+00
R32593 n0_5866_5601 n0_5958_5601 5.257143e-01
R32594 n0_5958_5601 n0_6054_5601 5.485714e-01
R32595 n0_6054_5601 n0_6146_5601 5.257143e-01
R32596 n0_6146_5601 n0_8116_5601 1.125714e+01
R32597 n0_8116_5601 n0_8208_5601 5.257143e-01
R32598 n0_8208_5601 n0_8304_5601 5.485714e-01
R32599 n0_8304_5601 n0_8396_5601 5.257143e-01
R32600 n0_8396_5601 n0_10366_5601 1.125714e+01
R32601 n0_10366_5601 n0_10458_5601 5.257143e-01
R32602 n0_10458_5601 n0_10554_5601 5.485714e-01
R32603 n0_10554_5601 n0_10646_5601 5.257143e-01
R32604 n0_10646_5601 n0_12616_5601 1.125714e+01
R32605 n0_12616_5601 n0_12708_5601 5.257143e-01
R32606 n0_12708_5601 n0_12804_5601 5.485714e-01
R32607 n0_12804_5601 n0_12896_5601 5.257143e-01
R32608 n0_12896_5601 n0_14866_5601 1.125714e+01
R32609 n0_14866_5601 n0_14958_5601 5.257143e-01
R32610 n0_14958_5601 n0_15054_5601 5.485714e-01
R32611 n0_15054_5601 n0_15146_5601 5.257143e-01
R32612 n0_15146_5601 n0_15991_5601 4.828571e+00
R32613 n0_15991_5601 n0_16179_5601 1.074286e+00
R32614 n0_16179_5601 n0_17116_5601 5.354286e+00
R32615 n0_17116_5601 n0_17304_5601 1.074286e+00
R32616 n0_17304_5601 n0_18241_5601 5.354286e+00
R32617 n0_18241_5601 n0_18429_5601 1.074286e+00
R32618 n0_18429_5601 n0_19366_5601 5.354286e+00
R32619 n0_19366_5601 n0_19554_5601 1.074286e+00
R32620 n0_19554_5601 n0_20491_5601 5.354286e+00
R32621 n0_20491_5601 n0_20679_5601 1.074286e+00
R32622 n0_241_5634 n0_429_5634 1.074286e+00
R32623 n0_429_5634 n0_1366_5634 5.354286e+00
R32624 n0_1366_5634 n0_1554_5634 1.074286e+00
R32625 n0_1554_5634 n0_2491_5634 5.354286e+00
R32626 n0_2491_5634 n0_2679_5634 1.074286e+00
R32627 n0_2679_5634 n0_3616_5634 5.354286e+00
R32628 n0_3616_5634 n0_3804_5634 1.074286e+00
R32629 n0_3804_5634 n0_4741_5634 5.354286e+00
R32630 n0_4741_5634 n0_4929_5634 1.074286e+00
R32631 n0_4929_5634 n0_5866_5634 5.354286e+00
R32632 n0_5866_5634 n0_5958_5634 5.257143e-01
R32633 n0_5958_5634 n0_6054_5634 5.485714e-01
R32634 n0_6054_5634 n0_6146_5634 5.257143e-01
R32635 n0_6146_5634 n0_8116_5634 1.125714e+01
R32636 n0_8116_5634 n0_8208_5634 5.257143e-01
R32637 n0_8208_5634 n0_8304_5634 5.485714e-01
R32638 n0_8304_5634 n0_8396_5634 5.257143e-01
R32639 n0_8396_5634 n0_10366_5634 1.125714e+01
R32640 n0_10366_5634 n0_10458_5634 5.257143e-01
R32641 n0_10458_5634 n0_10554_5634 5.485714e-01
R32642 n0_10554_5634 n0_10646_5634 5.257143e-01
R32643 n0_10646_5634 n0_12616_5634 1.125714e+01
R32644 n0_12616_5634 n0_12708_5634 5.257143e-01
R32645 n0_12708_5634 n0_12804_5634 5.485714e-01
R32646 n0_12804_5634 n0_12896_5634 5.257143e-01
R32647 n0_12896_5634 n0_14866_5634 1.125714e+01
R32648 n0_14866_5634 n0_14958_5634 5.257143e-01
R32649 n0_14958_5634 n0_15054_5634 5.485714e-01
R32650 n0_15054_5634 n0_15146_5634 5.257143e-01
R32651 n0_15146_5634 n0_15991_5634 4.828571e+00
R32652 n0_15991_5634 n0_16179_5634 1.074286e+00
R32653 n0_16179_5634 n0_17116_5634 5.354286e+00
R32654 n0_17116_5634 n0_17304_5634 1.074286e+00
R32655 n0_17304_5634 n0_18241_5634 5.354286e+00
R32656 n0_18241_5634 n0_18429_5634 1.074286e+00
R32657 n0_18429_5634 n0_19366_5634 5.354286e+00
R32658 n0_19366_5634 n0_19554_5634 1.074286e+00
R32659 n0_19554_5634 n0_20491_5634 5.354286e+00
R32660 n0_20491_5634 n0_20679_5634 1.074286e+00
R32661 n0_241_5817 n0_429_5817 1.074286e+00
R32662 n0_429_5817 n0_1366_5817 5.354286e+00
R32663 n0_1366_5817 n0_1554_5817 1.074286e+00
R32664 n0_1554_5817 n0_2491_5817 5.354286e+00
R32665 n0_2491_5817 n0_2679_5817 1.074286e+00
R32666 n0_2679_5817 n0_3616_5817 5.354286e+00
R32667 n0_3616_5817 n0_3804_5817 1.074286e+00
R32668 n0_3804_5817 n0_4741_5817 5.354286e+00
R32669 n0_4741_5817 n0_4929_5817 1.074286e+00
R32670 n0_4929_5817 n0_5866_5817 5.354286e+00
R32671 n0_5866_5817 n0_5958_5817 5.257143e-01
R32672 n0_5958_5817 n0_6054_5817 5.485714e-01
R32673 n0_6054_5817 n0_6146_5817 5.257143e-01
R32674 n0_6146_5817 n0_8116_5817 1.125714e+01
R32675 n0_8116_5817 n0_8208_5817 5.257143e-01
R32676 n0_8208_5817 n0_8304_5817 5.485714e-01
R32677 n0_8304_5817 n0_8396_5817 5.257143e-01
R32678 n0_8396_5817 n0_10366_5817 1.125714e+01
R32679 n0_10366_5817 n0_10458_5817 5.257143e-01
R32680 n0_10458_5817 n0_10554_5817 5.485714e-01
R32681 n0_10554_5817 n0_10646_5817 5.257143e-01
R32682 n0_10646_5817 n0_12616_5817 1.125714e+01
R32683 n0_12616_5817 n0_12708_5817 5.257143e-01
R32684 n0_12708_5817 n0_12804_5817 5.485714e-01
R32685 n0_12804_5817 n0_12896_5817 5.257143e-01
R32686 n0_12896_5817 n0_14866_5817 1.125714e+01
R32687 n0_14866_5817 n0_14958_5817 5.257143e-01
R32688 n0_14958_5817 n0_15054_5817 5.485714e-01
R32689 n0_15054_5817 n0_15146_5817 5.257143e-01
R32690 n0_15146_5817 n0_15991_5817 4.828571e+00
R32691 n0_15991_5817 n0_16179_5817 1.074286e+00
R32692 n0_16179_5817 n0_17116_5817 5.354286e+00
R32693 n0_17116_5817 n0_17304_5817 1.074286e+00
R32694 n0_17304_5817 n0_18241_5817 5.354286e+00
R32695 n0_18241_5817 n0_18429_5817 1.074286e+00
R32696 n0_18429_5817 n0_19366_5817 5.354286e+00
R32697 n0_19366_5817 n0_19554_5817 1.074286e+00
R32698 n0_19554_5817 n0_20491_5817 5.354286e+00
R32699 n0_20491_5817 n0_20679_5817 1.074286e+00
R32700 n0_241_5850 n0_429_5850 1.074286e+00
R32701 n0_429_5850 n0_1366_5850 5.354286e+00
R32702 n0_1366_5850 n0_1554_5850 1.074286e+00
R32703 n0_1554_5850 n0_2491_5850 5.354286e+00
R32704 n0_2491_5850 n0_2679_5850 1.074286e+00
R32705 n0_2679_5850 n0_3616_5850 5.354286e+00
R32706 n0_3616_5850 n0_3804_5850 1.074286e+00
R32707 n0_3804_5850 n0_4741_5850 5.354286e+00
R32708 n0_4741_5850 n0_4929_5850 1.074286e+00
R32709 n0_4929_5850 n0_5866_5850 5.354286e+00
R32710 n0_5866_5850 n0_5958_5850 5.257143e-01
R32711 n0_5958_5850 n0_6054_5850 5.485714e-01
R32712 n0_6054_5850 n0_6146_5850 5.257143e-01
R32713 n0_6146_5850 n0_8116_5850 1.125714e+01
R32714 n0_8116_5850 n0_8208_5850 5.257143e-01
R32715 n0_8208_5850 n0_8304_5850 5.485714e-01
R32716 n0_8304_5850 n0_8396_5850 5.257143e-01
R32717 n0_8396_5850 n0_10366_5850 1.125714e+01
R32718 n0_10366_5850 n0_10458_5850 5.257143e-01
R32719 n0_10458_5850 n0_10554_5850 5.485714e-01
R32720 n0_10554_5850 n0_10646_5850 5.257143e-01
R32721 n0_10646_5850 n0_12616_5850 1.125714e+01
R32722 n0_12616_5850 n0_12708_5850 5.257143e-01
R32723 n0_12708_5850 n0_12804_5850 5.485714e-01
R32724 n0_12804_5850 n0_12896_5850 5.257143e-01
R32725 n0_12896_5850 n0_14866_5850 1.125714e+01
R32726 n0_14866_5850 n0_14958_5850 5.257143e-01
R32727 n0_14958_5850 n0_15054_5850 5.485714e-01
R32728 n0_15054_5850 n0_15146_5850 5.257143e-01
R32729 n0_15146_5850 n0_15991_5850 4.828571e+00
R32730 n0_15991_5850 n0_16179_5850 1.074286e+00
R32731 n0_16179_5850 n0_17116_5850 5.354286e+00
R32732 n0_17116_5850 n0_17304_5850 1.074286e+00
R32733 n0_17304_5850 n0_18241_5850 5.354286e+00
R32734 n0_18241_5850 n0_18429_5850 1.074286e+00
R32735 n0_18429_5850 n0_19366_5850 5.354286e+00
R32736 n0_19366_5850 n0_19554_5850 1.074286e+00
R32737 n0_19554_5850 n0_20491_5850 5.354286e+00
R32738 n0_20491_5850 n0_20679_5850 1.074286e+00
R32739 n0_241_6033 n0_380_6033 7.942857e-01
R32740 n0_380_6033 n0_429_6033 2.800000e-01
R32741 n0_429_6033 n0_1366_6033 5.354286e+00
R32742 n0_1366_6033 n0_1505_6033 7.942857e-01
R32743 n0_1505_6033 n0_1554_6033 2.800000e-01
R32744 n0_1554_6033 n0_2491_6033 5.354286e+00
R32745 n0_2491_6033 n0_2630_6033 7.942857e-01
R32746 n0_2630_6033 n0_2679_6033 2.800000e-01
R32747 n0_2679_6033 n0_3616_6033 5.354286e+00
R32748 n0_3616_6033 n0_3755_6033 7.942857e-01
R32749 n0_3755_6033 n0_3804_6033 2.800000e-01
R32750 n0_3804_6033 n0_4741_6033 5.354286e+00
R32751 n0_4741_6033 n0_4880_6033 7.942857e-01
R32752 n0_4880_6033 n0_4929_6033 2.800000e-01
R32753 n0_4929_6033 n0_5866_6033 5.354286e+00
R32754 n0_5866_6033 n0_5958_6033 5.257143e-01
R32755 n0_5958_6033 n0_6005_6033 2.685714e-01
R32756 n0_6005_6033 n0_6054_6033 2.800000e-01
R32757 n0_6054_6033 n0_6146_6033 5.257143e-01
R32758 n0_6146_6033 n0_8116_6033 1.125714e+01
R32759 n0_8116_6033 n0_8208_6033 5.257143e-01
R32760 n0_8208_6033 n0_8255_6033 2.685714e-01
R32761 n0_8255_6033 n0_8304_6033 2.800000e-01
R32762 n0_8304_6033 n0_8396_6033 5.257143e-01
R32763 n0_8396_6033 n0_10366_6033 1.125714e+01
R32764 n0_10366_6033 n0_10458_6033 5.257143e-01
R32765 n0_10458_6033 n0_10505_6033 2.685714e-01
R32766 n0_10505_6033 n0_10554_6033 2.800000e-01
R32767 n0_10554_6033 n0_10646_6033 5.257143e-01
R32768 n0_10646_6033 n0_12616_6033 1.125714e+01
R32769 n0_12616_6033 n0_12708_6033 5.257143e-01
R32770 n0_12708_6033 n0_12755_6033 2.685714e-01
R32771 n0_12755_6033 n0_12804_6033 2.800000e-01
R32772 n0_12804_6033 n0_12896_6033 5.257143e-01
R32773 n0_12896_6033 n0_14866_6033 1.125714e+01
R32774 n0_14866_6033 n0_14958_6033 5.257143e-01
R32775 n0_14958_6033 n0_15005_6033 2.685714e-01
R32776 n0_15005_6033 n0_15054_6033 2.800000e-01
R32777 n0_15054_6033 n0_15146_6033 5.257143e-01
R32778 n0_15146_6033 n0_15991_6033 4.828571e+00
R32779 n0_15991_6033 n0_16130_6033 7.942857e-01
R32780 n0_16130_6033 n0_16179_6033 2.800000e-01
R32781 n0_16179_6033 n0_17116_6033 5.354286e+00
R32782 n0_17116_6033 n0_17255_6033 7.942857e-01
R32783 n0_17255_6033 n0_17304_6033 2.800000e-01
R32784 n0_17304_6033 n0_18241_6033 5.354286e+00
R32785 n0_18241_6033 n0_18380_6033 7.942857e-01
R32786 n0_18380_6033 n0_18429_6033 2.800000e-01
R32787 n0_18429_6033 n0_19366_6033 5.354286e+00
R32788 n0_19366_6033 n0_19505_6033 7.942857e-01
R32789 n0_19505_6033 n0_19554_6033 2.800000e-01
R32790 n0_19554_6033 n0_20491_6033 5.354286e+00
R32791 n0_20491_6033 n0_20630_6033 7.942857e-01
R32792 n0_20630_6033 n0_20679_6033 2.800000e-01
R32793 n0_241_6066 n0_380_6066 7.942857e-01
R32794 n0_380_6066 n0_429_6066 2.800000e-01
R32795 n0_429_6066 n0_1366_6066 5.354286e+00
R32796 n0_1366_6066 n0_1505_6066 7.942857e-01
R32797 n0_1505_6066 n0_1554_6066 2.800000e-01
R32798 n0_1554_6066 n0_2491_6066 5.354286e+00
R32799 n0_2491_6066 n0_2630_6066 7.942857e-01
R32800 n0_2630_6066 n0_2679_6066 2.800000e-01
R32801 n0_2679_6066 n0_3616_6066 5.354286e+00
R32802 n0_3616_6066 n0_3755_6066 7.942857e-01
R32803 n0_3755_6066 n0_3804_6066 2.800000e-01
R32804 n0_3804_6066 n0_4741_6066 5.354286e+00
R32805 n0_4741_6066 n0_4880_6066 7.942857e-01
R32806 n0_4880_6066 n0_4929_6066 2.800000e-01
R32807 n0_4929_6066 n0_5866_6066 5.354286e+00
R32808 n0_5866_6066 n0_5958_6066 5.257143e-01
R32809 n0_5958_6066 n0_6005_6066 2.685714e-01
R32810 n0_6005_6066 n0_6054_6066 2.800000e-01
R32811 n0_6054_6066 n0_6146_6066 5.257143e-01
R32812 n0_6146_6066 n0_8116_6066 1.125714e+01
R32813 n0_8116_6066 n0_8208_6066 5.257143e-01
R32814 n0_8208_6066 n0_8255_6066 2.685714e-01
R32815 n0_8255_6066 n0_8304_6066 2.800000e-01
R32816 n0_8304_6066 n0_8396_6066 5.257143e-01
R32817 n0_8396_6066 n0_10366_6066 1.125714e+01
R32818 n0_10366_6066 n0_10458_6066 5.257143e-01
R32819 n0_10458_6066 n0_10505_6066 2.685714e-01
R32820 n0_10505_6066 n0_10554_6066 2.800000e-01
R32821 n0_10554_6066 n0_10646_6066 5.257143e-01
R32822 n0_10646_6066 n0_12616_6066 1.125714e+01
R32823 n0_12616_6066 n0_12708_6066 5.257143e-01
R32824 n0_12708_6066 n0_12755_6066 2.685714e-01
R32825 n0_12755_6066 n0_12804_6066 2.800000e-01
R32826 n0_12804_6066 n0_12896_6066 5.257143e-01
R32827 n0_12896_6066 n0_14866_6066 1.125714e+01
R32828 n0_14866_6066 n0_14958_6066 5.257143e-01
R32829 n0_14958_6066 n0_15005_6066 2.685714e-01
R32830 n0_15005_6066 n0_15054_6066 2.800000e-01
R32831 n0_15054_6066 n0_15146_6066 5.257143e-01
R32832 n0_15146_6066 n0_15991_6066 4.828571e+00
R32833 n0_15991_6066 n0_16130_6066 7.942857e-01
R32834 n0_16130_6066 n0_16179_6066 2.800000e-01
R32835 n0_16179_6066 n0_17116_6066 5.354286e+00
R32836 n0_17116_6066 n0_17255_6066 7.942857e-01
R32837 n0_17255_6066 n0_17304_6066 2.800000e-01
R32838 n0_17304_6066 n0_18241_6066 5.354286e+00
R32839 n0_18241_6066 n0_18380_6066 7.942857e-01
R32840 n0_18380_6066 n0_18429_6066 2.800000e-01
R32841 n0_18429_6066 n0_19366_6066 5.354286e+00
R32842 n0_19366_6066 n0_19505_6066 7.942857e-01
R32843 n0_19505_6066 n0_19554_6066 2.800000e-01
R32844 n0_19554_6066 n0_20491_6066 5.354286e+00
R32845 n0_20491_6066 n0_20630_6066 7.942857e-01
R32846 n0_20630_6066 n0_20679_6066 2.800000e-01
R32847 n0_241_6249 n0_429_6249 1.074286e+00
R32848 n0_429_6249 n0_1366_6249 5.354286e+00
R32849 n0_1366_6249 n0_1554_6249 1.074286e+00
R32850 n0_1554_6249 n0_2491_6249 5.354286e+00
R32851 n0_2491_6249 n0_2679_6249 1.074286e+00
R32852 n0_2679_6249 n0_3616_6249 5.354286e+00
R32853 n0_3616_6249 n0_3804_6249 1.074286e+00
R32854 n0_3804_6249 n0_4741_6249 5.354286e+00
R32855 n0_4741_6249 n0_4929_6249 1.074286e+00
R32856 n0_4929_6249 n0_5866_6249 5.354286e+00
R32857 n0_5866_6249 n0_6054_6249 1.074286e+00
R32858 n0_6054_6249 n0_8116_6249 1.178286e+01
R32859 n0_8116_6249 n0_8208_6249 5.257143e-01
R32860 n0_8208_6249 n0_8304_6249 5.485714e-01
R32861 n0_8304_6249 n0_8396_6249 5.257143e-01
R32862 n0_8396_6249 n0_10366_6249 1.125714e+01
R32863 n0_10366_6249 n0_10458_6249 5.257143e-01
R32864 n0_10458_6249 n0_10554_6249 5.485714e-01
R32865 n0_10554_6249 n0_10646_6249 5.257143e-01
R32866 n0_10646_6249 n0_12616_6249 1.125714e+01
R32867 n0_12616_6249 n0_12708_6249 5.257143e-01
R32868 n0_12708_6249 n0_12804_6249 5.485714e-01
R32869 n0_12804_6249 n0_12896_6249 5.257143e-01
R32870 n0_12896_6249 n0_14866_6249 1.125714e+01
R32871 n0_14866_6249 n0_15054_6249 1.074286e+00
R32872 n0_15054_6249 n0_15991_6249 5.354286e+00
R32873 n0_15991_6249 n0_16179_6249 1.074286e+00
R32874 n0_16179_6249 n0_17116_6249 5.354286e+00
R32875 n0_17116_6249 n0_17304_6249 1.074286e+00
R32876 n0_17304_6249 n0_18241_6249 5.354286e+00
R32877 n0_18241_6249 n0_18429_6249 1.074286e+00
R32878 n0_18429_6249 n0_19366_6249 5.354286e+00
R32879 n0_19366_6249 n0_19554_6249 1.074286e+00
R32880 n0_19554_6249 n0_20491_6249 5.354286e+00
R32881 n0_20491_6249 n0_20679_6249 1.074286e+00
R32882 n0_241_6282 n0_429_6282 1.074286e+00
R32883 n0_429_6282 n0_1366_6282 5.354286e+00
R32884 n0_1366_6282 n0_1554_6282 1.074286e+00
R32885 n0_1554_6282 n0_2491_6282 5.354286e+00
R32886 n0_2491_6282 n0_2679_6282 1.074286e+00
R32887 n0_2679_6282 n0_3616_6282 5.354286e+00
R32888 n0_3616_6282 n0_3804_6282 1.074286e+00
R32889 n0_3804_6282 n0_4741_6282 5.354286e+00
R32890 n0_4741_6282 n0_4929_6282 1.074286e+00
R32891 n0_4929_6282 n0_5866_6282 5.354286e+00
R32892 n0_5866_6282 n0_6054_6282 1.074286e+00
R32893 n0_6054_6282 n0_8116_6282 1.178286e+01
R32894 n0_8116_6282 n0_8208_6282 5.257143e-01
R32895 n0_8208_6282 n0_8304_6282 5.485714e-01
R32896 n0_8304_6282 n0_8396_6282 5.257143e-01
R32897 n0_8396_6282 n0_10366_6282 1.125714e+01
R32898 n0_10366_6282 n0_10458_6282 5.257143e-01
R32899 n0_10458_6282 n0_10554_6282 5.485714e-01
R32900 n0_10554_6282 n0_10646_6282 5.257143e-01
R32901 n0_10646_6282 n0_12616_6282 1.125714e+01
R32902 n0_12616_6282 n0_12708_6282 5.257143e-01
R32903 n0_12708_6282 n0_12804_6282 5.485714e-01
R32904 n0_12804_6282 n0_12896_6282 5.257143e-01
R32905 n0_12896_6282 n0_14866_6282 1.125714e+01
R32906 n0_14866_6282 n0_15054_6282 1.074286e+00
R32907 n0_15054_6282 n0_15991_6282 5.354286e+00
R32908 n0_15991_6282 n0_16179_6282 1.074286e+00
R32909 n0_16179_6282 n0_17116_6282 5.354286e+00
R32910 n0_17116_6282 n0_17304_6282 1.074286e+00
R32911 n0_17304_6282 n0_18241_6282 5.354286e+00
R32912 n0_18241_6282 n0_18429_6282 1.074286e+00
R32913 n0_18429_6282 n0_19366_6282 5.354286e+00
R32914 n0_19366_6282 n0_19554_6282 1.074286e+00
R32915 n0_19554_6282 n0_20491_6282 5.354286e+00
R32916 n0_20491_6282 n0_20679_6282 1.074286e+00
R32917 n0_241_6465 n0_429_6465 1.074286e+00
R32918 n0_429_6465 n0_1366_6465 5.354286e+00
R32919 n0_1366_6465 n0_1554_6465 1.074286e+00
R32920 n0_1554_6465 n0_2491_6465 5.354286e+00
R32921 n0_2491_6465 n0_2679_6465 1.074286e+00
R32922 n0_2679_6465 n0_3616_6465 5.354286e+00
R32923 n0_3616_6465 n0_3804_6465 1.074286e+00
R32924 n0_3804_6465 n0_4741_6465 5.354286e+00
R32925 n0_4741_6465 n0_4929_6465 1.074286e+00
R32926 n0_4929_6465 n0_5866_6465 5.354286e+00
R32927 n0_5866_6465 n0_6054_6465 1.074286e+00
R32928 n0_6054_6465 n0_8116_6465 1.178286e+01
R32929 n0_8116_6465 n0_8208_6465 5.257143e-01
R32930 n0_8208_6465 n0_8304_6465 5.485714e-01
R32931 n0_8304_6465 n0_8396_6465 5.257143e-01
R32932 n0_8396_6465 n0_10366_6465 1.125714e+01
R32933 n0_10366_6465 n0_10458_6465 5.257143e-01
R32934 n0_10458_6465 n0_10554_6465 5.485714e-01
R32935 n0_10554_6465 n0_10646_6465 5.257143e-01
R32936 n0_10646_6465 n0_12616_6465 1.125714e+01
R32937 n0_12616_6465 n0_12708_6465 5.257143e-01
R32938 n0_12708_6465 n0_12804_6465 5.485714e-01
R32939 n0_12804_6465 n0_12896_6465 5.257143e-01
R32940 n0_12896_6465 n0_14866_6465 1.125714e+01
R32941 n0_14866_6465 n0_15054_6465 1.074286e+00
R32942 n0_15054_6465 n0_15991_6465 5.354286e+00
R32943 n0_15991_6465 n0_16179_6465 1.074286e+00
R32944 n0_16179_6465 n0_17116_6465 5.354286e+00
R32945 n0_17116_6465 n0_17304_6465 1.074286e+00
R32946 n0_17304_6465 n0_18241_6465 5.354286e+00
R32947 n0_18241_6465 n0_18429_6465 1.074286e+00
R32948 n0_18429_6465 n0_19366_6465 5.354286e+00
R32949 n0_19366_6465 n0_19554_6465 1.074286e+00
R32950 n0_19554_6465 n0_20491_6465 5.354286e+00
R32951 n0_20491_6465 n0_20679_6465 1.074286e+00
R32952 n0_241_6498 n0_429_6498 1.074286e+00
R32953 n0_429_6498 n0_1366_6498 5.354286e+00
R32954 n0_1366_6498 n0_1554_6498 1.074286e+00
R32955 n0_1554_6498 n0_2491_6498 5.354286e+00
R32956 n0_2491_6498 n0_2679_6498 1.074286e+00
R32957 n0_2679_6498 n0_3616_6498 5.354286e+00
R32958 n0_3616_6498 n0_3804_6498 1.074286e+00
R32959 n0_3804_6498 n0_4741_6498 5.354286e+00
R32960 n0_4741_6498 n0_4929_6498 1.074286e+00
R32961 n0_4929_6498 n0_5866_6498 5.354286e+00
R32962 n0_5866_6498 n0_6054_6498 1.074286e+00
R32963 n0_6054_6498 n0_8116_6498 1.178286e+01
R32964 n0_8116_6498 n0_8208_6498 5.257143e-01
R32965 n0_8208_6498 n0_8304_6498 5.485714e-01
R32966 n0_8304_6498 n0_8396_6498 5.257143e-01
R32967 n0_8396_6498 n0_10366_6498 1.125714e+01
R32968 n0_10366_6498 n0_10458_6498 5.257143e-01
R32969 n0_10458_6498 n0_10554_6498 5.485714e-01
R32970 n0_10554_6498 n0_10646_6498 5.257143e-01
R32971 n0_10646_6498 n0_12616_6498 1.125714e+01
R32972 n0_12616_6498 n0_12708_6498 5.257143e-01
R32973 n0_12708_6498 n0_12804_6498 5.485714e-01
R32974 n0_12804_6498 n0_12896_6498 5.257143e-01
R32975 n0_12896_6498 n0_14866_6498 1.125714e+01
R32976 n0_14866_6498 n0_15054_6498 1.074286e+00
R32977 n0_15054_6498 n0_15991_6498 5.354286e+00
R32978 n0_15991_6498 n0_16179_6498 1.074286e+00
R32979 n0_16179_6498 n0_17116_6498 5.354286e+00
R32980 n0_17116_6498 n0_17304_6498 1.074286e+00
R32981 n0_17304_6498 n0_18241_6498 5.354286e+00
R32982 n0_18241_6498 n0_18429_6498 1.074286e+00
R32983 n0_18429_6498 n0_19366_6498 5.354286e+00
R32984 n0_19366_6498 n0_19554_6498 1.074286e+00
R32985 n0_19554_6498 n0_20491_6498 5.354286e+00
R32986 n0_20491_6498 n0_20679_6498 1.074286e+00
R32987 n0_241_6681 n0_429_6681 1.074286e+00
R32988 n0_429_6681 n0_1366_6681 5.354286e+00
R32989 n0_1366_6681 n0_1554_6681 1.074286e+00
R32990 n0_1554_6681 n0_2491_6681 5.354286e+00
R32991 n0_2491_6681 n0_2679_6681 1.074286e+00
R32992 n0_2679_6681 n0_3616_6681 5.354286e+00
R32993 n0_3616_6681 n0_3804_6681 1.074286e+00
R32994 n0_3804_6681 n0_4741_6681 5.354286e+00
R32995 n0_4741_6681 n0_4929_6681 1.074286e+00
R32996 n0_4929_6681 n0_5866_6681 5.354286e+00
R32997 n0_5866_6681 n0_6054_6681 1.074286e+00
R32998 n0_6054_6681 n0_8116_6681 1.178286e+01
R32999 n0_8116_6681 n0_8208_6681 5.257143e-01
R33000 n0_8208_6681 n0_8304_6681 5.485714e-01
R33001 n0_8304_6681 n0_8396_6681 5.257143e-01
R33002 n0_8396_6681 n0_10366_6681 1.125714e+01
R33003 n0_10366_6681 n0_10458_6681 5.257143e-01
R33004 n0_10458_6681 n0_10554_6681 5.485714e-01
R33005 n0_10554_6681 n0_10646_6681 5.257143e-01
R33006 n0_10646_6681 n0_12616_6681 1.125714e+01
R33007 n0_12616_6681 n0_12708_6681 5.257143e-01
R33008 n0_12708_6681 n0_12804_6681 5.485714e-01
R33009 n0_12804_6681 n0_12896_6681 5.257143e-01
R33010 n0_12896_6681 n0_14866_6681 1.125714e+01
R33011 n0_14866_6681 n0_15054_6681 1.074286e+00
R33012 n0_15054_6681 n0_15991_6681 5.354286e+00
R33013 n0_15991_6681 n0_16179_6681 1.074286e+00
R33014 n0_16179_6681 n0_17116_6681 5.354286e+00
R33015 n0_17116_6681 n0_17304_6681 1.074286e+00
R33016 n0_17304_6681 n0_18241_6681 5.354286e+00
R33017 n0_18241_6681 n0_18429_6681 1.074286e+00
R33018 n0_18429_6681 n0_19366_6681 5.354286e+00
R33019 n0_19366_6681 n0_19554_6681 1.074286e+00
R33020 n0_19554_6681 n0_20491_6681 5.354286e+00
R33021 n0_20491_6681 n0_20679_6681 1.074286e+00
R33022 n0_241_6714 n0_429_6714 1.074286e+00
R33023 n0_429_6714 n0_1366_6714 5.354286e+00
R33024 n0_1366_6714 n0_1554_6714 1.074286e+00
R33025 n0_1554_6714 n0_2491_6714 5.354286e+00
R33026 n0_2491_6714 n0_2679_6714 1.074286e+00
R33027 n0_2679_6714 n0_3616_6714 5.354286e+00
R33028 n0_3616_6714 n0_3804_6714 1.074286e+00
R33029 n0_3804_6714 n0_4741_6714 5.354286e+00
R33030 n0_4741_6714 n0_4929_6714 1.074286e+00
R33031 n0_4929_6714 n0_5866_6714 5.354286e+00
R33032 n0_5866_6714 n0_6054_6714 1.074286e+00
R33033 n0_6054_6714 n0_8116_6714 1.178286e+01
R33034 n0_8116_6714 n0_8208_6714 5.257143e-01
R33035 n0_8208_6714 n0_8304_6714 5.485714e-01
R33036 n0_8304_6714 n0_8396_6714 5.257143e-01
R33037 n0_8396_6714 n0_10366_6714 1.125714e+01
R33038 n0_10366_6714 n0_10458_6714 5.257143e-01
R33039 n0_10458_6714 n0_10554_6714 5.485714e-01
R33040 n0_10554_6714 n0_10646_6714 5.257143e-01
R33041 n0_10646_6714 n0_12616_6714 1.125714e+01
R33042 n0_12616_6714 n0_12708_6714 5.257143e-01
R33043 n0_12708_6714 n0_12804_6714 5.485714e-01
R33044 n0_12804_6714 n0_12896_6714 5.257143e-01
R33045 n0_12896_6714 n0_14866_6714 1.125714e+01
R33046 n0_14866_6714 n0_15054_6714 1.074286e+00
R33047 n0_15054_6714 n0_15991_6714 5.354286e+00
R33048 n0_15991_6714 n0_16179_6714 1.074286e+00
R33049 n0_16179_6714 n0_17116_6714 5.354286e+00
R33050 n0_17116_6714 n0_17304_6714 1.074286e+00
R33051 n0_17304_6714 n0_18241_6714 5.354286e+00
R33052 n0_18241_6714 n0_18429_6714 1.074286e+00
R33053 n0_18429_6714 n0_19366_6714 5.354286e+00
R33054 n0_19366_6714 n0_19554_6714 1.074286e+00
R33055 n0_19554_6714 n0_20491_6714 5.354286e+00
R33056 n0_20491_6714 n0_20679_6714 1.074286e+00
R33057 n0_241_6897 n0_429_6897 1.074286e+00
R33058 n0_429_6897 n0_1366_6897 5.354286e+00
R33059 n0_1366_6897 n0_1554_6897 1.074286e+00
R33060 n0_1554_6897 n0_2491_6897 5.354286e+00
R33061 n0_2491_6897 n0_2679_6897 1.074286e+00
R33062 n0_2679_6897 n0_3616_6897 5.354286e+00
R33063 n0_3616_6897 n0_3804_6897 1.074286e+00
R33064 n0_3804_6897 n0_4741_6897 5.354286e+00
R33065 n0_4741_6897 n0_4929_6897 1.074286e+00
R33066 n0_4929_6897 n0_5866_6897 5.354286e+00
R33067 n0_5866_6897 n0_6054_6897 1.074286e+00
R33068 n0_6054_6897 n0_8116_6897 1.178286e+01
R33069 n0_8116_6897 n0_8208_6897 5.257143e-01
R33070 n0_8208_6897 n0_8304_6897 5.485714e-01
R33071 n0_8304_6897 n0_8396_6897 5.257143e-01
R33072 n0_8396_6897 n0_10366_6897 1.125714e+01
R33073 n0_10366_6897 n0_10458_6897 5.257143e-01
R33074 n0_10458_6897 n0_10554_6897 5.485714e-01
R33075 n0_10554_6897 n0_10646_6897 5.257143e-01
R33076 n0_10646_6897 n0_12616_6897 1.125714e+01
R33077 n0_12616_6897 n0_12708_6897 5.257143e-01
R33078 n0_12708_6897 n0_12804_6897 5.485714e-01
R33079 n0_12804_6897 n0_12896_6897 5.257143e-01
R33080 n0_12896_6897 n0_14866_6897 1.125714e+01
R33081 n0_14866_6897 n0_15054_6897 1.074286e+00
R33082 n0_15054_6897 n0_15991_6897 5.354286e+00
R33083 n0_15991_6897 n0_16179_6897 1.074286e+00
R33084 n0_16179_6897 n0_17116_6897 5.354286e+00
R33085 n0_17116_6897 n0_17304_6897 1.074286e+00
R33086 n0_17304_6897 n0_18241_6897 5.354286e+00
R33087 n0_18241_6897 n0_18429_6897 1.074286e+00
R33088 n0_18429_6897 n0_19366_6897 5.354286e+00
R33089 n0_19366_6897 n0_19554_6897 1.074286e+00
R33090 n0_19554_6897 n0_20491_6897 5.354286e+00
R33091 n0_20491_6897 n0_20679_6897 1.074286e+00
R33092 n0_241_6930 n0_429_6930 1.074286e+00
R33093 n0_429_6930 n0_1366_6930 5.354286e+00
R33094 n0_1366_6930 n0_1554_6930 1.074286e+00
R33095 n0_1554_6930 n0_2491_6930 5.354286e+00
R33096 n0_2491_6930 n0_2679_6930 1.074286e+00
R33097 n0_2679_6930 n0_3616_6930 5.354286e+00
R33098 n0_3616_6930 n0_3804_6930 1.074286e+00
R33099 n0_3804_6930 n0_4741_6930 5.354286e+00
R33100 n0_4741_6930 n0_4929_6930 1.074286e+00
R33101 n0_4929_6930 n0_5866_6930 5.354286e+00
R33102 n0_5866_6930 n0_6054_6930 1.074286e+00
R33103 n0_6054_6930 n0_8116_6930 1.178286e+01
R33104 n0_8116_6930 n0_8208_6930 5.257143e-01
R33105 n0_8208_6930 n0_8304_6930 5.485714e-01
R33106 n0_8304_6930 n0_8396_6930 5.257143e-01
R33107 n0_8396_6930 n0_10366_6930 1.125714e+01
R33108 n0_10366_6930 n0_10458_6930 5.257143e-01
R33109 n0_10458_6930 n0_10554_6930 5.485714e-01
R33110 n0_10554_6930 n0_10646_6930 5.257143e-01
R33111 n0_10646_6930 n0_12616_6930 1.125714e+01
R33112 n0_12616_6930 n0_12708_6930 5.257143e-01
R33113 n0_12708_6930 n0_12804_6930 5.485714e-01
R33114 n0_12804_6930 n0_12896_6930 5.257143e-01
R33115 n0_12896_6930 n0_14866_6930 1.125714e+01
R33116 n0_14866_6930 n0_15054_6930 1.074286e+00
R33117 n0_15054_6930 n0_15991_6930 5.354286e+00
R33118 n0_15991_6930 n0_16179_6930 1.074286e+00
R33119 n0_16179_6930 n0_17116_6930 5.354286e+00
R33120 n0_17116_6930 n0_17304_6930 1.074286e+00
R33121 n0_17304_6930 n0_18241_6930 5.354286e+00
R33122 n0_18241_6930 n0_18429_6930 1.074286e+00
R33123 n0_18429_6930 n0_19366_6930 5.354286e+00
R33124 n0_19366_6930 n0_19554_6930 1.074286e+00
R33125 n0_19554_6930 n0_20491_6930 5.354286e+00
R33126 n0_20491_6930 n0_20679_6930 1.074286e+00
R33127 n0_241_7113 n0_429_7113 1.074286e+00
R33128 n0_429_7113 n0_1366_7113 5.354286e+00
R33129 n0_1366_7113 n0_1554_7113 1.074286e+00
R33130 n0_1554_7113 n0_2491_7113 5.354286e+00
R33131 n0_2491_7113 n0_2679_7113 1.074286e+00
R33132 n0_2679_7113 n0_3616_7113 5.354286e+00
R33133 n0_3616_7113 n0_3804_7113 1.074286e+00
R33134 n0_3804_7113 n0_4741_7113 5.354286e+00
R33135 n0_4741_7113 n0_4929_7113 1.074286e+00
R33136 n0_4929_7113 n0_5866_7113 5.354286e+00
R33137 n0_5866_7113 n0_6054_7113 1.074286e+00
R33138 n0_6054_7113 n0_8116_7113 1.178286e+01
R33139 n0_8116_7113 n0_8208_7113 5.257143e-01
R33140 n0_8208_7113 n0_8304_7113 5.485714e-01
R33141 n0_8304_7113 n0_8396_7113 5.257143e-01
R33142 n0_8396_7113 n0_10366_7113 1.125714e+01
R33143 n0_10366_7113 n0_10458_7113 5.257143e-01
R33144 n0_10458_7113 n0_10554_7113 5.485714e-01
R33145 n0_10554_7113 n0_10646_7113 5.257143e-01
R33146 n0_10646_7113 n0_12616_7113 1.125714e+01
R33147 n0_12616_7113 n0_12708_7113 5.257143e-01
R33148 n0_12708_7113 n0_12804_7113 5.485714e-01
R33149 n0_12804_7113 n0_12896_7113 5.257143e-01
R33150 n0_12896_7113 n0_14866_7113 1.125714e+01
R33151 n0_14866_7113 n0_15054_7113 1.074286e+00
R33152 n0_15054_7113 n0_15991_7113 5.354286e+00
R33153 n0_15991_7113 n0_16179_7113 1.074286e+00
R33154 n0_16179_7113 n0_17116_7113 5.354286e+00
R33155 n0_17116_7113 n0_17304_7113 1.074286e+00
R33156 n0_17304_7113 n0_18241_7113 5.354286e+00
R33157 n0_18241_7113 n0_18429_7113 1.074286e+00
R33158 n0_18429_7113 n0_19366_7113 5.354286e+00
R33159 n0_19366_7113 n0_19554_7113 1.074286e+00
R33160 n0_19554_7113 n0_20491_7113 5.354286e+00
R33161 n0_20491_7113 n0_20679_7113 1.074286e+00
R33162 n0_241_7146 n0_1366_7146 6.428571e+00
R33163 n0_1366_7146 n0_2491_7146 6.428571e+00
R33164 n0_2491_7146 n0_3616_7146 6.428571e+00
R33165 n0_3616_7146 n0_4741_7146 6.428571e+00
R33166 n0_4741_7146 n0_5866_7146 6.428571e+00
R33167 n0_5866_7146 n0_8116_7146 1.285714e+01
R33168 n0_8116_7146 n0_8208_7146 5.257143e-01
R33169 n0_8208_7146 n0_8255_7146 2.685714e-01
R33170 n0_8255_7146 n0_8304_7146 2.800000e-01
R33171 n0_8304_7146 n0_8396_7146 5.257143e-01
R33172 n0_8396_7146 n0_10366_7146 1.125714e+01
R33173 n0_10366_7146 n0_10458_7146 5.257143e-01
R33174 n0_10458_7146 n0_10505_7146 2.685714e-01
R33175 n0_10505_7146 n0_10554_7146 2.800000e-01
R33176 n0_10554_7146 n0_10646_7146 5.257143e-01
R33177 n0_10646_7146 n0_12616_7146 1.125714e+01
R33178 n0_12616_7146 n0_12708_7146 5.257143e-01
R33179 n0_12708_7146 n0_12755_7146 2.685714e-01
R33180 n0_12755_7146 n0_12804_7146 2.800000e-01
R33181 n0_12804_7146 n0_12896_7146 5.257143e-01
R33182 n0_12896_7146 n0_14866_7146 1.125714e+01
R33183 n0_14866_7146 n0_15991_7146 6.428571e+00
R33184 n0_15991_7146 n0_17116_7146 6.428571e+00
R33185 n0_17116_7146 n0_18241_7146 6.428571e+00
R33186 n0_18241_7146 n0_19366_7146 6.428571e+00
R33187 n0_19366_7146 n0_20491_7146 6.428571e+00
R33188 n0_241_7329 n0_429_7329 1.074286e+00
R33189 n0_429_7329 n0_1366_7329 5.354286e+00
R33190 n0_1366_7329 n0_1554_7329 1.074286e+00
R33191 n0_1554_7329 n0_2491_7329 5.354286e+00
R33192 n0_2491_7329 n0_2679_7329 1.074286e+00
R33193 n0_2679_7329 n0_3616_7329 5.354286e+00
R33194 n0_3616_7329 n0_3804_7329 1.074286e+00
R33195 n0_3804_7329 n0_4741_7329 5.354286e+00
R33196 n0_4741_7329 n0_4929_7329 1.074286e+00
R33197 n0_4929_7329 n0_5866_7329 5.354286e+00
R33198 n0_5866_7329 n0_6054_7329 1.074286e+00
R33199 n0_6054_7329 n0_6991_7329 5.354286e+00
R33200 n0_6991_7329 n0_7179_7329 1.074286e+00
R33201 n0_7179_7329 n0_8116_7329 5.354286e+00
R33202 n0_8116_7329 n0_8208_7329 5.257143e-01
R33203 n0_8208_7329 n0_8304_7329 5.485714e-01
R33204 n0_8304_7329 n0_8396_7329 5.257143e-01
R33205 n0_8396_7329 n0_10366_7329 1.125714e+01
R33206 n0_10366_7329 n0_10458_7329 5.257143e-01
R33207 n0_10458_7329 n0_10554_7329 5.485714e-01
R33208 n0_10554_7329 n0_10646_7329 5.257143e-01
R33209 n0_10646_7329 n0_12616_7329 1.125714e+01
R33210 n0_12616_7329 n0_12708_7329 5.257143e-01
R33211 n0_12708_7329 n0_12804_7329 5.485714e-01
R33212 n0_12804_7329 n0_12896_7329 5.257143e-01
R33213 n0_12896_7329 n0_13741_7329 4.828571e+00
R33214 n0_13741_7329 n0_13929_7329 1.074286e+00
R33215 n0_13929_7329 n0_14866_7329 5.354286e+00
R33216 n0_14866_7329 n0_15054_7329 1.074286e+00
R33217 n0_15054_7329 n0_15991_7329 5.354286e+00
R33218 n0_15991_7329 n0_16179_7329 1.074286e+00
R33219 n0_16179_7329 n0_17116_7329 5.354286e+00
R33220 n0_17116_7329 n0_17304_7329 1.074286e+00
R33221 n0_17304_7329 n0_18241_7329 5.354286e+00
R33222 n0_18241_7329 n0_18429_7329 1.074286e+00
R33223 n0_18429_7329 n0_19366_7329 5.354286e+00
R33224 n0_19366_7329 n0_19554_7329 1.074286e+00
R33225 n0_19554_7329 n0_20491_7329 5.354286e+00
R33226 n0_20491_7329 n0_20679_7329 1.074286e+00
R33227 n0_241_7362 n0_429_7362 1.074286e+00
R33228 n0_429_7362 n0_1366_7362 5.354286e+00
R33229 n0_1366_7362 n0_1554_7362 1.074286e+00
R33230 n0_1554_7362 n0_2491_7362 5.354286e+00
R33231 n0_2491_7362 n0_2679_7362 1.074286e+00
R33232 n0_2679_7362 n0_3616_7362 5.354286e+00
R33233 n0_3616_7362 n0_3804_7362 1.074286e+00
R33234 n0_3804_7362 n0_4741_7362 5.354286e+00
R33235 n0_4741_7362 n0_4929_7362 1.074286e+00
R33236 n0_4929_7362 n0_5866_7362 5.354286e+00
R33237 n0_5866_7362 n0_6054_7362 1.074286e+00
R33238 n0_6054_7362 n0_6991_7362 5.354286e+00
R33239 n0_6991_7362 n0_7179_7362 1.074286e+00
R33240 n0_7179_7362 n0_8116_7362 5.354286e+00
R33241 n0_8116_7362 n0_8208_7362 5.257143e-01
R33242 n0_8208_7362 n0_8304_7362 5.485714e-01
R33243 n0_8304_7362 n0_8396_7362 5.257143e-01
R33244 n0_8396_7362 n0_10366_7362 1.125714e+01
R33245 n0_10366_7362 n0_10458_7362 5.257143e-01
R33246 n0_10458_7362 n0_10554_7362 5.485714e-01
R33247 n0_10554_7362 n0_10646_7362 5.257143e-01
R33248 n0_10646_7362 n0_12616_7362 1.125714e+01
R33249 n0_12616_7362 n0_12708_7362 5.257143e-01
R33250 n0_12708_7362 n0_12804_7362 5.485714e-01
R33251 n0_12804_7362 n0_12896_7362 5.257143e-01
R33252 n0_12896_7362 n0_13741_7362 4.828571e+00
R33253 n0_13741_7362 n0_13929_7362 1.074286e+00
R33254 n0_13929_7362 n0_14866_7362 5.354286e+00
R33255 n0_14866_7362 n0_15054_7362 1.074286e+00
R33256 n0_15054_7362 n0_15991_7362 5.354286e+00
R33257 n0_15991_7362 n0_16179_7362 1.074286e+00
R33258 n0_16179_7362 n0_17116_7362 5.354286e+00
R33259 n0_17116_7362 n0_17304_7362 1.074286e+00
R33260 n0_17304_7362 n0_18241_7362 5.354286e+00
R33261 n0_18241_7362 n0_18429_7362 1.074286e+00
R33262 n0_18429_7362 n0_19366_7362 5.354286e+00
R33263 n0_19366_7362 n0_19554_7362 1.074286e+00
R33264 n0_19554_7362 n0_20491_7362 5.354286e+00
R33265 n0_20491_7362 n0_20679_7362 1.074286e+00
R33266 n0_241_7545 n0_429_7545 1.074286e+00
R33267 n0_429_7545 n0_1366_7545 5.354286e+00
R33268 n0_1366_7545 n0_1554_7545 1.074286e+00
R33269 n0_1554_7545 n0_2491_7545 5.354286e+00
R33270 n0_2491_7545 n0_2679_7545 1.074286e+00
R33271 n0_2679_7545 n0_3616_7545 5.354286e+00
R33272 n0_3616_7545 n0_3804_7545 1.074286e+00
R33273 n0_3804_7545 n0_4741_7545 5.354286e+00
R33274 n0_4741_7545 n0_4929_7545 1.074286e+00
R33275 n0_4929_7545 n0_5866_7545 5.354286e+00
R33276 n0_5866_7545 n0_6054_7545 1.074286e+00
R33277 n0_6054_7545 n0_6991_7545 5.354286e+00
R33278 n0_6991_7545 n0_7179_7545 1.074286e+00
R33279 n0_7179_7545 n0_8116_7545 5.354286e+00
R33280 n0_8116_7545 n0_8208_7545 5.257143e-01
R33281 n0_8208_7545 n0_8304_7545 5.485714e-01
R33282 n0_8304_7545 n0_8396_7545 5.257143e-01
R33283 n0_8396_7545 n0_10366_7545 1.125714e+01
R33284 n0_10366_7545 n0_10458_7545 5.257143e-01
R33285 n0_10458_7545 n0_10554_7545 5.485714e-01
R33286 n0_10554_7545 n0_10646_7545 5.257143e-01
R33287 n0_10646_7545 n0_12616_7545 1.125714e+01
R33288 n0_12616_7545 n0_12708_7545 5.257143e-01
R33289 n0_12708_7545 n0_12804_7545 5.485714e-01
R33290 n0_12804_7545 n0_12896_7545 5.257143e-01
R33291 n0_12896_7545 n0_13741_7545 4.828571e+00
R33292 n0_13741_7545 n0_13929_7545 1.074286e+00
R33293 n0_13929_7545 n0_14866_7545 5.354286e+00
R33294 n0_14866_7545 n0_15054_7545 1.074286e+00
R33295 n0_15054_7545 n0_15991_7545 5.354286e+00
R33296 n0_15991_7545 n0_16179_7545 1.074286e+00
R33297 n0_16179_7545 n0_17116_7545 5.354286e+00
R33298 n0_17116_7545 n0_17304_7545 1.074286e+00
R33299 n0_17304_7545 n0_18241_7545 5.354286e+00
R33300 n0_18241_7545 n0_18429_7545 1.074286e+00
R33301 n0_18429_7545 n0_19366_7545 5.354286e+00
R33302 n0_19366_7545 n0_19554_7545 1.074286e+00
R33303 n0_19554_7545 n0_20491_7545 5.354286e+00
R33304 n0_20491_7545 n0_20679_7545 1.074286e+00
R33305 n0_241_7578 n0_429_7578 1.074286e+00
R33306 n0_429_7578 n0_1366_7578 5.354286e+00
R33307 n0_1366_7578 n0_1554_7578 1.074286e+00
R33308 n0_1554_7578 n0_2491_7578 5.354286e+00
R33309 n0_2491_7578 n0_2679_7578 1.074286e+00
R33310 n0_2679_7578 n0_3616_7578 5.354286e+00
R33311 n0_3616_7578 n0_3804_7578 1.074286e+00
R33312 n0_3804_7578 n0_4741_7578 5.354286e+00
R33313 n0_4741_7578 n0_4929_7578 1.074286e+00
R33314 n0_4929_7578 n0_5866_7578 5.354286e+00
R33315 n0_5866_7578 n0_6054_7578 1.074286e+00
R33316 n0_6054_7578 n0_6991_7578 5.354286e+00
R33317 n0_6991_7578 n0_7179_7578 1.074286e+00
R33318 n0_7179_7578 n0_8116_7578 5.354286e+00
R33319 n0_8116_7578 n0_8208_7578 5.257143e-01
R33320 n0_8208_7578 n0_8304_7578 5.485714e-01
R33321 n0_8304_7578 n0_8396_7578 5.257143e-01
R33322 n0_8396_7578 n0_10366_7578 1.125714e+01
R33323 n0_10366_7578 n0_10458_7578 5.257143e-01
R33324 n0_10458_7578 n0_10554_7578 5.485714e-01
R33325 n0_10554_7578 n0_10646_7578 5.257143e-01
R33326 n0_10646_7578 n0_12616_7578 1.125714e+01
R33327 n0_12616_7578 n0_12708_7578 5.257143e-01
R33328 n0_12708_7578 n0_12804_7578 5.485714e-01
R33329 n0_12804_7578 n0_12896_7578 5.257143e-01
R33330 n0_12896_7578 n0_13741_7578 4.828571e+00
R33331 n0_13741_7578 n0_13929_7578 1.074286e+00
R33332 n0_13929_7578 n0_14866_7578 5.354286e+00
R33333 n0_14866_7578 n0_15054_7578 1.074286e+00
R33334 n0_15054_7578 n0_15991_7578 5.354286e+00
R33335 n0_15991_7578 n0_16179_7578 1.074286e+00
R33336 n0_16179_7578 n0_17116_7578 5.354286e+00
R33337 n0_17116_7578 n0_17304_7578 1.074286e+00
R33338 n0_17304_7578 n0_18241_7578 5.354286e+00
R33339 n0_18241_7578 n0_18429_7578 1.074286e+00
R33340 n0_18429_7578 n0_19366_7578 5.354286e+00
R33341 n0_19366_7578 n0_19554_7578 1.074286e+00
R33342 n0_19554_7578 n0_20491_7578 5.354286e+00
R33343 n0_20491_7578 n0_20679_7578 1.074286e+00
R33344 n0_241_7761 n0_429_7761 1.074286e+00
R33345 n0_429_7761 n0_1366_7761 5.354286e+00
R33346 n0_1366_7761 n0_1554_7761 1.074286e+00
R33347 n0_1554_7761 n0_2491_7761 5.354286e+00
R33348 n0_2491_7761 n0_2679_7761 1.074286e+00
R33349 n0_2679_7761 n0_3616_7761 5.354286e+00
R33350 n0_3616_7761 n0_3804_7761 1.074286e+00
R33351 n0_3804_7761 n0_4741_7761 5.354286e+00
R33352 n0_4741_7761 n0_4929_7761 1.074286e+00
R33353 n0_4929_7761 n0_5866_7761 5.354286e+00
R33354 n0_5866_7761 n0_6054_7761 1.074286e+00
R33355 n0_6054_7761 n0_6991_7761 5.354286e+00
R33356 n0_6991_7761 n0_7179_7761 1.074286e+00
R33357 n0_7179_7761 n0_8116_7761 5.354286e+00
R33358 n0_8116_7761 n0_8208_7761 5.257143e-01
R33359 n0_8208_7761 n0_8304_7761 5.485714e-01
R33360 n0_8304_7761 n0_8396_7761 5.257143e-01
R33361 n0_8396_7761 n0_10366_7761 1.125714e+01
R33362 n0_10366_7761 n0_10458_7761 5.257143e-01
R33363 n0_10458_7761 n0_10554_7761 5.485714e-01
R33364 n0_10554_7761 n0_10646_7761 5.257143e-01
R33365 n0_10646_7761 n0_12616_7761 1.125714e+01
R33366 n0_12616_7761 n0_12708_7761 5.257143e-01
R33367 n0_12708_7761 n0_12804_7761 5.485714e-01
R33368 n0_12804_7761 n0_12896_7761 5.257143e-01
R33369 n0_12896_7761 n0_13741_7761 4.828571e+00
R33370 n0_13741_7761 n0_13929_7761 1.074286e+00
R33371 n0_13929_7761 n0_14866_7761 5.354286e+00
R33372 n0_14866_7761 n0_15054_7761 1.074286e+00
R33373 n0_15054_7761 n0_15991_7761 5.354286e+00
R33374 n0_15991_7761 n0_16179_7761 1.074286e+00
R33375 n0_16179_7761 n0_17116_7761 5.354286e+00
R33376 n0_17116_7761 n0_17304_7761 1.074286e+00
R33377 n0_17304_7761 n0_18241_7761 5.354286e+00
R33378 n0_18241_7761 n0_18429_7761 1.074286e+00
R33379 n0_18429_7761 n0_19366_7761 5.354286e+00
R33380 n0_19366_7761 n0_19554_7761 1.074286e+00
R33381 n0_19554_7761 n0_20491_7761 5.354286e+00
R33382 n0_20491_7761 n0_20679_7761 1.074286e+00
R33383 n0_241_7794 n0_429_7794 1.074286e+00
R33384 n0_429_7794 n0_1366_7794 5.354286e+00
R33385 n0_1366_7794 n0_1554_7794 1.074286e+00
R33386 n0_1554_7794 n0_2491_7794 5.354286e+00
R33387 n0_2491_7794 n0_2679_7794 1.074286e+00
R33388 n0_2679_7794 n0_3616_7794 5.354286e+00
R33389 n0_3616_7794 n0_3804_7794 1.074286e+00
R33390 n0_3804_7794 n0_4741_7794 5.354286e+00
R33391 n0_4741_7794 n0_4929_7794 1.074286e+00
R33392 n0_4929_7794 n0_5866_7794 5.354286e+00
R33393 n0_5866_7794 n0_6054_7794 1.074286e+00
R33394 n0_6054_7794 n0_6991_7794 5.354286e+00
R33395 n0_6991_7794 n0_7179_7794 1.074286e+00
R33396 n0_7179_7794 n0_8116_7794 5.354286e+00
R33397 n0_8116_7794 n0_8208_7794 5.257143e-01
R33398 n0_8208_7794 n0_8304_7794 5.485714e-01
R33399 n0_8304_7794 n0_8396_7794 5.257143e-01
R33400 n0_8396_7794 n0_10366_7794 1.125714e+01
R33401 n0_10366_7794 n0_10458_7794 5.257143e-01
R33402 n0_10458_7794 n0_10554_7794 5.485714e-01
R33403 n0_10554_7794 n0_10646_7794 5.257143e-01
R33404 n0_10646_7794 n0_12616_7794 1.125714e+01
R33405 n0_12616_7794 n0_12708_7794 5.257143e-01
R33406 n0_12708_7794 n0_12804_7794 5.485714e-01
R33407 n0_12804_7794 n0_12896_7794 5.257143e-01
R33408 n0_12896_7794 n0_13741_7794 4.828571e+00
R33409 n0_13741_7794 n0_13929_7794 1.074286e+00
R33410 n0_13929_7794 n0_14866_7794 5.354286e+00
R33411 n0_14866_7794 n0_15054_7794 1.074286e+00
R33412 n0_15054_7794 n0_15991_7794 5.354286e+00
R33413 n0_15991_7794 n0_16179_7794 1.074286e+00
R33414 n0_16179_7794 n0_17116_7794 5.354286e+00
R33415 n0_17116_7794 n0_17304_7794 1.074286e+00
R33416 n0_17304_7794 n0_18241_7794 5.354286e+00
R33417 n0_18241_7794 n0_18429_7794 1.074286e+00
R33418 n0_18429_7794 n0_19366_7794 5.354286e+00
R33419 n0_19366_7794 n0_19554_7794 1.074286e+00
R33420 n0_19554_7794 n0_20491_7794 5.354286e+00
R33421 n0_20491_7794 n0_20679_7794 1.074286e+00
R33422 n0_241_7977 n0_429_7977 1.074286e+00
R33423 n0_429_7977 n0_1366_7977 5.354286e+00
R33424 n0_1366_7977 n0_1554_7977 1.074286e+00
R33425 n0_1554_7977 n0_2491_7977 5.354286e+00
R33426 n0_2491_7977 n0_2679_7977 1.074286e+00
R33427 n0_2679_7977 n0_3616_7977 5.354286e+00
R33428 n0_3616_7977 n0_3804_7977 1.074286e+00
R33429 n0_3804_7977 n0_4741_7977 5.354286e+00
R33430 n0_4741_7977 n0_4929_7977 1.074286e+00
R33431 n0_4929_7977 n0_5866_7977 5.354286e+00
R33432 n0_5866_7977 n0_6054_7977 1.074286e+00
R33433 n0_6054_7977 n0_6991_7977 5.354286e+00
R33434 n0_6991_7977 n0_7179_7977 1.074286e+00
R33435 n0_7179_7977 n0_8116_7977 5.354286e+00
R33436 n0_8116_7977 n0_8208_7977 5.257143e-01
R33437 n0_8208_7977 n0_8304_7977 5.485714e-01
R33438 n0_8304_7977 n0_8396_7977 5.257143e-01
R33439 n0_8396_7977 n0_10366_7977 1.125714e+01
R33440 n0_10366_7977 n0_10458_7977 5.257143e-01
R33441 n0_10458_7977 n0_10554_7977 5.485714e-01
R33442 n0_10554_7977 n0_10646_7977 5.257143e-01
R33443 n0_10646_7977 n0_12616_7977 1.125714e+01
R33444 n0_12616_7977 n0_12708_7977 5.257143e-01
R33445 n0_12708_7977 n0_12804_7977 5.485714e-01
R33446 n0_12804_7977 n0_12896_7977 5.257143e-01
R33447 n0_12896_7977 n0_13741_7977 4.828571e+00
R33448 n0_13741_7977 n0_13929_7977 1.074286e+00
R33449 n0_13929_7977 n0_14866_7977 5.354286e+00
R33450 n0_14866_7977 n0_15054_7977 1.074286e+00
R33451 n0_15054_7977 n0_15991_7977 5.354286e+00
R33452 n0_15991_7977 n0_16179_7977 1.074286e+00
R33453 n0_16179_7977 n0_17116_7977 5.354286e+00
R33454 n0_17116_7977 n0_17304_7977 1.074286e+00
R33455 n0_17304_7977 n0_18241_7977 5.354286e+00
R33456 n0_18241_7977 n0_18429_7977 1.074286e+00
R33457 n0_18429_7977 n0_19366_7977 5.354286e+00
R33458 n0_19366_7977 n0_19554_7977 1.074286e+00
R33459 n0_19554_7977 n0_20491_7977 5.354286e+00
R33460 n0_20491_7977 n0_20679_7977 1.074286e+00
R33461 n0_241_8010 n0_429_8010 1.074286e+00
R33462 n0_429_8010 n0_1366_8010 5.354286e+00
R33463 n0_1366_8010 n0_1554_8010 1.074286e+00
R33464 n0_1554_8010 n0_2491_8010 5.354286e+00
R33465 n0_2491_8010 n0_2679_8010 1.074286e+00
R33466 n0_2679_8010 n0_3616_8010 5.354286e+00
R33467 n0_3616_8010 n0_3804_8010 1.074286e+00
R33468 n0_3804_8010 n0_4741_8010 5.354286e+00
R33469 n0_4741_8010 n0_4929_8010 1.074286e+00
R33470 n0_4929_8010 n0_5866_8010 5.354286e+00
R33471 n0_5866_8010 n0_6054_8010 1.074286e+00
R33472 n0_6054_8010 n0_6991_8010 5.354286e+00
R33473 n0_6991_8010 n0_7179_8010 1.074286e+00
R33474 n0_7179_8010 n0_8116_8010 5.354286e+00
R33475 n0_8116_8010 n0_8208_8010 5.257143e-01
R33476 n0_8208_8010 n0_8304_8010 5.485714e-01
R33477 n0_8304_8010 n0_8396_8010 5.257143e-01
R33478 n0_8396_8010 n0_10366_8010 1.125714e+01
R33479 n0_10366_8010 n0_10458_8010 5.257143e-01
R33480 n0_10458_8010 n0_10554_8010 5.485714e-01
R33481 n0_10554_8010 n0_10646_8010 5.257143e-01
R33482 n0_10646_8010 n0_12616_8010 1.125714e+01
R33483 n0_12616_8010 n0_12708_8010 5.257143e-01
R33484 n0_12708_8010 n0_12804_8010 5.485714e-01
R33485 n0_12804_8010 n0_12896_8010 5.257143e-01
R33486 n0_12896_8010 n0_13741_8010 4.828571e+00
R33487 n0_13741_8010 n0_13929_8010 1.074286e+00
R33488 n0_13929_8010 n0_14866_8010 5.354286e+00
R33489 n0_14866_8010 n0_15054_8010 1.074286e+00
R33490 n0_15054_8010 n0_15991_8010 5.354286e+00
R33491 n0_15991_8010 n0_16179_8010 1.074286e+00
R33492 n0_16179_8010 n0_17116_8010 5.354286e+00
R33493 n0_17116_8010 n0_17304_8010 1.074286e+00
R33494 n0_17304_8010 n0_18241_8010 5.354286e+00
R33495 n0_18241_8010 n0_18429_8010 1.074286e+00
R33496 n0_18429_8010 n0_19366_8010 5.354286e+00
R33497 n0_19366_8010 n0_19554_8010 1.074286e+00
R33498 n0_19554_8010 n0_20491_8010 5.354286e+00
R33499 n0_20491_8010 n0_20679_8010 1.074286e+00
R33500 n0_241_8193 n0_429_8193 1.074286e+00
R33501 n0_429_8193 n0_1366_8193 5.354286e+00
R33502 n0_1366_8193 n0_1554_8193 1.074286e+00
R33503 n0_1554_8193 n0_2491_8193 5.354286e+00
R33504 n0_2491_8193 n0_2679_8193 1.074286e+00
R33505 n0_2679_8193 n0_3616_8193 5.354286e+00
R33506 n0_3616_8193 n0_3804_8193 1.074286e+00
R33507 n0_3804_8193 n0_4741_8193 5.354286e+00
R33508 n0_4741_8193 n0_4929_8193 1.074286e+00
R33509 n0_4929_8193 n0_5866_8193 5.354286e+00
R33510 n0_5866_8193 n0_6054_8193 1.074286e+00
R33511 n0_6054_8193 n0_6991_8193 5.354286e+00
R33512 n0_6991_8193 n0_7179_8193 1.074286e+00
R33513 n0_7179_8193 n0_8116_8193 5.354286e+00
R33514 n0_8116_8193 n0_8208_8193 5.257143e-01
R33515 n0_8208_8193 n0_8304_8193 5.485714e-01
R33516 n0_8304_8193 n0_8396_8193 5.257143e-01
R33517 n0_8396_8193 n0_10366_8193 1.125714e+01
R33518 n0_10366_8193 n0_10458_8193 5.257143e-01
R33519 n0_10458_8193 n0_10554_8193 5.485714e-01
R33520 n0_10554_8193 n0_10646_8193 5.257143e-01
R33521 n0_10646_8193 n0_12616_8193 1.125714e+01
R33522 n0_12616_8193 n0_12708_8193 5.257143e-01
R33523 n0_12708_8193 n0_12804_8193 5.485714e-01
R33524 n0_12804_8193 n0_12896_8193 5.257143e-01
R33525 n0_12896_8193 n0_13741_8193 4.828571e+00
R33526 n0_13741_8193 n0_13929_8193 1.074286e+00
R33527 n0_13929_8193 n0_14866_8193 5.354286e+00
R33528 n0_14866_8193 n0_15054_8193 1.074286e+00
R33529 n0_15054_8193 n0_15991_8193 5.354286e+00
R33530 n0_15991_8193 n0_16179_8193 1.074286e+00
R33531 n0_16179_8193 n0_17116_8193 5.354286e+00
R33532 n0_17116_8193 n0_17304_8193 1.074286e+00
R33533 n0_17304_8193 n0_18241_8193 5.354286e+00
R33534 n0_18241_8193 n0_18429_8193 1.074286e+00
R33535 n0_18429_8193 n0_19366_8193 5.354286e+00
R33536 n0_19366_8193 n0_19554_8193 1.074286e+00
R33537 n0_19554_8193 n0_20491_8193 5.354286e+00
R33538 n0_20491_8193 n0_20679_8193 1.074286e+00
R33539 n0_241_8226 n0_429_8226 1.074286e+00
R33540 n0_429_8226 n0_1366_8226 5.354286e+00
R33541 n0_1366_8226 n0_1554_8226 1.074286e+00
R33542 n0_1554_8226 n0_2491_8226 5.354286e+00
R33543 n0_2491_8226 n0_2679_8226 1.074286e+00
R33544 n0_2679_8226 n0_3616_8226 5.354286e+00
R33545 n0_3616_8226 n0_3804_8226 1.074286e+00
R33546 n0_3804_8226 n0_4741_8226 5.354286e+00
R33547 n0_4741_8226 n0_4929_8226 1.074286e+00
R33548 n0_4929_8226 n0_5866_8226 5.354286e+00
R33549 n0_5866_8226 n0_6054_8226 1.074286e+00
R33550 n0_6054_8226 n0_6991_8226 5.354286e+00
R33551 n0_6991_8226 n0_7179_8226 1.074286e+00
R33552 n0_7179_8226 n0_8116_8226 5.354286e+00
R33553 n0_8116_8226 n0_8208_8226 5.257143e-01
R33554 n0_8208_8226 n0_8304_8226 5.485714e-01
R33555 n0_8304_8226 n0_8396_8226 5.257143e-01
R33556 n0_8396_8226 n0_10366_8226 1.125714e+01
R33557 n0_10366_8226 n0_10458_8226 5.257143e-01
R33558 n0_10458_8226 n0_10554_8226 5.485714e-01
R33559 n0_10554_8226 n0_10646_8226 5.257143e-01
R33560 n0_10646_8226 n0_12616_8226 1.125714e+01
R33561 n0_12616_8226 n0_12708_8226 5.257143e-01
R33562 n0_12708_8226 n0_12804_8226 5.485714e-01
R33563 n0_12804_8226 n0_12896_8226 5.257143e-01
R33564 n0_12896_8226 n0_13741_8226 4.828571e+00
R33565 n0_13741_8226 n0_13929_8226 1.074286e+00
R33566 n0_13929_8226 n0_14866_8226 5.354286e+00
R33567 n0_14866_8226 n0_15054_8226 1.074286e+00
R33568 n0_15054_8226 n0_15991_8226 5.354286e+00
R33569 n0_15991_8226 n0_16179_8226 1.074286e+00
R33570 n0_16179_8226 n0_17116_8226 5.354286e+00
R33571 n0_17116_8226 n0_17304_8226 1.074286e+00
R33572 n0_17304_8226 n0_18241_8226 5.354286e+00
R33573 n0_18241_8226 n0_18429_8226 1.074286e+00
R33574 n0_18429_8226 n0_19366_8226 5.354286e+00
R33575 n0_19366_8226 n0_19554_8226 1.074286e+00
R33576 n0_19554_8226 n0_20491_8226 5.354286e+00
R33577 n0_20491_8226 n0_20679_8226 1.074286e+00
R33578 n0_241_8409 n0_380_8409 7.942857e-01
R33579 n0_380_8409 n0_429_8409 2.800000e-01
R33580 n0_429_8409 n0_1366_8409 5.354286e+00
R33581 n0_1366_8409 n0_1505_8409 7.942857e-01
R33582 n0_1505_8409 n0_1554_8409 2.800000e-01
R33583 n0_1554_8409 n0_2491_8409 5.354286e+00
R33584 n0_2491_8409 n0_2630_8409 7.942857e-01
R33585 n0_2630_8409 n0_2679_8409 2.800000e-01
R33586 n0_2679_8409 n0_3616_8409 5.354286e+00
R33587 n0_3616_8409 n0_3755_8409 7.942857e-01
R33588 n0_3755_8409 n0_3804_8409 2.800000e-01
R33589 n0_3804_8409 n0_4741_8409 5.354286e+00
R33590 n0_4741_8409 n0_4880_8409 7.942857e-01
R33591 n0_4880_8409 n0_4929_8409 2.800000e-01
R33592 n0_4929_8409 n0_5866_8409 5.354286e+00
R33593 n0_5866_8409 n0_6005_8409 7.942857e-01
R33594 n0_6005_8409 n0_6054_8409 2.800000e-01
R33595 n0_6054_8409 n0_6991_8409 5.354286e+00
R33596 n0_6991_8409 n0_7130_8409 7.942857e-01
R33597 n0_7130_8409 n0_7179_8409 2.800000e-01
R33598 n0_7179_8409 n0_8116_8409 5.354286e+00
R33599 n0_8116_8409 n0_8208_8409 5.257143e-01
R33600 n0_8208_8409 n0_8255_8409 2.685714e-01
R33601 n0_8255_8409 n0_8304_8409 2.800000e-01
R33602 n0_8304_8409 n0_10366_8409 1.178286e+01
R33603 n0_10366_8409 n0_10458_8409 5.257143e-01
R33604 n0_10458_8409 n0_10505_8409 2.685714e-01
R33605 n0_10505_8409 n0_10554_8409 2.800000e-01
R33606 n0_10554_8409 n0_10646_8409 5.257143e-01
R33607 n0_10646_8409 n0_12616_8409 1.125714e+01
R33608 n0_12616_8409 n0_12708_8409 5.257143e-01
R33609 n0_12708_8409 n0_12755_8409 2.685714e-01
R33610 n0_12755_8409 n0_12804_8409 2.800000e-01
R33611 n0_12804_8409 n0_13741_8409 5.354286e+00
R33612 n0_13741_8409 n0_13880_8409 7.942857e-01
R33613 n0_13880_8409 n0_13929_8409 2.800000e-01
R33614 n0_13929_8409 n0_14866_8409 5.354286e+00
R33615 n0_14866_8409 n0_15005_8409 7.942857e-01
R33616 n0_15005_8409 n0_15054_8409 2.800000e-01
R33617 n0_15054_8409 n0_15991_8409 5.354286e+00
R33618 n0_15991_8409 n0_16130_8409 7.942857e-01
R33619 n0_16130_8409 n0_16179_8409 2.800000e-01
R33620 n0_16179_8409 n0_17116_8409 5.354286e+00
R33621 n0_17116_8409 n0_17255_8409 7.942857e-01
R33622 n0_17255_8409 n0_17304_8409 2.800000e-01
R33623 n0_17304_8409 n0_18241_8409 5.354286e+00
R33624 n0_18241_8409 n0_18380_8409 7.942857e-01
R33625 n0_18380_8409 n0_18429_8409 2.800000e-01
R33626 n0_18429_8409 n0_19366_8409 5.354286e+00
R33627 n0_19366_8409 n0_19505_8409 7.942857e-01
R33628 n0_19505_8409 n0_19554_8409 2.800000e-01
R33629 n0_19554_8409 n0_20491_8409 5.354286e+00
R33630 n0_20491_8409 n0_20630_8409 7.942857e-01
R33631 n0_20630_8409 n0_20679_8409 2.800000e-01
R33632 n0_241_8442 n0_429_8442 1.074286e+00
R33633 n0_429_8442 n0_1366_8442 5.354286e+00
R33634 n0_1366_8442 n0_1554_8442 1.074286e+00
R33635 n0_1554_8442 n0_2491_8442 5.354286e+00
R33636 n0_2491_8442 n0_2679_8442 1.074286e+00
R33637 n0_2679_8442 n0_3616_8442 5.354286e+00
R33638 n0_3616_8442 n0_3804_8442 1.074286e+00
R33639 n0_3804_8442 n0_4741_8442 5.354286e+00
R33640 n0_4741_8442 n0_4929_8442 1.074286e+00
R33641 n0_4929_8442 n0_5866_8442 5.354286e+00
R33642 n0_5866_8442 n0_6054_8442 1.074286e+00
R33643 n0_6054_8442 n0_6991_8442 5.354286e+00
R33644 n0_6991_8442 n0_7179_8442 1.074286e+00
R33645 n0_7179_8442 n0_8116_8442 5.354286e+00
R33646 n0_8116_8442 n0_8208_8442 5.257143e-01
R33647 n0_8208_8442 n0_8304_8442 5.485714e-01
R33648 n0_8304_8442 n0_10366_8442 1.178286e+01
R33649 n0_10366_8442 n0_10458_8442 5.257143e-01
R33650 n0_10458_8442 n0_10554_8442 5.485714e-01
R33651 n0_10554_8442 n0_10646_8442 5.257143e-01
R33652 n0_10646_8442 n0_12616_8442 1.125714e+01
R33653 n0_12616_8442 n0_12708_8442 5.257143e-01
R33654 n0_12708_8442 n0_12804_8442 5.485714e-01
R33655 n0_12804_8442 n0_13741_8442 5.354286e+00
R33656 n0_13741_8442 n0_13929_8442 1.074286e+00
R33657 n0_13929_8442 n0_14866_8442 5.354286e+00
R33658 n0_14866_8442 n0_15054_8442 1.074286e+00
R33659 n0_15054_8442 n0_15991_8442 5.354286e+00
R33660 n0_15991_8442 n0_16179_8442 1.074286e+00
R33661 n0_16179_8442 n0_17116_8442 5.354286e+00
R33662 n0_17116_8442 n0_17304_8442 1.074286e+00
R33663 n0_17304_8442 n0_18241_8442 5.354286e+00
R33664 n0_18241_8442 n0_18429_8442 1.074286e+00
R33665 n0_18429_8442 n0_19366_8442 5.354286e+00
R33666 n0_19366_8442 n0_19554_8442 1.074286e+00
R33667 n0_19554_8442 n0_20491_8442 5.354286e+00
R33668 n0_20491_8442 n0_20679_8442 1.074286e+00
R33669 n0_241_8625 n0_429_8625 1.074286e+00
R33670 n0_429_8625 n0_1366_8625 5.354286e+00
R33671 n0_1366_8625 n0_1554_8625 1.074286e+00
R33672 n0_1554_8625 n0_2491_8625 5.354286e+00
R33673 n0_2491_8625 n0_2679_8625 1.074286e+00
R33674 n0_2679_8625 n0_3616_8625 5.354286e+00
R33675 n0_3616_8625 n0_3804_8625 1.074286e+00
R33676 n0_3804_8625 n0_4741_8625 5.354286e+00
R33677 n0_4741_8625 n0_4929_8625 1.074286e+00
R33678 n0_4929_8625 n0_5866_8625 5.354286e+00
R33679 n0_5866_8625 n0_6054_8625 1.074286e+00
R33680 n0_6054_8625 n0_6991_8625 5.354286e+00
R33681 n0_6991_8625 n0_7179_8625 1.074286e+00
R33682 n0_7179_8625 n0_8116_8625 5.354286e+00
R33683 n0_8116_8625 n0_8304_8625 1.074286e+00
R33684 n0_8304_8625 n0_10366_8625 1.178286e+01
R33685 n0_10366_8625 n0_10458_8625 5.257143e-01
R33686 n0_10458_8625 n0_10554_8625 5.485714e-01
R33687 n0_10554_8625 n0_10646_8625 5.257143e-01
R33688 n0_10646_8625 n0_12616_8625 1.125714e+01
R33689 n0_12616_8625 n0_12804_8625 1.074286e+00
R33690 n0_12804_8625 n0_13741_8625 5.354286e+00
R33691 n0_13741_8625 n0_13929_8625 1.074286e+00
R33692 n0_13929_8625 n0_14866_8625 5.354286e+00
R33693 n0_14866_8625 n0_15054_8625 1.074286e+00
R33694 n0_15054_8625 n0_15991_8625 5.354286e+00
R33695 n0_15991_8625 n0_16179_8625 1.074286e+00
R33696 n0_16179_8625 n0_17116_8625 5.354286e+00
R33697 n0_17116_8625 n0_17304_8625 1.074286e+00
R33698 n0_17304_8625 n0_18241_8625 5.354286e+00
R33699 n0_18241_8625 n0_18429_8625 1.074286e+00
R33700 n0_18429_8625 n0_19366_8625 5.354286e+00
R33701 n0_19366_8625 n0_19554_8625 1.074286e+00
R33702 n0_19554_8625 n0_20491_8625 5.354286e+00
R33703 n0_20491_8625 n0_20679_8625 1.074286e+00
R33704 n0_241_8658 n0_429_8658 1.074286e+00
R33705 n0_429_8658 n0_1366_8658 5.354286e+00
R33706 n0_1366_8658 n0_1554_8658 1.074286e+00
R33707 n0_1554_8658 n0_2491_8658 5.354286e+00
R33708 n0_2491_8658 n0_2679_8658 1.074286e+00
R33709 n0_2679_8658 n0_3616_8658 5.354286e+00
R33710 n0_3616_8658 n0_3804_8658 1.074286e+00
R33711 n0_3804_8658 n0_4741_8658 5.354286e+00
R33712 n0_4741_8658 n0_4929_8658 1.074286e+00
R33713 n0_4929_8658 n0_5866_8658 5.354286e+00
R33714 n0_5866_8658 n0_6054_8658 1.074286e+00
R33715 n0_6054_8658 n0_6991_8658 5.354286e+00
R33716 n0_6991_8658 n0_7179_8658 1.074286e+00
R33717 n0_7179_8658 n0_8116_8658 5.354286e+00
R33718 n0_8116_8658 n0_8304_8658 1.074286e+00
R33719 n0_8304_8658 n0_10366_8658 1.178286e+01
R33720 n0_10366_8658 n0_10458_8658 5.257143e-01
R33721 n0_10458_8658 n0_10554_8658 5.485714e-01
R33722 n0_10554_8658 n0_10646_8658 5.257143e-01
R33723 n0_10646_8658 n0_12616_8658 1.125714e+01
R33724 n0_12616_8658 n0_12804_8658 1.074286e+00
R33725 n0_12804_8658 n0_13741_8658 5.354286e+00
R33726 n0_13741_8658 n0_13929_8658 1.074286e+00
R33727 n0_13929_8658 n0_14866_8658 5.354286e+00
R33728 n0_14866_8658 n0_15054_8658 1.074286e+00
R33729 n0_15054_8658 n0_15991_8658 5.354286e+00
R33730 n0_15991_8658 n0_16179_8658 1.074286e+00
R33731 n0_16179_8658 n0_17116_8658 5.354286e+00
R33732 n0_17116_8658 n0_17304_8658 1.074286e+00
R33733 n0_17304_8658 n0_18241_8658 5.354286e+00
R33734 n0_18241_8658 n0_18429_8658 1.074286e+00
R33735 n0_18429_8658 n0_19366_8658 5.354286e+00
R33736 n0_19366_8658 n0_19554_8658 1.074286e+00
R33737 n0_19554_8658 n0_20491_8658 5.354286e+00
R33738 n0_20491_8658 n0_20679_8658 1.074286e+00
R33739 n0_241_8841 n0_429_8841 1.074286e+00
R33740 n0_429_8841 n0_1366_8841 5.354286e+00
R33741 n0_1366_8841 n0_1554_8841 1.074286e+00
R33742 n0_1554_8841 n0_2491_8841 5.354286e+00
R33743 n0_2491_8841 n0_2679_8841 1.074286e+00
R33744 n0_2679_8841 n0_3616_8841 5.354286e+00
R33745 n0_3616_8841 n0_3804_8841 1.074286e+00
R33746 n0_3804_8841 n0_4741_8841 5.354286e+00
R33747 n0_4741_8841 n0_4929_8841 1.074286e+00
R33748 n0_4929_8841 n0_5866_8841 5.354286e+00
R33749 n0_5866_8841 n0_6054_8841 1.074286e+00
R33750 n0_6054_8841 n0_6991_8841 5.354286e+00
R33751 n0_6991_8841 n0_7179_8841 1.074286e+00
R33752 n0_7179_8841 n0_8116_8841 5.354286e+00
R33753 n0_8116_8841 n0_8304_8841 1.074286e+00
R33754 n0_8304_8841 n0_10366_8841 1.178286e+01
R33755 n0_10366_8841 n0_10458_8841 5.257143e-01
R33756 n0_10458_8841 n0_10554_8841 5.485714e-01
R33757 n0_10554_8841 n0_10646_8841 5.257143e-01
R33758 n0_10646_8841 n0_12616_8841 1.125714e+01
R33759 n0_12616_8841 n0_12804_8841 1.074286e+00
R33760 n0_12804_8841 n0_13741_8841 5.354286e+00
R33761 n0_13741_8841 n0_13929_8841 1.074286e+00
R33762 n0_13929_8841 n0_14866_8841 5.354286e+00
R33763 n0_14866_8841 n0_15054_8841 1.074286e+00
R33764 n0_15054_8841 n0_15991_8841 5.354286e+00
R33765 n0_15991_8841 n0_16179_8841 1.074286e+00
R33766 n0_16179_8841 n0_17116_8841 5.354286e+00
R33767 n0_17116_8841 n0_17304_8841 1.074286e+00
R33768 n0_17304_8841 n0_18241_8841 5.354286e+00
R33769 n0_18241_8841 n0_18429_8841 1.074286e+00
R33770 n0_18429_8841 n0_19366_8841 5.354286e+00
R33771 n0_19366_8841 n0_19554_8841 1.074286e+00
R33772 n0_19554_8841 n0_20491_8841 5.354286e+00
R33773 n0_20491_8841 n0_20679_8841 1.074286e+00
R33774 n0_241_8874 n0_429_8874 1.074286e+00
R33775 n0_429_8874 n0_1366_8874 5.354286e+00
R33776 n0_1366_8874 n0_1554_8874 1.074286e+00
R33777 n0_1554_8874 n0_2491_8874 5.354286e+00
R33778 n0_2491_8874 n0_2679_8874 1.074286e+00
R33779 n0_2679_8874 n0_3616_8874 5.354286e+00
R33780 n0_3616_8874 n0_3804_8874 1.074286e+00
R33781 n0_3804_8874 n0_4741_8874 5.354286e+00
R33782 n0_4741_8874 n0_4929_8874 1.074286e+00
R33783 n0_4929_8874 n0_5866_8874 5.354286e+00
R33784 n0_5866_8874 n0_6054_8874 1.074286e+00
R33785 n0_6054_8874 n0_6991_8874 5.354286e+00
R33786 n0_6991_8874 n0_7179_8874 1.074286e+00
R33787 n0_7179_8874 n0_8116_8874 5.354286e+00
R33788 n0_8116_8874 n0_8304_8874 1.074286e+00
R33789 n0_8304_8874 n0_10366_8874 1.178286e+01
R33790 n0_10366_8874 n0_10458_8874 5.257143e-01
R33791 n0_10458_8874 n0_10554_8874 5.485714e-01
R33792 n0_10554_8874 n0_10646_8874 5.257143e-01
R33793 n0_10646_8874 n0_12616_8874 1.125714e+01
R33794 n0_12616_8874 n0_12804_8874 1.074286e+00
R33795 n0_12804_8874 n0_13741_8874 5.354286e+00
R33796 n0_13741_8874 n0_13929_8874 1.074286e+00
R33797 n0_13929_8874 n0_14866_8874 5.354286e+00
R33798 n0_14866_8874 n0_15054_8874 1.074286e+00
R33799 n0_15054_8874 n0_15991_8874 5.354286e+00
R33800 n0_15991_8874 n0_16179_8874 1.074286e+00
R33801 n0_16179_8874 n0_17116_8874 5.354286e+00
R33802 n0_17116_8874 n0_17304_8874 1.074286e+00
R33803 n0_17304_8874 n0_18241_8874 5.354286e+00
R33804 n0_18241_8874 n0_18429_8874 1.074286e+00
R33805 n0_18429_8874 n0_19366_8874 5.354286e+00
R33806 n0_19366_8874 n0_19554_8874 1.074286e+00
R33807 n0_19554_8874 n0_20491_8874 5.354286e+00
R33808 n0_20491_8874 n0_20679_8874 1.074286e+00
R33809 n0_241_9057 n0_429_9057 1.074286e+00
R33810 n0_429_9057 n0_1366_9057 5.354286e+00
R33811 n0_1366_9057 n0_1554_9057 1.074286e+00
R33812 n0_1554_9057 n0_2491_9057 5.354286e+00
R33813 n0_2491_9057 n0_2679_9057 1.074286e+00
R33814 n0_2679_9057 n0_3616_9057 5.354286e+00
R33815 n0_3616_9057 n0_3804_9057 1.074286e+00
R33816 n0_3804_9057 n0_4741_9057 5.354286e+00
R33817 n0_4741_9057 n0_4929_9057 1.074286e+00
R33818 n0_4929_9057 n0_5866_9057 5.354286e+00
R33819 n0_5866_9057 n0_6054_9057 1.074286e+00
R33820 n0_6054_9057 n0_6991_9057 5.354286e+00
R33821 n0_6991_9057 n0_7179_9057 1.074286e+00
R33822 n0_7179_9057 n0_8116_9057 5.354286e+00
R33823 n0_8116_9057 n0_8304_9057 1.074286e+00
R33824 n0_8304_9057 n0_10366_9057 1.178286e+01
R33825 n0_10366_9057 n0_10458_9057 5.257143e-01
R33826 n0_10458_9057 n0_10554_9057 5.485714e-01
R33827 n0_10554_9057 n0_10646_9057 5.257143e-01
R33828 n0_10646_9057 n0_12616_9057 1.125714e+01
R33829 n0_12616_9057 n0_12804_9057 1.074286e+00
R33830 n0_12804_9057 n0_13741_9057 5.354286e+00
R33831 n0_13741_9057 n0_13929_9057 1.074286e+00
R33832 n0_13929_9057 n0_14866_9057 5.354286e+00
R33833 n0_14866_9057 n0_15054_9057 1.074286e+00
R33834 n0_15054_9057 n0_15991_9057 5.354286e+00
R33835 n0_15991_9057 n0_16179_9057 1.074286e+00
R33836 n0_16179_9057 n0_17116_9057 5.354286e+00
R33837 n0_17116_9057 n0_17304_9057 1.074286e+00
R33838 n0_17304_9057 n0_18241_9057 5.354286e+00
R33839 n0_18241_9057 n0_18429_9057 1.074286e+00
R33840 n0_18429_9057 n0_19366_9057 5.354286e+00
R33841 n0_19366_9057 n0_19554_9057 1.074286e+00
R33842 n0_19554_9057 n0_20491_9057 5.354286e+00
R33843 n0_20491_9057 n0_20679_9057 1.074286e+00
R33844 n0_241_9090 n0_429_9090 1.074286e+00
R33845 n0_429_9090 n0_1366_9090 5.354286e+00
R33846 n0_1366_9090 n0_1554_9090 1.074286e+00
R33847 n0_1554_9090 n0_2491_9090 5.354286e+00
R33848 n0_2491_9090 n0_2679_9090 1.074286e+00
R33849 n0_2679_9090 n0_3616_9090 5.354286e+00
R33850 n0_3616_9090 n0_3804_9090 1.074286e+00
R33851 n0_3804_9090 n0_4741_9090 5.354286e+00
R33852 n0_4741_9090 n0_4929_9090 1.074286e+00
R33853 n0_4929_9090 n0_5866_9090 5.354286e+00
R33854 n0_5866_9090 n0_6054_9090 1.074286e+00
R33855 n0_6054_9090 n0_6991_9090 5.354286e+00
R33856 n0_6991_9090 n0_7179_9090 1.074286e+00
R33857 n0_7179_9090 n0_8116_9090 5.354286e+00
R33858 n0_8116_9090 n0_8304_9090 1.074286e+00
R33859 n0_8304_9090 n0_10366_9090 1.178286e+01
R33860 n0_10366_9090 n0_10458_9090 5.257143e-01
R33861 n0_10458_9090 n0_10554_9090 5.485714e-01
R33862 n0_10554_9090 n0_10646_9090 5.257143e-01
R33863 n0_10646_9090 n0_12616_9090 1.125714e+01
R33864 n0_12616_9090 n0_12804_9090 1.074286e+00
R33865 n0_12804_9090 n0_13741_9090 5.354286e+00
R33866 n0_13741_9090 n0_13929_9090 1.074286e+00
R33867 n0_13929_9090 n0_14866_9090 5.354286e+00
R33868 n0_14866_9090 n0_15054_9090 1.074286e+00
R33869 n0_15054_9090 n0_15991_9090 5.354286e+00
R33870 n0_15991_9090 n0_16179_9090 1.074286e+00
R33871 n0_16179_9090 n0_17116_9090 5.354286e+00
R33872 n0_17116_9090 n0_17304_9090 1.074286e+00
R33873 n0_17304_9090 n0_18241_9090 5.354286e+00
R33874 n0_18241_9090 n0_18429_9090 1.074286e+00
R33875 n0_18429_9090 n0_19366_9090 5.354286e+00
R33876 n0_19366_9090 n0_19554_9090 1.074286e+00
R33877 n0_19554_9090 n0_20491_9090 5.354286e+00
R33878 n0_20491_9090 n0_20679_9090 1.074286e+00
R33879 n0_241_12081 n0_429_12081 1.074286e+00
R33880 n0_429_12081 n0_1366_12081 5.354286e+00
R33881 n0_1366_12081 n0_1554_12081 1.074286e+00
R33882 n0_1554_12081 n0_2491_12081 5.354286e+00
R33883 n0_2491_12081 n0_2679_12081 1.074286e+00
R33884 n0_2679_12081 n0_3616_12081 5.354286e+00
R33885 n0_3616_12081 n0_3804_12081 1.074286e+00
R33886 n0_3804_12081 n0_4741_12081 5.354286e+00
R33887 n0_4741_12081 n0_4929_12081 1.074286e+00
R33888 n0_4929_12081 n0_5866_12081 5.354286e+00
R33889 n0_5866_12081 n0_6054_12081 1.074286e+00
R33890 n0_6054_12081 n0_6991_12081 5.354286e+00
R33891 n0_6991_12081 n0_7179_12081 1.074286e+00
R33892 n0_7179_12081 n0_8116_12081 5.354286e+00
R33893 n0_8116_12081 n0_8304_12081 1.074286e+00
R33894 n0_8304_12081 n0_10366_12081 1.178286e+01
R33895 n0_10366_12081 n0_10458_12081 5.257143e-01
R33896 n0_10458_12081 n0_10554_12081 5.485714e-01
R33897 n0_10554_12081 n0_10646_12081 5.257143e-01
R33898 n0_10646_12081 n0_12616_12081 1.125714e+01
R33899 n0_12616_12081 n0_12804_12081 1.074286e+00
R33900 n0_12804_12081 n0_13741_12081 5.354286e+00
R33901 n0_13741_12081 n0_13929_12081 1.074286e+00
R33902 n0_13929_12081 n0_14866_12081 5.354286e+00
R33903 n0_14866_12081 n0_15054_12081 1.074286e+00
R33904 n0_15054_12081 n0_15991_12081 5.354286e+00
R33905 n0_15991_12081 n0_16179_12081 1.074286e+00
R33906 n0_16179_12081 n0_17116_12081 5.354286e+00
R33907 n0_17116_12081 n0_17304_12081 1.074286e+00
R33908 n0_17304_12081 n0_18241_12081 5.354286e+00
R33909 n0_18241_12081 n0_18429_12081 1.074286e+00
R33910 n0_18429_12081 n0_19366_12081 5.354286e+00
R33911 n0_19366_12081 n0_19554_12081 1.074286e+00
R33912 n0_19554_12081 n0_20491_12081 5.354286e+00
R33913 n0_20491_12081 n0_20679_12081 1.074286e+00
R33914 n0_241_12114 n0_429_12114 1.074286e+00
R33915 n0_429_12114 n0_1366_12114 5.354286e+00
R33916 n0_1366_12114 n0_1554_12114 1.074286e+00
R33917 n0_1554_12114 n0_2491_12114 5.354286e+00
R33918 n0_2491_12114 n0_2679_12114 1.074286e+00
R33919 n0_2679_12114 n0_3616_12114 5.354286e+00
R33920 n0_3616_12114 n0_3804_12114 1.074286e+00
R33921 n0_3804_12114 n0_4741_12114 5.354286e+00
R33922 n0_4741_12114 n0_4929_12114 1.074286e+00
R33923 n0_4929_12114 n0_5866_12114 5.354286e+00
R33924 n0_5866_12114 n0_6054_12114 1.074286e+00
R33925 n0_6054_12114 n0_6991_12114 5.354286e+00
R33926 n0_6991_12114 n0_7179_12114 1.074286e+00
R33927 n0_7179_12114 n0_8116_12114 5.354286e+00
R33928 n0_8116_12114 n0_8304_12114 1.074286e+00
R33929 n0_8304_12114 n0_10366_12114 1.178286e+01
R33930 n0_10366_12114 n0_10458_12114 5.257143e-01
R33931 n0_10458_12114 n0_10554_12114 5.485714e-01
R33932 n0_10554_12114 n0_10646_12114 5.257143e-01
R33933 n0_10646_12114 n0_12616_12114 1.125714e+01
R33934 n0_12616_12114 n0_12804_12114 1.074286e+00
R33935 n0_12804_12114 n0_13741_12114 5.354286e+00
R33936 n0_13741_12114 n0_13929_12114 1.074286e+00
R33937 n0_13929_12114 n0_14866_12114 5.354286e+00
R33938 n0_14866_12114 n0_15054_12114 1.074286e+00
R33939 n0_15054_12114 n0_15991_12114 5.354286e+00
R33940 n0_15991_12114 n0_16179_12114 1.074286e+00
R33941 n0_16179_12114 n0_17116_12114 5.354286e+00
R33942 n0_17116_12114 n0_17304_12114 1.074286e+00
R33943 n0_17304_12114 n0_18241_12114 5.354286e+00
R33944 n0_18241_12114 n0_18429_12114 1.074286e+00
R33945 n0_18429_12114 n0_19366_12114 5.354286e+00
R33946 n0_19366_12114 n0_19554_12114 1.074286e+00
R33947 n0_19554_12114 n0_20491_12114 5.354286e+00
R33948 n0_20491_12114 n0_20679_12114 1.074286e+00
R33949 n0_241_12297 n0_429_12297 1.074286e+00
R33950 n0_429_12297 n0_1366_12297 5.354286e+00
R33951 n0_1366_12297 n0_1554_12297 1.074286e+00
R33952 n0_1554_12297 n0_2491_12297 5.354286e+00
R33953 n0_2491_12297 n0_2679_12297 1.074286e+00
R33954 n0_2679_12297 n0_3616_12297 5.354286e+00
R33955 n0_3616_12297 n0_3804_12297 1.074286e+00
R33956 n0_3804_12297 n0_4741_12297 5.354286e+00
R33957 n0_4741_12297 n0_4929_12297 1.074286e+00
R33958 n0_4929_12297 n0_5866_12297 5.354286e+00
R33959 n0_5866_12297 n0_6054_12297 1.074286e+00
R33960 n0_6054_12297 n0_6991_12297 5.354286e+00
R33961 n0_6991_12297 n0_7179_12297 1.074286e+00
R33962 n0_7179_12297 n0_8116_12297 5.354286e+00
R33963 n0_8116_12297 n0_8304_12297 1.074286e+00
R33964 n0_8304_12297 n0_10366_12297 1.178286e+01
R33965 n0_10366_12297 n0_10458_12297 5.257143e-01
R33966 n0_10458_12297 n0_10554_12297 5.485714e-01
R33967 n0_10554_12297 n0_10646_12297 5.257143e-01
R33968 n0_10646_12297 n0_12616_12297 1.125714e+01
R33969 n0_12616_12297 n0_12804_12297 1.074286e+00
R33970 n0_12804_12297 n0_13741_12297 5.354286e+00
R33971 n0_13741_12297 n0_13929_12297 1.074286e+00
R33972 n0_13929_12297 n0_14866_12297 5.354286e+00
R33973 n0_14866_12297 n0_15054_12297 1.074286e+00
R33974 n0_15054_12297 n0_15991_12297 5.354286e+00
R33975 n0_15991_12297 n0_16179_12297 1.074286e+00
R33976 n0_16179_12297 n0_17116_12297 5.354286e+00
R33977 n0_17116_12297 n0_17304_12297 1.074286e+00
R33978 n0_17304_12297 n0_18241_12297 5.354286e+00
R33979 n0_18241_12297 n0_18429_12297 1.074286e+00
R33980 n0_18429_12297 n0_19366_12297 5.354286e+00
R33981 n0_19366_12297 n0_19554_12297 1.074286e+00
R33982 n0_19554_12297 n0_20491_12297 5.354286e+00
R33983 n0_20491_12297 n0_20679_12297 1.074286e+00
R33984 n0_241_12330 n0_429_12330 1.074286e+00
R33985 n0_429_12330 n0_1366_12330 5.354286e+00
R33986 n0_1366_12330 n0_1554_12330 1.074286e+00
R33987 n0_1554_12330 n0_2491_12330 5.354286e+00
R33988 n0_2491_12330 n0_2679_12330 1.074286e+00
R33989 n0_2679_12330 n0_3616_12330 5.354286e+00
R33990 n0_3616_12330 n0_3804_12330 1.074286e+00
R33991 n0_3804_12330 n0_4741_12330 5.354286e+00
R33992 n0_4741_12330 n0_4929_12330 1.074286e+00
R33993 n0_4929_12330 n0_5866_12330 5.354286e+00
R33994 n0_5866_12330 n0_6054_12330 1.074286e+00
R33995 n0_6054_12330 n0_6991_12330 5.354286e+00
R33996 n0_6991_12330 n0_7179_12330 1.074286e+00
R33997 n0_7179_12330 n0_8116_12330 5.354286e+00
R33998 n0_8116_12330 n0_8304_12330 1.074286e+00
R33999 n0_8304_12330 n0_10366_12330 1.178286e+01
R34000 n0_10366_12330 n0_10458_12330 5.257143e-01
R34001 n0_10458_12330 n0_10554_12330 5.485714e-01
R34002 n0_10554_12330 n0_10646_12330 5.257143e-01
R34003 n0_10646_12330 n0_12616_12330 1.125714e+01
R34004 n0_12616_12330 n0_12804_12330 1.074286e+00
R34005 n0_12804_12330 n0_13741_12330 5.354286e+00
R34006 n0_13741_12330 n0_13929_12330 1.074286e+00
R34007 n0_13929_12330 n0_14866_12330 5.354286e+00
R34008 n0_14866_12330 n0_15054_12330 1.074286e+00
R34009 n0_15054_12330 n0_15991_12330 5.354286e+00
R34010 n0_15991_12330 n0_16179_12330 1.074286e+00
R34011 n0_16179_12330 n0_17116_12330 5.354286e+00
R34012 n0_17116_12330 n0_17304_12330 1.074286e+00
R34013 n0_17304_12330 n0_18241_12330 5.354286e+00
R34014 n0_18241_12330 n0_18429_12330 1.074286e+00
R34015 n0_18429_12330 n0_19366_12330 5.354286e+00
R34016 n0_19366_12330 n0_19554_12330 1.074286e+00
R34017 n0_19554_12330 n0_20491_12330 5.354286e+00
R34018 n0_20491_12330 n0_20679_12330 1.074286e+00
R34019 n0_241_12513 n0_429_12513 1.074286e+00
R34020 n0_429_12513 n0_1366_12513 5.354286e+00
R34021 n0_1366_12513 n0_1554_12513 1.074286e+00
R34022 n0_1554_12513 n0_2491_12513 5.354286e+00
R34023 n0_2491_12513 n0_2679_12513 1.074286e+00
R34024 n0_2679_12513 n0_3616_12513 5.354286e+00
R34025 n0_3616_12513 n0_3804_12513 1.074286e+00
R34026 n0_3804_12513 n0_4741_12513 5.354286e+00
R34027 n0_4741_12513 n0_4929_12513 1.074286e+00
R34028 n0_4929_12513 n0_5866_12513 5.354286e+00
R34029 n0_5866_12513 n0_6054_12513 1.074286e+00
R34030 n0_6054_12513 n0_6991_12513 5.354286e+00
R34031 n0_6991_12513 n0_7179_12513 1.074286e+00
R34032 n0_7179_12513 n0_8116_12513 5.354286e+00
R34033 n0_8116_12513 n0_8304_12513 1.074286e+00
R34034 n0_8304_12513 n0_10366_12513 1.178286e+01
R34035 n0_10366_12513 n0_10458_12513 5.257143e-01
R34036 n0_10458_12513 n0_10554_12513 5.485714e-01
R34037 n0_10554_12513 n0_10646_12513 5.257143e-01
R34038 n0_10646_12513 n0_12616_12513 1.125714e+01
R34039 n0_12616_12513 n0_12804_12513 1.074286e+00
R34040 n0_12804_12513 n0_13741_12513 5.354286e+00
R34041 n0_13741_12513 n0_13929_12513 1.074286e+00
R34042 n0_13929_12513 n0_14866_12513 5.354286e+00
R34043 n0_14866_12513 n0_15054_12513 1.074286e+00
R34044 n0_15054_12513 n0_15991_12513 5.354286e+00
R34045 n0_15991_12513 n0_16179_12513 1.074286e+00
R34046 n0_16179_12513 n0_17116_12513 5.354286e+00
R34047 n0_17116_12513 n0_17304_12513 1.074286e+00
R34048 n0_17304_12513 n0_18241_12513 5.354286e+00
R34049 n0_18241_12513 n0_18429_12513 1.074286e+00
R34050 n0_18429_12513 n0_19366_12513 5.354286e+00
R34051 n0_19366_12513 n0_19554_12513 1.074286e+00
R34052 n0_19554_12513 n0_20491_12513 5.354286e+00
R34053 n0_20491_12513 n0_20679_12513 1.074286e+00
R34054 n0_241_12546 n0_429_12546 1.074286e+00
R34055 n0_429_12546 n0_1366_12546 5.354286e+00
R34056 n0_1366_12546 n0_1554_12546 1.074286e+00
R34057 n0_1554_12546 n0_2491_12546 5.354286e+00
R34058 n0_2491_12546 n0_2679_12546 1.074286e+00
R34059 n0_2679_12546 n0_3616_12546 5.354286e+00
R34060 n0_3616_12546 n0_3804_12546 1.074286e+00
R34061 n0_3804_12546 n0_4741_12546 5.354286e+00
R34062 n0_4741_12546 n0_4929_12546 1.074286e+00
R34063 n0_4929_12546 n0_5866_12546 5.354286e+00
R34064 n0_5866_12546 n0_6054_12546 1.074286e+00
R34065 n0_6054_12546 n0_6991_12546 5.354286e+00
R34066 n0_6991_12546 n0_7179_12546 1.074286e+00
R34067 n0_7179_12546 n0_8116_12546 5.354286e+00
R34068 n0_8116_12546 n0_8304_12546 1.074286e+00
R34069 n0_8304_12546 n0_10366_12546 1.178286e+01
R34070 n0_10366_12546 n0_10458_12546 5.257143e-01
R34071 n0_10458_12546 n0_10554_12546 5.485714e-01
R34072 n0_10554_12546 n0_10646_12546 5.257143e-01
R34073 n0_10646_12546 n0_12616_12546 1.125714e+01
R34074 n0_12616_12546 n0_12804_12546 1.074286e+00
R34075 n0_12804_12546 n0_13741_12546 5.354286e+00
R34076 n0_13741_12546 n0_13929_12546 1.074286e+00
R34077 n0_13929_12546 n0_14866_12546 5.354286e+00
R34078 n0_14866_12546 n0_15054_12546 1.074286e+00
R34079 n0_15054_12546 n0_15991_12546 5.354286e+00
R34080 n0_15991_12546 n0_16179_12546 1.074286e+00
R34081 n0_16179_12546 n0_17116_12546 5.354286e+00
R34082 n0_17116_12546 n0_17304_12546 1.074286e+00
R34083 n0_17304_12546 n0_18241_12546 5.354286e+00
R34084 n0_18241_12546 n0_18429_12546 1.074286e+00
R34085 n0_18429_12546 n0_19366_12546 5.354286e+00
R34086 n0_19366_12546 n0_19554_12546 1.074286e+00
R34087 n0_19554_12546 n0_20491_12546 5.354286e+00
R34088 n0_20491_12546 n0_20679_12546 1.074286e+00
R34089 n0_241_12729 n0_429_12729 1.074286e+00
R34090 n0_429_12729 n0_1366_12729 5.354286e+00
R34091 n0_1366_12729 n0_1554_12729 1.074286e+00
R34092 n0_1554_12729 n0_2491_12729 5.354286e+00
R34093 n0_2491_12729 n0_2679_12729 1.074286e+00
R34094 n0_2679_12729 n0_3616_12729 5.354286e+00
R34095 n0_3616_12729 n0_3804_12729 1.074286e+00
R34096 n0_3804_12729 n0_4741_12729 5.354286e+00
R34097 n0_4741_12729 n0_4929_12729 1.074286e+00
R34098 n0_4929_12729 n0_5866_12729 5.354286e+00
R34099 n0_5866_12729 n0_6054_12729 1.074286e+00
R34100 n0_6054_12729 n0_6991_12729 5.354286e+00
R34101 n0_6991_12729 n0_7179_12729 1.074286e+00
R34102 n0_7179_12729 n0_8116_12729 5.354286e+00
R34103 n0_8116_12729 n0_8304_12729 1.074286e+00
R34104 n0_8304_12729 n0_10366_12729 1.178286e+01
R34105 n0_10366_12729 n0_10458_12729 5.257143e-01
R34106 n0_10458_12729 n0_10554_12729 5.485714e-01
R34107 n0_10554_12729 n0_10646_12729 5.257143e-01
R34108 n0_10646_12729 n0_12616_12729 1.125714e+01
R34109 n0_12616_12729 n0_12804_12729 1.074286e+00
R34110 n0_12804_12729 n0_13741_12729 5.354286e+00
R34111 n0_13741_12729 n0_13929_12729 1.074286e+00
R34112 n0_13929_12729 n0_14866_12729 5.354286e+00
R34113 n0_14866_12729 n0_15054_12729 1.074286e+00
R34114 n0_15054_12729 n0_15991_12729 5.354286e+00
R34115 n0_15991_12729 n0_16179_12729 1.074286e+00
R34116 n0_16179_12729 n0_17116_12729 5.354286e+00
R34117 n0_17116_12729 n0_17304_12729 1.074286e+00
R34118 n0_17304_12729 n0_18241_12729 5.354286e+00
R34119 n0_18241_12729 n0_18429_12729 1.074286e+00
R34120 n0_18429_12729 n0_19366_12729 5.354286e+00
R34121 n0_19366_12729 n0_19554_12729 1.074286e+00
R34122 n0_19554_12729 n0_20491_12729 5.354286e+00
R34123 n0_20491_12729 n0_20679_12729 1.074286e+00
R34124 n0_241_12762 n0_429_12762 1.074286e+00
R34125 n0_429_12762 n0_1366_12762 5.354286e+00
R34126 n0_1366_12762 n0_1554_12762 1.074286e+00
R34127 n0_1554_12762 n0_2491_12762 5.354286e+00
R34128 n0_2491_12762 n0_2679_12762 1.074286e+00
R34129 n0_2679_12762 n0_3616_12762 5.354286e+00
R34130 n0_3616_12762 n0_3804_12762 1.074286e+00
R34131 n0_3804_12762 n0_4741_12762 5.354286e+00
R34132 n0_4741_12762 n0_4929_12762 1.074286e+00
R34133 n0_4929_12762 n0_5866_12762 5.354286e+00
R34134 n0_5866_12762 n0_6054_12762 1.074286e+00
R34135 n0_6054_12762 n0_6991_12762 5.354286e+00
R34136 n0_6991_12762 n0_7179_12762 1.074286e+00
R34137 n0_7179_12762 n0_8116_12762 5.354286e+00
R34138 n0_8116_12762 n0_8208_12762 5.257143e-01
R34139 n0_8208_12762 n0_8304_12762 5.485714e-01
R34140 n0_8304_12762 n0_10366_12762 1.178286e+01
R34141 n0_10366_12762 n0_10458_12762 5.257143e-01
R34142 n0_10458_12762 n0_10554_12762 5.485714e-01
R34143 n0_10554_12762 n0_10646_12762 5.257143e-01
R34144 n0_10646_12762 n0_12616_12762 1.125714e+01
R34145 n0_12616_12762 n0_12708_12762 5.257143e-01
R34146 n0_12708_12762 n0_12804_12762 5.485714e-01
R34147 n0_12804_12762 n0_13741_12762 5.354286e+00
R34148 n0_13741_12762 n0_13929_12762 1.074286e+00
R34149 n0_13929_12762 n0_14866_12762 5.354286e+00
R34150 n0_14866_12762 n0_15054_12762 1.074286e+00
R34151 n0_15054_12762 n0_15991_12762 5.354286e+00
R34152 n0_15991_12762 n0_16179_12762 1.074286e+00
R34153 n0_16179_12762 n0_17116_12762 5.354286e+00
R34154 n0_17116_12762 n0_17304_12762 1.074286e+00
R34155 n0_17304_12762 n0_18241_12762 5.354286e+00
R34156 n0_18241_12762 n0_18429_12762 1.074286e+00
R34157 n0_18429_12762 n0_19366_12762 5.354286e+00
R34158 n0_19366_12762 n0_19554_12762 1.074286e+00
R34159 n0_19554_12762 n0_20491_12762 5.354286e+00
R34160 n0_20491_12762 n0_20679_12762 1.074286e+00
R34161 n0_241_12945 n0_429_12945 1.074286e+00
R34162 n0_429_12945 n0_1366_12945 5.354286e+00
R34163 n0_1366_12945 n0_1554_12945 1.074286e+00
R34164 n0_1554_12945 n0_2491_12945 5.354286e+00
R34165 n0_2491_12945 n0_2679_12945 1.074286e+00
R34166 n0_2679_12945 n0_3616_12945 5.354286e+00
R34167 n0_3616_12945 n0_3804_12945 1.074286e+00
R34168 n0_3804_12945 n0_4741_12945 5.354286e+00
R34169 n0_4741_12945 n0_4929_12945 1.074286e+00
R34170 n0_4929_12945 n0_5866_12945 5.354286e+00
R34171 n0_5866_12945 n0_6054_12945 1.074286e+00
R34172 n0_6054_12945 n0_6991_12945 5.354286e+00
R34173 n0_6991_12945 n0_7179_12945 1.074286e+00
R34174 n0_7179_12945 n0_8116_12945 5.354286e+00
R34175 n0_8116_12945 n0_8208_12945 5.257143e-01
R34176 n0_8208_12945 n0_8304_12945 5.485714e-01
R34177 n0_8304_12945 n0_8396_12945 5.257143e-01
R34178 n0_8396_12945 n0_10366_12945 1.125714e+01
R34179 n0_10366_12945 n0_10458_12945 5.257143e-01
R34180 n0_10458_12945 n0_10554_12945 5.485714e-01
R34181 n0_10554_12945 n0_10646_12945 5.257143e-01
R34182 n0_10646_12945 n0_12616_12945 1.125714e+01
R34183 n0_12616_12945 n0_12708_12945 5.257143e-01
R34184 n0_12708_12945 n0_12804_12945 5.485714e-01
R34185 n0_12804_12945 n0_12896_12945 5.257143e-01
R34186 n0_12896_12945 n0_13741_12945 4.828571e+00
R34187 n0_13741_12945 n0_13929_12945 1.074286e+00
R34188 n0_13929_12945 n0_14866_12945 5.354286e+00
R34189 n0_14866_12945 n0_15054_12945 1.074286e+00
R34190 n0_15054_12945 n0_15991_12945 5.354286e+00
R34191 n0_15991_12945 n0_16179_12945 1.074286e+00
R34192 n0_16179_12945 n0_17116_12945 5.354286e+00
R34193 n0_17116_12945 n0_17304_12945 1.074286e+00
R34194 n0_17304_12945 n0_18241_12945 5.354286e+00
R34195 n0_18241_12945 n0_18429_12945 1.074286e+00
R34196 n0_18429_12945 n0_19366_12945 5.354286e+00
R34197 n0_19366_12945 n0_19554_12945 1.074286e+00
R34198 n0_19554_12945 n0_20491_12945 5.354286e+00
R34199 n0_20491_12945 n0_20679_12945 1.074286e+00
R34200 n0_241_12978 n0_429_12978 1.074286e+00
R34201 n0_429_12978 n0_1366_12978 5.354286e+00
R34202 n0_1366_12978 n0_1554_12978 1.074286e+00
R34203 n0_1554_12978 n0_2491_12978 5.354286e+00
R34204 n0_2491_12978 n0_2679_12978 1.074286e+00
R34205 n0_2679_12978 n0_3616_12978 5.354286e+00
R34206 n0_3616_12978 n0_3804_12978 1.074286e+00
R34207 n0_3804_12978 n0_4741_12978 5.354286e+00
R34208 n0_4741_12978 n0_4929_12978 1.074286e+00
R34209 n0_4929_12978 n0_5866_12978 5.354286e+00
R34210 n0_5866_12978 n0_6054_12978 1.074286e+00
R34211 n0_6054_12978 n0_6991_12978 5.354286e+00
R34212 n0_6991_12978 n0_7179_12978 1.074286e+00
R34213 n0_7179_12978 n0_8116_12978 5.354286e+00
R34214 n0_8116_12978 n0_8208_12978 5.257143e-01
R34215 n0_8208_12978 n0_8304_12978 5.485714e-01
R34216 n0_8304_12978 n0_8396_12978 5.257143e-01
R34217 n0_8396_12978 n0_10366_12978 1.125714e+01
R34218 n0_10366_12978 n0_10458_12978 5.257143e-01
R34219 n0_10458_12978 n0_10554_12978 5.485714e-01
R34220 n0_10554_12978 n0_10646_12978 5.257143e-01
R34221 n0_10646_12978 n0_12616_12978 1.125714e+01
R34222 n0_12616_12978 n0_12708_12978 5.257143e-01
R34223 n0_12708_12978 n0_12804_12978 5.485714e-01
R34224 n0_12804_12978 n0_12896_12978 5.257143e-01
R34225 n0_12896_12978 n0_13741_12978 4.828571e+00
R34226 n0_13741_12978 n0_13929_12978 1.074286e+00
R34227 n0_13929_12978 n0_14866_12978 5.354286e+00
R34228 n0_14866_12978 n0_15054_12978 1.074286e+00
R34229 n0_15054_12978 n0_15991_12978 5.354286e+00
R34230 n0_15991_12978 n0_16179_12978 1.074286e+00
R34231 n0_16179_12978 n0_17116_12978 5.354286e+00
R34232 n0_17116_12978 n0_17304_12978 1.074286e+00
R34233 n0_17304_12978 n0_18241_12978 5.354286e+00
R34234 n0_18241_12978 n0_18429_12978 1.074286e+00
R34235 n0_18429_12978 n0_19366_12978 5.354286e+00
R34236 n0_19366_12978 n0_19554_12978 1.074286e+00
R34237 n0_19554_12978 n0_20491_12978 5.354286e+00
R34238 n0_20491_12978 n0_20679_12978 1.074286e+00
R34239 n0_241_13161 n0_429_13161 1.074286e+00
R34240 n0_429_13161 n0_1366_13161 5.354286e+00
R34241 n0_1366_13161 n0_1554_13161 1.074286e+00
R34242 n0_1554_13161 n0_2491_13161 5.354286e+00
R34243 n0_2491_13161 n0_2679_13161 1.074286e+00
R34244 n0_2679_13161 n0_3616_13161 5.354286e+00
R34245 n0_3616_13161 n0_3804_13161 1.074286e+00
R34246 n0_3804_13161 n0_4741_13161 5.354286e+00
R34247 n0_4741_13161 n0_4929_13161 1.074286e+00
R34248 n0_4929_13161 n0_5866_13161 5.354286e+00
R34249 n0_5866_13161 n0_6054_13161 1.074286e+00
R34250 n0_6054_13161 n0_6991_13161 5.354286e+00
R34251 n0_6991_13161 n0_7179_13161 1.074286e+00
R34252 n0_7179_13161 n0_8116_13161 5.354286e+00
R34253 n0_8116_13161 n0_8208_13161 5.257143e-01
R34254 n0_8208_13161 n0_8304_13161 5.485714e-01
R34255 n0_8304_13161 n0_8396_13161 5.257143e-01
R34256 n0_8396_13161 n0_10366_13161 1.125714e+01
R34257 n0_10366_13161 n0_10458_13161 5.257143e-01
R34258 n0_10458_13161 n0_10554_13161 5.485714e-01
R34259 n0_10554_13161 n0_10646_13161 5.257143e-01
R34260 n0_10646_13161 n0_12616_13161 1.125714e+01
R34261 n0_12616_13161 n0_12708_13161 5.257143e-01
R34262 n0_12708_13161 n0_12804_13161 5.485714e-01
R34263 n0_12804_13161 n0_12896_13161 5.257143e-01
R34264 n0_12896_13161 n0_13741_13161 4.828571e+00
R34265 n0_13741_13161 n0_13929_13161 1.074286e+00
R34266 n0_13929_13161 n0_14866_13161 5.354286e+00
R34267 n0_14866_13161 n0_15054_13161 1.074286e+00
R34268 n0_15054_13161 n0_15991_13161 5.354286e+00
R34269 n0_15991_13161 n0_16179_13161 1.074286e+00
R34270 n0_16179_13161 n0_17116_13161 5.354286e+00
R34271 n0_17116_13161 n0_17304_13161 1.074286e+00
R34272 n0_17304_13161 n0_18241_13161 5.354286e+00
R34273 n0_18241_13161 n0_18429_13161 1.074286e+00
R34274 n0_18429_13161 n0_19366_13161 5.354286e+00
R34275 n0_19366_13161 n0_19554_13161 1.074286e+00
R34276 n0_19554_13161 n0_20491_13161 5.354286e+00
R34277 n0_20491_13161 n0_20679_13161 1.074286e+00
R34278 n0_241_13194 n0_429_13194 1.074286e+00
R34279 n0_429_13194 n0_1366_13194 5.354286e+00
R34280 n0_1366_13194 n0_1554_13194 1.074286e+00
R34281 n0_1554_13194 n0_2491_13194 5.354286e+00
R34282 n0_2491_13194 n0_2679_13194 1.074286e+00
R34283 n0_2679_13194 n0_3616_13194 5.354286e+00
R34284 n0_3616_13194 n0_3804_13194 1.074286e+00
R34285 n0_3804_13194 n0_4741_13194 5.354286e+00
R34286 n0_4741_13194 n0_4929_13194 1.074286e+00
R34287 n0_4929_13194 n0_5866_13194 5.354286e+00
R34288 n0_5866_13194 n0_6054_13194 1.074286e+00
R34289 n0_6054_13194 n0_6991_13194 5.354286e+00
R34290 n0_6991_13194 n0_7179_13194 1.074286e+00
R34291 n0_7179_13194 n0_8116_13194 5.354286e+00
R34292 n0_8116_13194 n0_8208_13194 5.257143e-01
R34293 n0_8208_13194 n0_8304_13194 5.485714e-01
R34294 n0_8304_13194 n0_8396_13194 5.257143e-01
R34295 n0_8396_13194 n0_10366_13194 1.125714e+01
R34296 n0_10366_13194 n0_10458_13194 5.257143e-01
R34297 n0_10458_13194 n0_10554_13194 5.485714e-01
R34298 n0_10554_13194 n0_10646_13194 5.257143e-01
R34299 n0_10646_13194 n0_12616_13194 1.125714e+01
R34300 n0_12616_13194 n0_12708_13194 5.257143e-01
R34301 n0_12708_13194 n0_12804_13194 5.485714e-01
R34302 n0_12804_13194 n0_12896_13194 5.257143e-01
R34303 n0_12896_13194 n0_13741_13194 4.828571e+00
R34304 n0_13741_13194 n0_13929_13194 1.074286e+00
R34305 n0_13929_13194 n0_14866_13194 5.354286e+00
R34306 n0_14866_13194 n0_15054_13194 1.074286e+00
R34307 n0_15054_13194 n0_15991_13194 5.354286e+00
R34308 n0_15991_13194 n0_16179_13194 1.074286e+00
R34309 n0_16179_13194 n0_17116_13194 5.354286e+00
R34310 n0_17116_13194 n0_17304_13194 1.074286e+00
R34311 n0_17304_13194 n0_18241_13194 5.354286e+00
R34312 n0_18241_13194 n0_18429_13194 1.074286e+00
R34313 n0_18429_13194 n0_19366_13194 5.354286e+00
R34314 n0_19366_13194 n0_19554_13194 1.074286e+00
R34315 n0_19554_13194 n0_20491_13194 5.354286e+00
R34316 n0_20491_13194 n0_20679_13194 1.074286e+00
R34317 n0_241_13377 n0_429_13377 1.074286e+00
R34318 n0_429_13377 n0_1366_13377 5.354286e+00
R34319 n0_1366_13377 n0_1554_13377 1.074286e+00
R34320 n0_1554_13377 n0_2491_13377 5.354286e+00
R34321 n0_2491_13377 n0_2679_13377 1.074286e+00
R34322 n0_2679_13377 n0_3616_13377 5.354286e+00
R34323 n0_3616_13377 n0_3804_13377 1.074286e+00
R34324 n0_3804_13377 n0_4741_13377 5.354286e+00
R34325 n0_4741_13377 n0_4929_13377 1.074286e+00
R34326 n0_4929_13377 n0_5866_13377 5.354286e+00
R34327 n0_5866_13377 n0_6054_13377 1.074286e+00
R34328 n0_6054_13377 n0_6991_13377 5.354286e+00
R34329 n0_6991_13377 n0_7179_13377 1.074286e+00
R34330 n0_7179_13377 n0_8116_13377 5.354286e+00
R34331 n0_8116_13377 n0_8208_13377 5.257143e-01
R34332 n0_8208_13377 n0_8304_13377 5.485714e-01
R34333 n0_8304_13377 n0_8396_13377 5.257143e-01
R34334 n0_8396_13377 n0_10366_13377 1.125714e+01
R34335 n0_10366_13377 n0_10458_13377 5.257143e-01
R34336 n0_10458_13377 n0_10554_13377 5.485714e-01
R34337 n0_10554_13377 n0_10646_13377 5.257143e-01
R34338 n0_10646_13377 n0_12616_13377 1.125714e+01
R34339 n0_12616_13377 n0_12708_13377 5.257143e-01
R34340 n0_12708_13377 n0_12804_13377 5.485714e-01
R34341 n0_12804_13377 n0_12896_13377 5.257143e-01
R34342 n0_12896_13377 n0_13741_13377 4.828571e+00
R34343 n0_13741_13377 n0_13929_13377 1.074286e+00
R34344 n0_13929_13377 n0_14866_13377 5.354286e+00
R34345 n0_14866_13377 n0_15054_13377 1.074286e+00
R34346 n0_15054_13377 n0_15991_13377 5.354286e+00
R34347 n0_15991_13377 n0_16179_13377 1.074286e+00
R34348 n0_16179_13377 n0_17116_13377 5.354286e+00
R34349 n0_17116_13377 n0_17304_13377 1.074286e+00
R34350 n0_17304_13377 n0_18241_13377 5.354286e+00
R34351 n0_18241_13377 n0_18429_13377 1.074286e+00
R34352 n0_18429_13377 n0_19366_13377 5.354286e+00
R34353 n0_19366_13377 n0_19554_13377 1.074286e+00
R34354 n0_19554_13377 n0_20491_13377 5.354286e+00
R34355 n0_20491_13377 n0_20679_13377 1.074286e+00
R34356 n0_241_13410 n0_429_13410 1.074286e+00
R34357 n0_429_13410 n0_1366_13410 5.354286e+00
R34358 n0_1366_13410 n0_1554_13410 1.074286e+00
R34359 n0_1554_13410 n0_2491_13410 5.354286e+00
R34360 n0_2491_13410 n0_2679_13410 1.074286e+00
R34361 n0_2679_13410 n0_3616_13410 5.354286e+00
R34362 n0_3616_13410 n0_3804_13410 1.074286e+00
R34363 n0_3804_13410 n0_4741_13410 5.354286e+00
R34364 n0_4741_13410 n0_4929_13410 1.074286e+00
R34365 n0_4929_13410 n0_5866_13410 5.354286e+00
R34366 n0_5866_13410 n0_6054_13410 1.074286e+00
R34367 n0_6054_13410 n0_6991_13410 5.354286e+00
R34368 n0_6991_13410 n0_7179_13410 1.074286e+00
R34369 n0_7179_13410 n0_8116_13410 5.354286e+00
R34370 n0_8116_13410 n0_8208_13410 5.257143e-01
R34371 n0_8208_13410 n0_8304_13410 5.485714e-01
R34372 n0_8304_13410 n0_8396_13410 5.257143e-01
R34373 n0_8396_13410 n0_10366_13410 1.125714e+01
R34374 n0_10366_13410 n0_10458_13410 5.257143e-01
R34375 n0_10458_13410 n0_10554_13410 5.485714e-01
R34376 n0_10554_13410 n0_10646_13410 5.257143e-01
R34377 n0_10646_13410 n0_12616_13410 1.125714e+01
R34378 n0_12616_13410 n0_12708_13410 5.257143e-01
R34379 n0_12708_13410 n0_12804_13410 5.485714e-01
R34380 n0_12804_13410 n0_12896_13410 5.257143e-01
R34381 n0_12896_13410 n0_13741_13410 4.828571e+00
R34382 n0_13741_13410 n0_13929_13410 1.074286e+00
R34383 n0_13929_13410 n0_14866_13410 5.354286e+00
R34384 n0_14866_13410 n0_15054_13410 1.074286e+00
R34385 n0_15054_13410 n0_15991_13410 5.354286e+00
R34386 n0_15991_13410 n0_16179_13410 1.074286e+00
R34387 n0_16179_13410 n0_17116_13410 5.354286e+00
R34388 n0_17116_13410 n0_17304_13410 1.074286e+00
R34389 n0_17304_13410 n0_18241_13410 5.354286e+00
R34390 n0_18241_13410 n0_18429_13410 1.074286e+00
R34391 n0_18429_13410 n0_19366_13410 5.354286e+00
R34392 n0_19366_13410 n0_19554_13410 1.074286e+00
R34393 n0_19554_13410 n0_20491_13410 5.354286e+00
R34394 n0_20491_13410 n0_20679_13410 1.074286e+00
R34395 n0_241_13593 n0_429_13593 1.074286e+00
R34396 n0_429_13593 n0_1366_13593 5.354286e+00
R34397 n0_1366_13593 n0_1554_13593 1.074286e+00
R34398 n0_1554_13593 n0_2491_13593 5.354286e+00
R34399 n0_2491_13593 n0_2679_13593 1.074286e+00
R34400 n0_2679_13593 n0_3616_13593 5.354286e+00
R34401 n0_3616_13593 n0_3804_13593 1.074286e+00
R34402 n0_3804_13593 n0_4741_13593 5.354286e+00
R34403 n0_4741_13593 n0_4929_13593 1.074286e+00
R34404 n0_4929_13593 n0_5866_13593 5.354286e+00
R34405 n0_5866_13593 n0_6054_13593 1.074286e+00
R34406 n0_6054_13593 n0_6991_13593 5.354286e+00
R34407 n0_6991_13593 n0_7179_13593 1.074286e+00
R34408 n0_7179_13593 n0_8116_13593 5.354286e+00
R34409 n0_8116_13593 n0_8208_13593 5.257143e-01
R34410 n0_8208_13593 n0_8304_13593 5.485714e-01
R34411 n0_8304_13593 n0_8396_13593 5.257143e-01
R34412 n0_8396_13593 n0_10366_13593 1.125714e+01
R34413 n0_10366_13593 n0_10458_13593 5.257143e-01
R34414 n0_10458_13593 n0_10554_13593 5.485714e-01
R34415 n0_10554_13593 n0_10646_13593 5.257143e-01
R34416 n0_10646_13593 n0_12616_13593 1.125714e+01
R34417 n0_12616_13593 n0_12708_13593 5.257143e-01
R34418 n0_12708_13593 n0_12804_13593 5.485714e-01
R34419 n0_12804_13593 n0_12896_13593 5.257143e-01
R34420 n0_12896_13593 n0_13741_13593 4.828571e+00
R34421 n0_13741_13593 n0_13929_13593 1.074286e+00
R34422 n0_13929_13593 n0_14866_13593 5.354286e+00
R34423 n0_14866_13593 n0_15054_13593 1.074286e+00
R34424 n0_15054_13593 n0_15991_13593 5.354286e+00
R34425 n0_15991_13593 n0_16179_13593 1.074286e+00
R34426 n0_16179_13593 n0_17116_13593 5.354286e+00
R34427 n0_17116_13593 n0_17304_13593 1.074286e+00
R34428 n0_17304_13593 n0_18241_13593 5.354286e+00
R34429 n0_18241_13593 n0_18429_13593 1.074286e+00
R34430 n0_18429_13593 n0_19366_13593 5.354286e+00
R34431 n0_19366_13593 n0_19554_13593 1.074286e+00
R34432 n0_19554_13593 n0_20491_13593 5.354286e+00
R34433 n0_20491_13593 n0_20679_13593 1.074286e+00
R34434 n0_241_13626 n0_429_13626 1.074286e+00
R34435 n0_429_13626 n0_1366_13626 5.354286e+00
R34436 n0_1366_13626 n0_1554_13626 1.074286e+00
R34437 n0_1554_13626 n0_2491_13626 5.354286e+00
R34438 n0_2491_13626 n0_2679_13626 1.074286e+00
R34439 n0_2679_13626 n0_3616_13626 5.354286e+00
R34440 n0_3616_13626 n0_3804_13626 1.074286e+00
R34441 n0_3804_13626 n0_4741_13626 5.354286e+00
R34442 n0_4741_13626 n0_4929_13626 1.074286e+00
R34443 n0_4929_13626 n0_5866_13626 5.354286e+00
R34444 n0_5866_13626 n0_6054_13626 1.074286e+00
R34445 n0_6054_13626 n0_6991_13626 5.354286e+00
R34446 n0_6991_13626 n0_7179_13626 1.074286e+00
R34447 n0_7179_13626 n0_8116_13626 5.354286e+00
R34448 n0_8116_13626 n0_8208_13626 5.257143e-01
R34449 n0_8208_13626 n0_8304_13626 5.485714e-01
R34450 n0_8304_13626 n0_8396_13626 5.257143e-01
R34451 n0_8396_13626 n0_10366_13626 1.125714e+01
R34452 n0_10366_13626 n0_10458_13626 5.257143e-01
R34453 n0_10458_13626 n0_10554_13626 5.485714e-01
R34454 n0_10554_13626 n0_10646_13626 5.257143e-01
R34455 n0_10646_13626 n0_12616_13626 1.125714e+01
R34456 n0_12616_13626 n0_12708_13626 5.257143e-01
R34457 n0_12708_13626 n0_12804_13626 5.485714e-01
R34458 n0_12804_13626 n0_12896_13626 5.257143e-01
R34459 n0_12896_13626 n0_13741_13626 4.828571e+00
R34460 n0_13741_13626 n0_13929_13626 1.074286e+00
R34461 n0_13929_13626 n0_14866_13626 5.354286e+00
R34462 n0_14866_13626 n0_15054_13626 1.074286e+00
R34463 n0_15054_13626 n0_15991_13626 5.354286e+00
R34464 n0_15991_13626 n0_16179_13626 1.074286e+00
R34465 n0_16179_13626 n0_17116_13626 5.354286e+00
R34466 n0_17116_13626 n0_17304_13626 1.074286e+00
R34467 n0_17304_13626 n0_18241_13626 5.354286e+00
R34468 n0_18241_13626 n0_18429_13626 1.074286e+00
R34469 n0_18429_13626 n0_19366_13626 5.354286e+00
R34470 n0_19366_13626 n0_19554_13626 1.074286e+00
R34471 n0_19554_13626 n0_20491_13626 5.354286e+00
R34472 n0_20491_13626 n0_20679_13626 1.074286e+00
R34473 n0_241_13809 n0_429_13809 1.074286e+00
R34474 n0_429_13809 n0_1366_13809 5.354286e+00
R34475 n0_1366_13809 n0_1554_13809 1.074286e+00
R34476 n0_1554_13809 n0_2491_13809 5.354286e+00
R34477 n0_2491_13809 n0_2679_13809 1.074286e+00
R34478 n0_2679_13809 n0_3616_13809 5.354286e+00
R34479 n0_3616_13809 n0_3804_13809 1.074286e+00
R34480 n0_3804_13809 n0_4741_13809 5.354286e+00
R34481 n0_4741_13809 n0_4929_13809 1.074286e+00
R34482 n0_4929_13809 n0_5866_13809 5.354286e+00
R34483 n0_5866_13809 n0_6054_13809 1.074286e+00
R34484 n0_6054_13809 n0_6991_13809 5.354286e+00
R34485 n0_6991_13809 n0_7179_13809 1.074286e+00
R34486 n0_7179_13809 n0_8116_13809 5.354286e+00
R34487 n0_8116_13809 n0_8208_13809 5.257143e-01
R34488 n0_8208_13809 n0_8304_13809 5.485714e-01
R34489 n0_8304_13809 n0_8396_13809 5.257143e-01
R34490 n0_8396_13809 n0_10366_13809 1.125714e+01
R34491 n0_10366_13809 n0_10458_13809 5.257143e-01
R34492 n0_10458_13809 n0_10554_13809 5.485714e-01
R34493 n0_10554_13809 n0_10646_13809 5.257143e-01
R34494 n0_10646_13809 n0_12616_13809 1.125714e+01
R34495 n0_12616_13809 n0_12708_13809 5.257143e-01
R34496 n0_12708_13809 n0_12804_13809 5.485714e-01
R34497 n0_12804_13809 n0_12896_13809 5.257143e-01
R34498 n0_12896_13809 n0_13741_13809 4.828571e+00
R34499 n0_13741_13809 n0_13929_13809 1.074286e+00
R34500 n0_13929_13809 n0_14866_13809 5.354286e+00
R34501 n0_14866_13809 n0_15054_13809 1.074286e+00
R34502 n0_15054_13809 n0_15991_13809 5.354286e+00
R34503 n0_15991_13809 n0_16179_13809 1.074286e+00
R34504 n0_16179_13809 n0_17116_13809 5.354286e+00
R34505 n0_17116_13809 n0_17304_13809 1.074286e+00
R34506 n0_17304_13809 n0_18241_13809 5.354286e+00
R34507 n0_18241_13809 n0_18429_13809 1.074286e+00
R34508 n0_18429_13809 n0_19366_13809 5.354286e+00
R34509 n0_19366_13809 n0_19554_13809 1.074286e+00
R34510 n0_19554_13809 n0_20491_13809 5.354286e+00
R34511 n0_20491_13809 n0_20679_13809 1.074286e+00
R34512 n0_241_13842 n0_429_13842 1.074286e+00
R34513 n0_429_13842 n0_1366_13842 5.354286e+00
R34514 n0_1366_13842 n0_1554_13842 1.074286e+00
R34515 n0_1554_13842 n0_2491_13842 5.354286e+00
R34516 n0_2491_13842 n0_2679_13842 1.074286e+00
R34517 n0_2679_13842 n0_3616_13842 5.354286e+00
R34518 n0_3616_13842 n0_3804_13842 1.074286e+00
R34519 n0_3804_13842 n0_4741_13842 5.354286e+00
R34520 n0_4741_13842 n0_4929_13842 1.074286e+00
R34521 n0_4929_13842 n0_5866_13842 5.354286e+00
R34522 n0_5866_13842 n0_6054_13842 1.074286e+00
R34523 n0_6054_13842 n0_6991_13842 5.354286e+00
R34524 n0_6991_13842 n0_7179_13842 1.074286e+00
R34525 n0_7179_13842 n0_8116_13842 5.354286e+00
R34526 n0_8116_13842 n0_8208_13842 5.257143e-01
R34527 n0_8208_13842 n0_8304_13842 5.485714e-01
R34528 n0_8304_13842 n0_8396_13842 5.257143e-01
R34529 n0_8396_13842 n0_10366_13842 1.125714e+01
R34530 n0_10366_13842 n0_10458_13842 5.257143e-01
R34531 n0_10458_13842 n0_10554_13842 5.485714e-01
R34532 n0_10554_13842 n0_10646_13842 5.257143e-01
R34533 n0_10646_13842 n0_12616_13842 1.125714e+01
R34534 n0_12616_13842 n0_12708_13842 5.257143e-01
R34535 n0_12708_13842 n0_12804_13842 5.485714e-01
R34536 n0_12804_13842 n0_12896_13842 5.257143e-01
R34537 n0_12896_13842 n0_13741_13842 4.828571e+00
R34538 n0_13741_13842 n0_13929_13842 1.074286e+00
R34539 n0_13929_13842 n0_14866_13842 5.354286e+00
R34540 n0_14866_13842 n0_15054_13842 1.074286e+00
R34541 n0_15054_13842 n0_15991_13842 5.354286e+00
R34542 n0_15991_13842 n0_16179_13842 1.074286e+00
R34543 n0_16179_13842 n0_17116_13842 5.354286e+00
R34544 n0_17116_13842 n0_17304_13842 1.074286e+00
R34545 n0_17304_13842 n0_18241_13842 5.354286e+00
R34546 n0_18241_13842 n0_18429_13842 1.074286e+00
R34547 n0_18429_13842 n0_19366_13842 5.354286e+00
R34548 n0_19366_13842 n0_19554_13842 1.074286e+00
R34549 n0_19554_13842 n0_20491_13842 5.354286e+00
R34550 n0_20491_13842 n0_20679_13842 1.074286e+00
R34551 n0_241_14025 n0_1366_14025 6.428571e+00
R34552 n0_1366_14025 n0_2491_14025 6.428571e+00
R34553 n0_2491_14025 n0_3616_14025 6.428571e+00
R34554 n0_3616_14025 n0_4741_14025 6.428571e+00
R34555 n0_4741_14025 n0_5866_14025 6.428571e+00
R34556 n0_5866_14025 n0_8116_14025 1.285714e+01
R34557 n0_8116_14025 n0_8208_14025 5.257143e-01
R34558 n0_8208_14025 n0_8255_14025 2.685714e-01
R34559 n0_8255_14025 n0_8304_14025 2.800000e-01
R34560 n0_8304_14025 n0_8396_14025 5.257143e-01
R34561 n0_8396_14025 n0_10366_14025 1.125714e+01
R34562 n0_10366_14025 n0_10458_14025 5.257143e-01
R34563 n0_10458_14025 n0_10505_14025 2.685714e-01
R34564 n0_10505_14025 n0_10554_14025 2.800000e-01
R34565 n0_10554_14025 n0_10646_14025 5.257143e-01
R34566 n0_10646_14025 n0_12616_14025 1.125714e+01
R34567 n0_12616_14025 n0_12708_14025 5.257143e-01
R34568 n0_12708_14025 n0_12755_14025 2.685714e-01
R34569 n0_12755_14025 n0_12804_14025 2.800000e-01
R34570 n0_12804_14025 n0_12896_14025 5.257143e-01
R34571 n0_12896_14025 n0_14866_14025 1.125714e+01
R34572 n0_14866_14025 n0_15991_14025 6.428571e+00
R34573 n0_15991_14025 n0_17116_14025 6.428571e+00
R34574 n0_17116_14025 n0_18241_14025 6.428571e+00
R34575 n0_18241_14025 n0_19366_14025 6.428571e+00
R34576 n0_19366_14025 n0_20491_14025 6.428571e+00
R34577 n0_241_14058 n0_1366_14058 6.428571e+00
R34578 n0_1366_14058 n0_2491_14058 6.428571e+00
R34579 n0_2491_14058 n0_3616_14058 6.428571e+00
R34580 n0_3616_14058 n0_4741_14058 6.428571e+00
R34581 n0_4741_14058 n0_5866_14058 6.428571e+00
R34582 n0_5866_14058 n0_8116_14058 1.285714e+01
R34583 n0_8116_14058 n0_8208_14058 5.257143e-01
R34584 n0_8208_14058 n0_8304_14058 5.485714e-01
R34585 n0_8304_14058 n0_8396_14058 5.257143e-01
R34586 n0_8396_14058 n0_10366_14058 1.125714e+01
R34587 n0_10366_14058 n0_10458_14058 5.257143e-01
R34588 n0_10458_14058 n0_10554_14058 5.485714e-01
R34589 n0_10554_14058 n0_10646_14058 5.257143e-01
R34590 n0_10646_14058 n0_12616_14058 1.125714e+01
R34591 n0_12616_14058 n0_12708_14058 5.257143e-01
R34592 n0_12708_14058 n0_12804_14058 5.485714e-01
R34593 n0_12804_14058 n0_12896_14058 5.257143e-01
R34594 n0_12896_14058 n0_14866_14058 1.125714e+01
R34595 n0_14866_14058 n0_15991_14058 6.428571e+00
R34596 n0_15991_14058 n0_17116_14058 6.428571e+00
R34597 n0_17116_14058 n0_18241_14058 6.428571e+00
R34598 n0_18241_14058 n0_19366_14058 6.428571e+00
R34599 n0_19366_14058 n0_20491_14058 6.428571e+00
R34600 n0_241_14241 n0_429_14241 1.074286e+00
R34601 n0_429_14241 n0_1366_14241 5.354286e+00
R34602 n0_1366_14241 n0_1554_14241 1.074286e+00
R34603 n0_1554_14241 n0_2491_14241 5.354286e+00
R34604 n0_2491_14241 n0_2679_14241 1.074286e+00
R34605 n0_2679_14241 n0_3616_14241 5.354286e+00
R34606 n0_3616_14241 n0_3804_14241 1.074286e+00
R34607 n0_3804_14241 n0_4741_14241 5.354286e+00
R34608 n0_4741_14241 n0_4929_14241 1.074286e+00
R34609 n0_4929_14241 n0_5866_14241 5.354286e+00
R34610 n0_5866_14241 n0_6054_14241 1.074286e+00
R34611 n0_6054_14241 n0_8116_14241 1.178286e+01
R34612 n0_8116_14241 n0_8208_14241 5.257143e-01
R34613 n0_8208_14241 n0_8304_14241 5.485714e-01
R34614 n0_8304_14241 n0_8396_14241 5.257143e-01
R34615 n0_8396_14241 n0_10366_14241 1.125714e+01
R34616 n0_10366_14241 n0_10458_14241 5.257143e-01
R34617 n0_10458_14241 n0_10554_14241 5.485714e-01
R34618 n0_10554_14241 n0_10646_14241 5.257143e-01
R34619 n0_10646_14241 n0_12616_14241 1.125714e+01
R34620 n0_12616_14241 n0_12708_14241 5.257143e-01
R34621 n0_12708_14241 n0_12804_14241 5.485714e-01
R34622 n0_12804_14241 n0_12896_14241 5.257143e-01
R34623 n0_12896_14241 n0_14866_14241 1.125714e+01
R34624 n0_14866_14241 n0_15054_14241 1.074286e+00
R34625 n0_15054_14241 n0_15991_14241 5.354286e+00
R34626 n0_15991_14241 n0_16179_14241 1.074286e+00
R34627 n0_16179_14241 n0_17116_14241 5.354286e+00
R34628 n0_17116_14241 n0_17304_14241 1.074286e+00
R34629 n0_17304_14241 n0_18241_14241 5.354286e+00
R34630 n0_18241_14241 n0_18429_14241 1.074286e+00
R34631 n0_18429_14241 n0_19366_14241 5.354286e+00
R34632 n0_19366_14241 n0_19554_14241 1.074286e+00
R34633 n0_19554_14241 n0_20491_14241 5.354286e+00
R34634 n0_20491_14241 n0_20679_14241 1.074286e+00
R34635 n0_241_14274 n0_429_14274 1.074286e+00
R34636 n0_429_14274 n0_1366_14274 5.354286e+00
R34637 n0_1366_14274 n0_1554_14274 1.074286e+00
R34638 n0_1554_14274 n0_2491_14274 5.354286e+00
R34639 n0_2491_14274 n0_2679_14274 1.074286e+00
R34640 n0_2679_14274 n0_3616_14274 5.354286e+00
R34641 n0_3616_14274 n0_3804_14274 1.074286e+00
R34642 n0_3804_14274 n0_4741_14274 5.354286e+00
R34643 n0_4741_14274 n0_4929_14274 1.074286e+00
R34644 n0_4929_14274 n0_5866_14274 5.354286e+00
R34645 n0_5866_14274 n0_6054_14274 1.074286e+00
R34646 n0_6054_14274 n0_8116_14274 1.178286e+01
R34647 n0_8116_14274 n0_8208_14274 5.257143e-01
R34648 n0_8208_14274 n0_8304_14274 5.485714e-01
R34649 n0_8304_14274 n0_8396_14274 5.257143e-01
R34650 n0_8396_14274 n0_10366_14274 1.125714e+01
R34651 n0_10366_14274 n0_10458_14274 5.257143e-01
R34652 n0_10458_14274 n0_10554_14274 5.485714e-01
R34653 n0_10554_14274 n0_10646_14274 5.257143e-01
R34654 n0_10646_14274 n0_12616_14274 1.125714e+01
R34655 n0_12616_14274 n0_12708_14274 5.257143e-01
R34656 n0_12708_14274 n0_12804_14274 5.485714e-01
R34657 n0_12804_14274 n0_12896_14274 5.257143e-01
R34658 n0_12896_14274 n0_14866_14274 1.125714e+01
R34659 n0_14866_14274 n0_15054_14274 1.074286e+00
R34660 n0_15054_14274 n0_15991_14274 5.354286e+00
R34661 n0_15991_14274 n0_16179_14274 1.074286e+00
R34662 n0_16179_14274 n0_17116_14274 5.354286e+00
R34663 n0_17116_14274 n0_17304_14274 1.074286e+00
R34664 n0_17304_14274 n0_18241_14274 5.354286e+00
R34665 n0_18241_14274 n0_18429_14274 1.074286e+00
R34666 n0_18429_14274 n0_19366_14274 5.354286e+00
R34667 n0_19366_14274 n0_19554_14274 1.074286e+00
R34668 n0_19554_14274 n0_20491_14274 5.354286e+00
R34669 n0_20491_14274 n0_20679_14274 1.074286e+00
R34670 n0_241_14457 n0_429_14457 1.074286e+00
R34671 n0_429_14457 n0_1366_14457 5.354286e+00
R34672 n0_1366_14457 n0_1554_14457 1.074286e+00
R34673 n0_1554_14457 n0_2491_14457 5.354286e+00
R34674 n0_2491_14457 n0_2679_14457 1.074286e+00
R34675 n0_2679_14457 n0_3616_14457 5.354286e+00
R34676 n0_3616_14457 n0_3804_14457 1.074286e+00
R34677 n0_3804_14457 n0_4741_14457 5.354286e+00
R34678 n0_4741_14457 n0_4929_14457 1.074286e+00
R34679 n0_4929_14457 n0_5866_14457 5.354286e+00
R34680 n0_5866_14457 n0_6054_14457 1.074286e+00
R34681 n0_6054_14457 n0_8116_14457 1.178286e+01
R34682 n0_8116_14457 n0_8208_14457 5.257143e-01
R34683 n0_8208_14457 n0_8304_14457 5.485714e-01
R34684 n0_8304_14457 n0_8396_14457 5.257143e-01
R34685 n0_8396_14457 n0_10366_14457 1.125714e+01
R34686 n0_10366_14457 n0_10458_14457 5.257143e-01
R34687 n0_10458_14457 n0_10554_14457 5.485714e-01
R34688 n0_10554_14457 n0_10646_14457 5.257143e-01
R34689 n0_10646_14457 n0_12616_14457 1.125714e+01
R34690 n0_12616_14457 n0_12708_14457 5.257143e-01
R34691 n0_12708_14457 n0_12804_14457 5.485714e-01
R34692 n0_12804_14457 n0_12896_14457 5.257143e-01
R34693 n0_12896_14457 n0_14866_14457 1.125714e+01
R34694 n0_14866_14457 n0_15054_14457 1.074286e+00
R34695 n0_15054_14457 n0_15991_14457 5.354286e+00
R34696 n0_15991_14457 n0_16179_14457 1.074286e+00
R34697 n0_16179_14457 n0_17116_14457 5.354286e+00
R34698 n0_17116_14457 n0_17304_14457 1.074286e+00
R34699 n0_17304_14457 n0_18241_14457 5.354286e+00
R34700 n0_18241_14457 n0_18429_14457 1.074286e+00
R34701 n0_18429_14457 n0_19366_14457 5.354286e+00
R34702 n0_19366_14457 n0_19554_14457 1.074286e+00
R34703 n0_19554_14457 n0_20491_14457 5.354286e+00
R34704 n0_20491_14457 n0_20679_14457 1.074286e+00
R34705 n0_241_14490 n0_429_14490 1.074286e+00
R34706 n0_429_14490 n0_1366_14490 5.354286e+00
R34707 n0_1366_14490 n0_1554_14490 1.074286e+00
R34708 n0_1554_14490 n0_2491_14490 5.354286e+00
R34709 n0_2491_14490 n0_2679_14490 1.074286e+00
R34710 n0_2679_14490 n0_3616_14490 5.354286e+00
R34711 n0_3616_14490 n0_3804_14490 1.074286e+00
R34712 n0_3804_14490 n0_4741_14490 5.354286e+00
R34713 n0_4741_14490 n0_4929_14490 1.074286e+00
R34714 n0_4929_14490 n0_5866_14490 5.354286e+00
R34715 n0_5866_14490 n0_6054_14490 1.074286e+00
R34716 n0_6054_14490 n0_8116_14490 1.178286e+01
R34717 n0_8116_14490 n0_8208_14490 5.257143e-01
R34718 n0_8208_14490 n0_8304_14490 5.485714e-01
R34719 n0_8304_14490 n0_8396_14490 5.257143e-01
R34720 n0_8396_14490 n0_10366_14490 1.125714e+01
R34721 n0_10366_14490 n0_10458_14490 5.257143e-01
R34722 n0_10458_14490 n0_10554_14490 5.485714e-01
R34723 n0_10554_14490 n0_10646_14490 5.257143e-01
R34724 n0_10646_14490 n0_12616_14490 1.125714e+01
R34725 n0_12616_14490 n0_12708_14490 5.257143e-01
R34726 n0_12708_14490 n0_12804_14490 5.485714e-01
R34727 n0_12804_14490 n0_12896_14490 5.257143e-01
R34728 n0_12896_14490 n0_14866_14490 1.125714e+01
R34729 n0_14866_14490 n0_15054_14490 1.074286e+00
R34730 n0_15054_14490 n0_15991_14490 5.354286e+00
R34731 n0_15991_14490 n0_16179_14490 1.074286e+00
R34732 n0_16179_14490 n0_17116_14490 5.354286e+00
R34733 n0_17116_14490 n0_17304_14490 1.074286e+00
R34734 n0_17304_14490 n0_18241_14490 5.354286e+00
R34735 n0_18241_14490 n0_18429_14490 1.074286e+00
R34736 n0_18429_14490 n0_19366_14490 5.354286e+00
R34737 n0_19366_14490 n0_19554_14490 1.074286e+00
R34738 n0_19554_14490 n0_20491_14490 5.354286e+00
R34739 n0_20491_14490 n0_20679_14490 1.074286e+00
R34740 n0_241_14673 n0_429_14673 1.074286e+00
R34741 n0_429_14673 n0_1366_14673 5.354286e+00
R34742 n0_1366_14673 n0_1554_14673 1.074286e+00
R34743 n0_1554_14673 n0_2491_14673 5.354286e+00
R34744 n0_2491_14673 n0_2679_14673 1.074286e+00
R34745 n0_2679_14673 n0_3616_14673 5.354286e+00
R34746 n0_3616_14673 n0_3804_14673 1.074286e+00
R34747 n0_3804_14673 n0_4741_14673 5.354286e+00
R34748 n0_4741_14673 n0_4929_14673 1.074286e+00
R34749 n0_4929_14673 n0_5866_14673 5.354286e+00
R34750 n0_5866_14673 n0_6054_14673 1.074286e+00
R34751 n0_6054_14673 n0_8116_14673 1.178286e+01
R34752 n0_8116_14673 n0_8208_14673 5.257143e-01
R34753 n0_8208_14673 n0_8304_14673 5.485714e-01
R34754 n0_8304_14673 n0_8396_14673 5.257143e-01
R34755 n0_8396_14673 n0_10366_14673 1.125714e+01
R34756 n0_10366_14673 n0_10458_14673 5.257143e-01
R34757 n0_10458_14673 n0_10554_14673 5.485714e-01
R34758 n0_10554_14673 n0_10646_14673 5.257143e-01
R34759 n0_10646_14673 n0_12616_14673 1.125714e+01
R34760 n0_12616_14673 n0_12708_14673 5.257143e-01
R34761 n0_12708_14673 n0_12804_14673 5.485714e-01
R34762 n0_12804_14673 n0_12896_14673 5.257143e-01
R34763 n0_12896_14673 n0_14866_14673 1.125714e+01
R34764 n0_14866_14673 n0_15054_14673 1.074286e+00
R34765 n0_15054_14673 n0_15991_14673 5.354286e+00
R34766 n0_15991_14673 n0_16179_14673 1.074286e+00
R34767 n0_16179_14673 n0_17116_14673 5.354286e+00
R34768 n0_17116_14673 n0_17304_14673 1.074286e+00
R34769 n0_17304_14673 n0_18241_14673 5.354286e+00
R34770 n0_18241_14673 n0_18429_14673 1.074286e+00
R34771 n0_18429_14673 n0_19366_14673 5.354286e+00
R34772 n0_19366_14673 n0_19554_14673 1.074286e+00
R34773 n0_19554_14673 n0_20491_14673 5.354286e+00
R34774 n0_20491_14673 n0_20679_14673 1.074286e+00
R34775 n0_241_14706 n0_429_14706 1.074286e+00
R34776 n0_429_14706 n0_1366_14706 5.354286e+00
R34777 n0_1366_14706 n0_1554_14706 1.074286e+00
R34778 n0_1554_14706 n0_2491_14706 5.354286e+00
R34779 n0_2491_14706 n0_2679_14706 1.074286e+00
R34780 n0_2679_14706 n0_3616_14706 5.354286e+00
R34781 n0_3616_14706 n0_3804_14706 1.074286e+00
R34782 n0_3804_14706 n0_4741_14706 5.354286e+00
R34783 n0_4741_14706 n0_4929_14706 1.074286e+00
R34784 n0_4929_14706 n0_5866_14706 5.354286e+00
R34785 n0_5866_14706 n0_6054_14706 1.074286e+00
R34786 n0_6054_14706 n0_8116_14706 1.178286e+01
R34787 n0_8116_14706 n0_8208_14706 5.257143e-01
R34788 n0_8208_14706 n0_8304_14706 5.485714e-01
R34789 n0_8304_14706 n0_8396_14706 5.257143e-01
R34790 n0_8396_14706 n0_10366_14706 1.125714e+01
R34791 n0_10366_14706 n0_10458_14706 5.257143e-01
R34792 n0_10458_14706 n0_10554_14706 5.485714e-01
R34793 n0_10554_14706 n0_10646_14706 5.257143e-01
R34794 n0_10646_14706 n0_12616_14706 1.125714e+01
R34795 n0_12616_14706 n0_12708_14706 5.257143e-01
R34796 n0_12708_14706 n0_12804_14706 5.485714e-01
R34797 n0_12804_14706 n0_12896_14706 5.257143e-01
R34798 n0_12896_14706 n0_14866_14706 1.125714e+01
R34799 n0_14866_14706 n0_15054_14706 1.074286e+00
R34800 n0_15054_14706 n0_15991_14706 5.354286e+00
R34801 n0_15991_14706 n0_16179_14706 1.074286e+00
R34802 n0_16179_14706 n0_17116_14706 5.354286e+00
R34803 n0_17116_14706 n0_17304_14706 1.074286e+00
R34804 n0_17304_14706 n0_18241_14706 5.354286e+00
R34805 n0_18241_14706 n0_18429_14706 1.074286e+00
R34806 n0_18429_14706 n0_19366_14706 5.354286e+00
R34807 n0_19366_14706 n0_19554_14706 1.074286e+00
R34808 n0_19554_14706 n0_20491_14706 5.354286e+00
R34809 n0_20491_14706 n0_20679_14706 1.074286e+00
R34810 n0_241_14889 n0_429_14889 1.074286e+00
R34811 n0_429_14889 n0_1366_14889 5.354286e+00
R34812 n0_1366_14889 n0_1554_14889 1.074286e+00
R34813 n0_1554_14889 n0_2491_14889 5.354286e+00
R34814 n0_2491_14889 n0_2679_14889 1.074286e+00
R34815 n0_2679_14889 n0_3616_14889 5.354286e+00
R34816 n0_3616_14889 n0_3804_14889 1.074286e+00
R34817 n0_3804_14889 n0_4741_14889 5.354286e+00
R34818 n0_4741_14889 n0_4929_14889 1.074286e+00
R34819 n0_4929_14889 n0_5866_14889 5.354286e+00
R34820 n0_5866_14889 n0_6054_14889 1.074286e+00
R34821 n0_6054_14889 n0_8116_14889 1.178286e+01
R34822 n0_8116_14889 n0_8208_14889 5.257143e-01
R34823 n0_8208_14889 n0_8304_14889 5.485714e-01
R34824 n0_8304_14889 n0_8396_14889 5.257143e-01
R34825 n0_8396_14889 n0_10366_14889 1.125714e+01
R34826 n0_10366_14889 n0_10458_14889 5.257143e-01
R34827 n0_10458_14889 n0_10554_14889 5.485714e-01
R34828 n0_10554_14889 n0_10646_14889 5.257143e-01
R34829 n0_10646_14889 n0_12616_14889 1.125714e+01
R34830 n0_12616_14889 n0_12708_14889 5.257143e-01
R34831 n0_12708_14889 n0_12804_14889 5.485714e-01
R34832 n0_12804_14889 n0_12896_14889 5.257143e-01
R34833 n0_12896_14889 n0_14866_14889 1.125714e+01
R34834 n0_14866_14889 n0_15054_14889 1.074286e+00
R34835 n0_15054_14889 n0_15991_14889 5.354286e+00
R34836 n0_15991_14889 n0_16179_14889 1.074286e+00
R34837 n0_16179_14889 n0_17116_14889 5.354286e+00
R34838 n0_17116_14889 n0_17304_14889 1.074286e+00
R34839 n0_17304_14889 n0_18241_14889 5.354286e+00
R34840 n0_18241_14889 n0_18429_14889 1.074286e+00
R34841 n0_18429_14889 n0_19366_14889 5.354286e+00
R34842 n0_19366_14889 n0_19554_14889 1.074286e+00
R34843 n0_19554_14889 n0_20491_14889 5.354286e+00
R34844 n0_20491_14889 n0_20679_14889 1.074286e+00
R34845 n0_241_14922 n0_429_14922 1.074286e+00
R34846 n0_429_14922 n0_1366_14922 5.354286e+00
R34847 n0_1366_14922 n0_1554_14922 1.074286e+00
R34848 n0_1554_14922 n0_2491_14922 5.354286e+00
R34849 n0_2491_14922 n0_2679_14922 1.074286e+00
R34850 n0_2679_14922 n0_3616_14922 5.354286e+00
R34851 n0_3616_14922 n0_3804_14922 1.074286e+00
R34852 n0_3804_14922 n0_4741_14922 5.354286e+00
R34853 n0_4741_14922 n0_4929_14922 1.074286e+00
R34854 n0_4929_14922 n0_5866_14922 5.354286e+00
R34855 n0_5866_14922 n0_6054_14922 1.074286e+00
R34856 n0_6054_14922 n0_8116_14922 1.178286e+01
R34857 n0_8116_14922 n0_8208_14922 5.257143e-01
R34858 n0_8208_14922 n0_8304_14922 5.485714e-01
R34859 n0_8304_14922 n0_8396_14922 5.257143e-01
R34860 n0_8396_14922 n0_10366_14922 1.125714e+01
R34861 n0_10366_14922 n0_10458_14922 5.257143e-01
R34862 n0_10458_14922 n0_10554_14922 5.485714e-01
R34863 n0_10554_14922 n0_10646_14922 5.257143e-01
R34864 n0_10646_14922 n0_12616_14922 1.125714e+01
R34865 n0_12616_14922 n0_12708_14922 5.257143e-01
R34866 n0_12708_14922 n0_12804_14922 5.485714e-01
R34867 n0_12804_14922 n0_12896_14922 5.257143e-01
R34868 n0_12896_14922 n0_14866_14922 1.125714e+01
R34869 n0_14866_14922 n0_15054_14922 1.074286e+00
R34870 n0_15054_14922 n0_15991_14922 5.354286e+00
R34871 n0_15991_14922 n0_16179_14922 1.074286e+00
R34872 n0_16179_14922 n0_17116_14922 5.354286e+00
R34873 n0_17116_14922 n0_17304_14922 1.074286e+00
R34874 n0_17304_14922 n0_18241_14922 5.354286e+00
R34875 n0_18241_14922 n0_18429_14922 1.074286e+00
R34876 n0_18429_14922 n0_19366_14922 5.354286e+00
R34877 n0_19366_14922 n0_19554_14922 1.074286e+00
R34878 n0_19554_14922 n0_20491_14922 5.354286e+00
R34879 n0_20491_14922 n0_20679_14922 1.074286e+00
R34880 n0_380_15105 n0_429_15105 2.800000e-01
R34881 n0_429_15105 n0_1505_15105 6.148571e+00
R34882 n0_1505_15105 n0_1554_15105 2.800000e-01
R34883 n0_1554_15105 n0_2630_15105 6.148571e+00
R34884 n0_2630_15105 n0_2679_15105 2.800000e-01
R34885 n0_2679_15105 n0_3755_15105 6.148571e+00
R34886 n0_3755_15105 n0_3804_15105 2.800000e-01
R34887 n0_3804_15105 n0_4880_15105 6.148571e+00
R34888 n0_4880_15105 n0_4929_15105 2.800000e-01
R34889 n0_4929_15105 n0_5958_15105 5.880000e+00
R34890 n0_5958_15105 n0_6005_15105 2.685714e-01
R34891 n0_6005_15105 n0_6054_15105 2.800000e-01
R34892 n0_6054_15105 n0_8208_15105 1.230857e+01
R34893 n0_8208_15105 n0_8255_15105 2.685714e-01
R34894 n0_8255_15105 n0_8304_15105 2.800000e-01
R34895 n0_8304_15105 n0_10458_15105 1.230857e+01
R34896 n0_10458_15105 n0_10505_15105 2.685714e-01
R34897 n0_10505_15105 n0_10554_15105 2.800000e-01
R34898 n0_10554_15105 n0_12708_15105 1.230857e+01
R34899 n0_12708_15105 n0_12755_15105 2.685714e-01
R34900 n0_12755_15105 n0_12804_15105 2.800000e-01
R34901 n0_12804_15105 n0_14958_15105 1.230857e+01
R34902 n0_14958_15105 n0_15005_15105 2.685714e-01
R34903 n0_15005_15105 n0_15054_15105 2.800000e-01
R34904 n0_15054_15105 n0_16130_15105 6.148571e+00
R34905 n0_16130_15105 n0_16179_15105 2.800000e-01
R34906 n0_16179_15105 n0_17255_15105 6.148571e+00
R34907 n0_17255_15105 n0_17304_15105 2.800000e-01
R34908 n0_17304_15105 n0_18380_15105 6.148571e+00
R34909 n0_18380_15105 n0_18429_15105 2.800000e-01
R34910 n0_18429_15105 n0_19505_15105 6.148571e+00
R34911 n0_19505_15105 n0_19554_15105 2.800000e-01
R34912 n0_19554_15105 n0_20630_15105 6.148571e+00
R34913 n0_20630_15105 n0_20679_15105 2.800000e-01
R34914 n0_241_15138 n0_380_15138 7.942857e-01
R34915 n0_380_15138 n0_429_15138 2.800000e-01
R34916 n0_429_15138 n0_1366_15138 5.354286e+00
R34917 n0_1366_15138 n0_1505_15138 7.942857e-01
R34918 n0_1505_15138 n0_1554_15138 2.800000e-01
R34919 n0_1554_15138 n0_2491_15138 5.354286e+00
R34920 n0_2491_15138 n0_2630_15138 7.942857e-01
R34921 n0_2630_15138 n0_2679_15138 2.800000e-01
R34922 n0_2679_15138 n0_3616_15138 5.354286e+00
R34923 n0_3616_15138 n0_3755_15138 7.942857e-01
R34924 n0_3755_15138 n0_3804_15138 2.800000e-01
R34925 n0_3804_15138 n0_4741_15138 5.354286e+00
R34926 n0_4741_15138 n0_4880_15138 7.942857e-01
R34927 n0_4880_15138 n0_4929_15138 2.800000e-01
R34928 n0_4929_15138 n0_5866_15138 5.354286e+00
R34929 n0_5866_15138 n0_5958_15138 5.257143e-01
R34930 n0_5958_15138 n0_6005_15138 2.685714e-01
R34931 n0_6005_15138 n0_6054_15138 2.800000e-01
R34932 n0_6054_15138 n0_6146_15138 5.257143e-01
R34933 n0_6146_15138 n0_8116_15138 1.125714e+01
R34934 n0_8116_15138 n0_8208_15138 5.257143e-01
R34935 n0_8208_15138 n0_8255_15138 2.685714e-01
R34936 n0_8255_15138 n0_8304_15138 2.800000e-01
R34937 n0_8304_15138 n0_8396_15138 5.257143e-01
R34938 n0_8396_15138 n0_10366_15138 1.125714e+01
R34939 n0_10366_15138 n0_10458_15138 5.257143e-01
R34940 n0_10458_15138 n0_10505_15138 2.685714e-01
R34941 n0_10505_15138 n0_10554_15138 2.800000e-01
R34942 n0_10554_15138 n0_10646_15138 5.257143e-01
R34943 n0_10646_15138 n0_12616_15138 1.125714e+01
R34944 n0_12616_15138 n0_12708_15138 5.257143e-01
R34945 n0_12708_15138 n0_12755_15138 2.685714e-01
R34946 n0_12755_15138 n0_12804_15138 2.800000e-01
R34947 n0_12804_15138 n0_12896_15138 5.257143e-01
R34948 n0_12896_15138 n0_14866_15138 1.125714e+01
R34949 n0_14866_15138 n0_14958_15138 5.257143e-01
R34950 n0_14958_15138 n0_15005_15138 2.685714e-01
R34951 n0_15005_15138 n0_15054_15138 2.800000e-01
R34952 n0_15054_15138 n0_15146_15138 5.257143e-01
R34953 n0_15146_15138 n0_15991_15138 4.828571e+00
R34954 n0_15991_15138 n0_16130_15138 7.942857e-01
R34955 n0_16130_15138 n0_16179_15138 2.800000e-01
R34956 n0_16179_15138 n0_17116_15138 5.354286e+00
R34957 n0_17116_15138 n0_17255_15138 7.942857e-01
R34958 n0_17255_15138 n0_17304_15138 2.800000e-01
R34959 n0_17304_15138 n0_18241_15138 5.354286e+00
R34960 n0_18241_15138 n0_18380_15138 7.942857e-01
R34961 n0_18380_15138 n0_18429_15138 2.800000e-01
R34962 n0_18429_15138 n0_19366_15138 5.354286e+00
R34963 n0_19366_15138 n0_19505_15138 7.942857e-01
R34964 n0_19505_15138 n0_19554_15138 2.800000e-01
R34965 n0_19554_15138 n0_20491_15138 5.354286e+00
R34966 n0_20491_15138 n0_20630_15138 7.942857e-01
R34967 n0_20630_15138 n0_20679_15138 2.800000e-01
R34968 n0_241_15321 n0_429_15321 1.074286e+00
R34969 n0_429_15321 n0_1366_15321 5.354286e+00
R34970 n0_1366_15321 n0_1554_15321 1.074286e+00
R34971 n0_1554_15321 n0_2491_15321 5.354286e+00
R34972 n0_2491_15321 n0_2679_15321 1.074286e+00
R34973 n0_2679_15321 n0_3616_15321 5.354286e+00
R34974 n0_3616_15321 n0_3804_15321 1.074286e+00
R34975 n0_3804_15321 n0_4741_15321 5.354286e+00
R34976 n0_4741_15321 n0_4929_15321 1.074286e+00
R34977 n0_4929_15321 n0_5866_15321 5.354286e+00
R34978 n0_5866_15321 n0_5958_15321 5.257143e-01
R34979 n0_5958_15321 n0_6054_15321 5.485714e-01
R34980 n0_6054_15321 n0_6146_15321 5.257143e-01
R34981 n0_6146_15321 n0_8116_15321 1.125714e+01
R34982 n0_8116_15321 n0_8208_15321 5.257143e-01
R34983 n0_8208_15321 n0_8304_15321 5.485714e-01
R34984 n0_8304_15321 n0_8396_15321 5.257143e-01
R34985 n0_8396_15321 n0_10366_15321 1.125714e+01
R34986 n0_10366_15321 n0_10458_15321 5.257143e-01
R34987 n0_10458_15321 n0_10554_15321 5.485714e-01
R34988 n0_10554_15321 n0_10646_15321 5.257143e-01
R34989 n0_10646_15321 n0_12616_15321 1.125714e+01
R34990 n0_12616_15321 n0_12708_15321 5.257143e-01
R34991 n0_12708_15321 n0_12804_15321 5.485714e-01
R34992 n0_12804_15321 n0_12896_15321 5.257143e-01
R34993 n0_12896_15321 n0_14866_15321 1.125714e+01
R34994 n0_14866_15321 n0_14958_15321 5.257143e-01
R34995 n0_14958_15321 n0_15054_15321 5.485714e-01
R34996 n0_15054_15321 n0_15146_15321 5.257143e-01
R34997 n0_15146_15321 n0_15991_15321 4.828571e+00
R34998 n0_15991_15321 n0_16179_15321 1.074286e+00
R34999 n0_16179_15321 n0_17116_15321 5.354286e+00
R35000 n0_17116_15321 n0_17304_15321 1.074286e+00
R35001 n0_17304_15321 n0_18241_15321 5.354286e+00
R35002 n0_18241_15321 n0_18429_15321 1.074286e+00
R35003 n0_18429_15321 n0_19366_15321 5.354286e+00
R35004 n0_19366_15321 n0_19554_15321 1.074286e+00
R35005 n0_19554_15321 n0_20491_15321 5.354286e+00
R35006 n0_20491_15321 n0_20679_15321 1.074286e+00
R35007 n0_241_15354 n0_429_15354 1.074286e+00
R35008 n0_429_15354 n0_1366_15354 5.354286e+00
R35009 n0_1366_15354 n0_1554_15354 1.074286e+00
R35010 n0_1554_15354 n0_2491_15354 5.354286e+00
R35011 n0_2491_15354 n0_2679_15354 1.074286e+00
R35012 n0_2679_15354 n0_3616_15354 5.354286e+00
R35013 n0_3616_15354 n0_3804_15354 1.074286e+00
R35014 n0_3804_15354 n0_4741_15354 5.354286e+00
R35015 n0_4741_15354 n0_4929_15354 1.074286e+00
R35016 n0_4929_15354 n0_5866_15354 5.354286e+00
R35017 n0_5866_15354 n0_5958_15354 5.257143e-01
R35018 n0_5958_15354 n0_6054_15354 5.485714e-01
R35019 n0_6054_15354 n0_6146_15354 5.257143e-01
R35020 n0_6146_15354 n0_8116_15354 1.125714e+01
R35021 n0_8116_15354 n0_8208_15354 5.257143e-01
R35022 n0_8208_15354 n0_8304_15354 5.485714e-01
R35023 n0_8304_15354 n0_8396_15354 5.257143e-01
R35024 n0_8396_15354 n0_10366_15354 1.125714e+01
R35025 n0_10366_15354 n0_10458_15354 5.257143e-01
R35026 n0_10458_15354 n0_10554_15354 5.485714e-01
R35027 n0_10554_15354 n0_10646_15354 5.257143e-01
R35028 n0_10646_15354 n0_12616_15354 1.125714e+01
R35029 n0_12616_15354 n0_12708_15354 5.257143e-01
R35030 n0_12708_15354 n0_12804_15354 5.485714e-01
R35031 n0_12804_15354 n0_12896_15354 5.257143e-01
R35032 n0_12896_15354 n0_14866_15354 1.125714e+01
R35033 n0_14866_15354 n0_14958_15354 5.257143e-01
R35034 n0_14958_15354 n0_15054_15354 5.485714e-01
R35035 n0_15054_15354 n0_15146_15354 5.257143e-01
R35036 n0_15146_15354 n0_15991_15354 4.828571e+00
R35037 n0_15991_15354 n0_16179_15354 1.074286e+00
R35038 n0_16179_15354 n0_17116_15354 5.354286e+00
R35039 n0_17116_15354 n0_17304_15354 1.074286e+00
R35040 n0_17304_15354 n0_18241_15354 5.354286e+00
R35041 n0_18241_15354 n0_18429_15354 1.074286e+00
R35042 n0_18429_15354 n0_19366_15354 5.354286e+00
R35043 n0_19366_15354 n0_19554_15354 1.074286e+00
R35044 n0_19554_15354 n0_20491_15354 5.354286e+00
R35045 n0_20491_15354 n0_20679_15354 1.074286e+00
R35046 n0_241_15537 n0_429_15537 1.074286e+00
R35047 n0_429_15537 n0_1366_15537 5.354286e+00
R35048 n0_1366_15537 n0_1554_15537 1.074286e+00
R35049 n0_1554_15537 n0_2491_15537 5.354286e+00
R35050 n0_2491_15537 n0_2679_15537 1.074286e+00
R35051 n0_2679_15537 n0_3616_15537 5.354286e+00
R35052 n0_3616_15537 n0_3804_15537 1.074286e+00
R35053 n0_3804_15537 n0_4741_15537 5.354286e+00
R35054 n0_4741_15537 n0_4929_15537 1.074286e+00
R35055 n0_4929_15537 n0_5866_15537 5.354286e+00
R35056 n0_5866_15537 n0_5958_15537 5.257143e-01
R35057 n0_5958_15537 n0_6054_15537 5.485714e-01
R35058 n0_6054_15537 n0_6146_15537 5.257143e-01
R35059 n0_6146_15537 n0_8116_15537 1.125714e+01
R35060 n0_8116_15537 n0_8208_15537 5.257143e-01
R35061 n0_8208_15537 n0_8304_15537 5.485714e-01
R35062 n0_8304_15537 n0_8396_15537 5.257143e-01
R35063 n0_8396_15537 n0_10366_15537 1.125714e+01
R35064 n0_10366_15537 n0_10458_15537 5.257143e-01
R35065 n0_10458_15537 n0_10554_15537 5.485714e-01
R35066 n0_10554_15537 n0_10646_15537 5.257143e-01
R35067 n0_10646_15537 n0_12616_15537 1.125714e+01
R35068 n0_12616_15537 n0_12708_15537 5.257143e-01
R35069 n0_12708_15537 n0_12804_15537 5.485714e-01
R35070 n0_12804_15537 n0_12896_15537 5.257143e-01
R35071 n0_12896_15537 n0_14866_15537 1.125714e+01
R35072 n0_14866_15537 n0_14958_15537 5.257143e-01
R35073 n0_14958_15537 n0_15054_15537 5.485714e-01
R35074 n0_15054_15537 n0_15146_15537 5.257143e-01
R35075 n0_15146_15537 n0_15991_15537 4.828571e+00
R35076 n0_15991_15537 n0_16179_15537 1.074286e+00
R35077 n0_16179_15537 n0_17116_15537 5.354286e+00
R35078 n0_17116_15537 n0_17304_15537 1.074286e+00
R35079 n0_17304_15537 n0_18241_15537 5.354286e+00
R35080 n0_18241_15537 n0_18429_15537 1.074286e+00
R35081 n0_18429_15537 n0_19366_15537 5.354286e+00
R35082 n0_19366_15537 n0_19554_15537 1.074286e+00
R35083 n0_19554_15537 n0_20491_15537 5.354286e+00
R35084 n0_20491_15537 n0_20679_15537 1.074286e+00
R35085 n0_241_15570 n0_429_15570 1.074286e+00
R35086 n0_429_15570 n0_1366_15570 5.354286e+00
R35087 n0_1366_15570 n0_1554_15570 1.074286e+00
R35088 n0_1554_15570 n0_2491_15570 5.354286e+00
R35089 n0_2491_15570 n0_2679_15570 1.074286e+00
R35090 n0_2679_15570 n0_3616_15570 5.354286e+00
R35091 n0_3616_15570 n0_3804_15570 1.074286e+00
R35092 n0_3804_15570 n0_4741_15570 5.354286e+00
R35093 n0_4741_15570 n0_4929_15570 1.074286e+00
R35094 n0_4929_15570 n0_5866_15570 5.354286e+00
R35095 n0_5866_15570 n0_5958_15570 5.257143e-01
R35096 n0_5958_15570 n0_6054_15570 5.485714e-01
R35097 n0_6054_15570 n0_6146_15570 5.257143e-01
R35098 n0_6146_15570 n0_8116_15570 1.125714e+01
R35099 n0_8116_15570 n0_8208_15570 5.257143e-01
R35100 n0_8208_15570 n0_8304_15570 5.485714e-01
R35101 n0_8304_15570 n0_8396_15570 5.257143e-01
R35102 n0_8396_15570 n0_10366_15570 1.125714e+01
R35103 n0_10366_15570 n0_10458_15570 5.257143e-01
R35104 n0_10458_15570 n0_10554_15570 5.485714e-01
R35105 n0_10554_15570 n0_10646_15570 5.257143e-01
R35106 n0_10646_15570 n0_12616_15570 1.125714e+01
R35107 n0_12616_15570 n0_12708_15570 5.257143e-01
R35108 n0_12708_15570 n0_12804_15570 5.485714e-01
R35109 n0_12804_15570 n0_12896_15570 5.257143e-01
R35110 n0_12896_15570 n0_14866_15570 1.125714e+01
R35111 n0_14866_15570 n0_14958_15570 5.257143e-01
R35112 n0_14958_15570 n0_15054_15570 5.485714e-01
R35113 n0_15054_15570 n0_15146_15570 5.257143e-01
R35114 n0_15146_15570 n0_15991_15570 4.828571e+00
R35115 n0_15991_15570 n0_16179_15570 1.074286e+00
R35116 n0_16179_15570 n0_17116_15570 5.354286e+00
R35117 n0_17116_15570 n0_17304_15570 1.074286e+00
R35118 n0_17304_15570 n0_18241_15570 5.354286e+00
R35119 n0_18241_15570 n0_18429_15570 1.074286e+00
R35120 n0_18429_15570 n0_19366_15570 5.354286e+00
R35121 n0_19366_15570 n0_19554_15570 1.074286e+00
R35122 n0_19554_15570 n0_20491_15570 5.354286e+00
R35123 n0_20491_15570 n0_20679_15570 1.074286e+00
R35124 n0_241_15753 n0_429_15753 1.074286e+00
R35125 n0_429_15753 n0_1366_15753 5.354286e+00
R35126 n0_1366_15753 n0_1554_15753 1.074286e+00
R35127 n0_1554_15753 n0_2491_15753 5.354286e+00
R35128 n0_2491_15753 n0_2679_15753 1.074286e+00
R35129 n0_2679_15753 n0_3616_15753 5.354286e+00
R35130 n0_3616_15753 n0_3804_15753 1.074286e+00
R35131 n0_3804_15753 n0_4741_15753 5.354286e+00
R35132 n0_4741_15753 n0_4929_15753 1.074286e+00
R35133 n0_4929_15753 n0_5866_15753 5.354286e+00
R35134 n0_5866_15753 n0_5958_15753 5.257143e-01
R35135 n0_5958_15753 n0_6054_15753 5.485714e-01
R35136 n0_6054_15753 n0_6146_15753 5.257143e-01
R35137 n0_6146_15753 n0_8116_15753 1.125714e+01
R35138 n0_8116_15753 n0_8208_15753 5.257143e-01
R35139 n0_8208_15753 n0_8304_15753 5.485714e-01
R35140 n0_8304_15753 n0_8396_15753 5.257143e-01
R35141 n0_8396_15753 n0_10366_15753 1.125714e+01
R35142 n0_10366_15753 n0_10458_15753 5.257143e-01
R35143 n0_10458_15753 n0_10554_15753 5.485714e-01
R35144 n0_10554_15753 n0_10646_15753 5.257143e-01
R35145 n0_10646_15753 n0_12616_15753 1.125714e+01
R35146 n0_12616_15753 n0_12708_15753 5.257143e-01
R35147 n0_12708_15753 n0_12804_15753 5.485714e-01
R35148 n0_12804_15753 n0_12896_15753 5.257143e-01
R35149 n0_12896_15753 n0_14866_15753 1.125714e+01
R35150 n0_14866_15753 n0_14958_15753 5.257143e-01
R35151 n0_14958_15753 n0_15054_15753 5.485714e-01
R35152 n0_15054_15753 n0_15146_15753 5.257143e-01
R35153 n0_15146_15753 n0_15991_15753 4.828571e+00
R35154 n0_15991_15753 n0_16179_15753 1.074286e+00
R35155 n0_16179_15753 n0_17116_15753 5.354286e+00
R35156 n0_17116_15753 n0_17304_15753 1.074286e+00
R35157 n0_17304_15753 n0_18241_15753 5.354286e+00
R35158 n0_18241_15753 n0_18429_15753 1.074286e+00
R35159 n0_18429_15753 n0_19366_15753 5.354286e+00
R35160 n0_19366_15753 n0_19554_15753 1.074286e+00
R35161 n0_19554_15753 n0_20491_15753 5.354286e+00
R35162 n0_20491_15753 n0_20679_15753 1.074286e+00
R35163 n0_241_15786 n0_429_15786 1.074286e+00
R35164 n0_429_15786 n0_1366_15786 5.354286e+00
R35165 n0_1366_15786 n0_1554_15786 1.074286e+00
R35166 n0_1554_15786 n0_2491_15786 5.354286e+00
R35167 n0_2491_15786 n0_2679_15786 1.074286e+00
R35168 n0_2679_15786 n0_3616_15786 5.354286e+00
R35169 n0_3616_15786 n0_3804_15786 1.074286e+00
R35170 n0_3804_15786 n0_4741_15786 5.354286e+00
R35171 n0_4741_15786 n0_4929_15786 1.074286e+00
R35172 n0_4929_15786 n0_5866_15786 5.354286e+00
R35173 n0_5866_15786 n0_5958_15786 5.257143e-01
R35174 n0_5958_15786 n0_6054_15786 5.485714e-01
R35175 n0_6054_15786 n0_6146_15786 5.257143e-01
R35176 n0_6146_15786 n0_8116_15786 1.125714e+01
R35177 n0_8116_15786 n0_8208_15786 5.257143e-01
R35178 n0_8208_15786 n0_8304_15786 5.485714e-01
R35179 n0_8304_15786 n0_8396_15786 5.257143e-01
R35180 n0_8396_15786 n0_10366_15786 1.125714e+01
R35181 n0_10366_15786 n0_10458_15786 5.257143e-01
R35182 n0_10458_15786 n0_10554_15786 5.485714e-01
R35183 n0_10554_15786 n0_10646_15786 5.257143e-01
R35184 n0_10646_15786 n0_12616_15786 1.125714e+01
R35185 n0_12616_15786 n0_12708_15786 5.257143e-01
R35186 n0_12708_15786 n0_12804_15786 5.485714e-01
R35187 n0_12804_15786 n0_12896_15786 5.257143e-01
R35188 n0_12896_15786 n0_14866_15786 1.125714e+01
R35189 n0_14866_15786 n0_14958_15786 5.257143e-01
R35190 n0_14958_15786 n0_15054_15786 5.485714e-01
R35191 n0_15054_15786 n0_15146_15786 5.257143e-01
R35192 n0_15146_15786 n0_15991_15786 4.828571e+00
R35193 n0_15991_15786 n0_16179_15786 1.074286e+00
R35194 n0_16179_15786 n0_17116_15786 5.354286e+00
R35195 n0_17116_15786 n0_17304_15786 1.074286e+00
R35196 n0_17304_15786 n0_18241_15786 5.354286e+00
R35197 n0_18241_15786 n0_18429_15786 1.074286e+00
R35198 n0_18429_15786 n0_19366_15786 5.354286e+00
R35199 n0_19366_15786 n0_19554_15786 1.074286e+00
R35200 n0_19554_15786 n0_20491_15786 5.354286e+00
R35201 n0_20491_15786 n0_20679_15786 1.074286e+00
R35202 n0_241_15969 n0_429_15969 1.074286e+00
R35203 n0_429_15969 n0_1366_15969 5.354286e+00
R35204 n0_1366_15969 n0_1554_15969 1.074286e+00
R35205 n0_1554_15969 n0_2491_15969 5.354286e+00
R35206 n0_2491_15969 n0_2679_15969 1.074286e+00
R35207 n0_2679_15969 n0_3616_15969 5.354286e+00
R35208 n0_3616_15969 n0_3804_15969 1.074286e+00
R35209 n0_3804_15969 n0_4741_15969 5.354286e+00
R35210 n0_4741_15969 n0_4929_15969 1.074286e+00
R35211 n0_4929_15969 n0_5866_15969 5.354286e+00
R35212 n0_5866_15969 n0_5958_15969 5.257143e-01
R35213 n0_5958_15969 n0_6054_15969 5.485714e-01
R35214 n0_6054_15969 n0_6146_15969 5.257143e-01
R35215 n0_6146_15969 n0_8116_15969 1.125714e+01
R35216 n0_8116_15969 n0_8208_15969 5.257143e-01
R35217 n0_8208_15969 n0_8304_15969 5.485714e-01
R35218 n0_8304_15969 n0_8396_15969 5.257143e-01
R35219 n0_8396_15969 n0_10366_15969 1.125714e+01
R35220 n0_10366_15969 n0_10458_15969 5.257143e-01
R35221 n0_10458_15969 n0_10554_15969 5.485714e-01
R35222 n0_10554_15969 n0_10646_15969 5.257143e-01
R35223 n0_10646_15969 n0_12616_15969 1.125714e+01
R35224 n0_12616_15969 n0_12708_15969 5.257143e-01
R35225 n0_12708_15969 n0_12804_15969 5.485714e-01
R35226 n0_12804_15969 n0_12896_15969 5.257143e-01
R35227 n0_12896_15969 n0_14866_15969 1.125714e+01
R35228 n0_14866_15969 n0_14958_15969 5.257143e-01
R35229 n0_14958_15969 n0_15054_15969 5.485714e-01
R35230 n0_15054_15969 n0_15146_15969 5.257143e-01
R35231 n0_15146_15969 n0_15991_15969 4.828571e+00
R35232 n0_15991_15969 n0_16179_15969 1.074286e+00
R35233 n0_16179_15969 n0_17116_15969 5.354286e+00
R35234 n0_17116_15969 n0_17304_15969 1.074286e+00
R35235 n0_17304_15969 n0_18241_15969 5.354286e+00
R35236 n0_18241_15969 n0_18429_15969 1.074286e+00
R35237 n0_18429_15969 n0_19366_15969 5.354286e+00
R35238 n0_19366_15969 n0_19554_15969 1.074286e+00
R35239 n0_19554_15969 n0_20491_15969 5.354286e+00
R35240 n0_20491_15969 n0_20679_15969 1.074286e+00
R35241 n0_241_16002 n0_429_16002 1.074286e+00
R35242 n0_429_16002 n0_1366_16002 5.354286e+00
R35243 n0_1366_16002 n0_1554_16002 1.074286e+00
R35244 n0_1554_16002 n0_2491_16002 5.354286e+00
R35245 n0_2491_16002 n0_2679_16002 1.074286e+00
R35246 n0_2679_16002 n0_3616_16002 5.354286e+00
R35247 n0_3616_16002 n0_3804_16002 1.074286e+00
R35248 n0_3804_16002 n0_4741_16002 5.354286e+00
R35249 n0_4741_16002 n0_4929_16002 1.074286e+00
R35250 n0_4929_16002 n0_5866_16002 5.354286e+00
R35251 n0_5866_16002 n0_5958_16002 5.257143e-01
R35252 n0_5958_16002 n0_6054_16002 5.485714e-01
R35253 n0_6054_16002 n0_6146_16002 5.257143e-01
R35254 n0_6146_16002 n0_8116_16002 1.125714e+01
R35255 n0_8116_16002 n0_8208_16002 5.257143e-01
R35256 n0_8208_16002 n0_8304_16002 5.485714e-01
R35257 n0_8304_16002 n0_8396_16002 5.257143e-01
R35258 n0_8396_16002 n0_10366_16002 1.125714e+01
R35259 n0_10366_16002 n0_10458_16002 5.257143e-01
R35260 n0_10458_16002 n0_10554_16002 5.485714e-01
R35261 n0_10554_16002 n0_10646_16002 5.257143e-01
R35262 n0_10646_16002 n0_12616_16002 1.125714e+01
R35263 n0_12616_16002 n0_12708_16002 5.257143e-01
R35264 n0_12708_16002 n0_12804_16002 5.485714e-01
R35265 n0_12804_16002 n0_12896_16002 5.257143e-01
R35266 n0_12896_16002 n0_14866_16002 1.125714e+01
R35267 n0_14866_16002 n0_14958_16002 5.257143e-01
R35268 n0_14958_16002 n0_15054_16002 5.485714e-01
R35269 n0_15054_16002 n0_15146_16002 5.257143e-01
R35270 n0_15146_16002 n0_15991_16002 4.828571e+00
R35271 n0_15991_16002 n0_16179_16002 1.074286e+00
R35272 n0_16179_16002 n0_17116_16002 5.354286e+00
R35273 n0_17116_16002 n0_17304_16002 1.074286e+00
R35274 n0_17304_16002 n0_18241_16002 5.354286e+00
R35275 n0_18241_16002 n0_18429_16002 1.074286e+00
R35276 n0_18429_16002 n0_19366_16002 5.354286e+00
R35277 n0_19366_16002 n0_19554_16002 1.074286e+00
R35278 n0_19554_16002 n0_20491_16002 5.354286e+00
R35279 n0_20491_16002 n0_20679_16002 1.074286e+00
R35280 n0_241_16185 n0_1366_16185 6.428571e+00
R35281 n0_1366_16185 n0_2491_16185 6.428571e+00
R35282 n0_2491_16185 n0_3616_16185 6.428571e+00
R35283 n0_3616_16185 n0_4741_16185 6.428571e+00
R35284 n0_4741_16185 n0_5866_16185 6.428571e+00
R35285 n0_5866_16185 n0_5958_16185 5.257143e-01
R35286 n0_5958_16185 n0_6005_16185 2.685714e-01
R35287 n0_6005_16185 n0_6054_16185 2.800000e-01
R35288 n0_6054_16185 n0_6146_16185 5.257143e-01
R35289 n0_6146_16185 n0_8116_16185 1.125714e+01
R35290 n0_8116_16185 n0_8208_16185 5.257143e-01
R35291 n0_8208_16185 n0_8255_16185 2.685714e-01
R35292 n0_8255_16185 n0_8304_16185 2.800000e-01
R35293 n0_8304_16185 n0_8396_16185 5.257143e-01
R35294 n0_8396_16185 n0_10366_16185 1.125714e+01
R35295 n0_10366_16185 n0_10458_16185 5.257143e-01
R35296 n0_10458_16185 n0_10505_16185 2.685714e-01
R35297 n0_10505_16185 n0_10554_16185 2.800000e-01
R35298 n0_10554_16185 n0_10646_16185 5.257143e-01
R35299 n0_10646_16185 n0_12616_16185 1.125714e+01
R35300 n0_12616_16185 n0_12708_16185 5.257143e-01
R35301 n0_12708_16185 n0_12755_16185 2.685714e-01
R35302 n0_12755_16185 n0_12804_16185 2.800000e-01
R35303 n0_12804_16185 n0_12896_16185 5.257143e-01
R35304 n0_12896_16185 n0_14866_16185 1.125714e+01
R35305 n0_14866_16185 n0_14958_16185 5.257143e-01
R35306 n0_14958_16185 n0_15005_16185 2.685714e-01
R35307 n0_15005_16185 n0_15054_16185 2.800000e-01
R35308 n0_15054_16185 n0_15146_16185 5.257143e-01
R35309 n0_15146_16185 n0_15991_16185 4.828571e+00
R35310 n0_15991_16185 n0_17116_16185 6.428571e+00
R35311 n0_17116_16185 n0_18241_16185 6.428571e+00
R35312 n0_18241_16185 n0_19366_16185 6.428571e+00
R35313 n0_19366_16185 n0_20491_16185 6.428571e+00
R35314 n0_241_16218 n0_1366_16218 6.428571e+00
R35315 n0_1366_16218 n0_2491_16218 6.428571e+00
R35316 n0_2491_16218 n0_3616_16218 6.428571e+00
R35317 n0_3616_16218 n0_5958_16218 1.338286e+01
R35318 n0_5958_16218 n0_6005_16218 2.685714e-01
R35319 n0_6005_16218 n0_6054_16218 2.800000e-01
R35320 n0_6054_16218 n0_8208_16218 1.230857e+01
R35321 n0_8208_16218 n0_8255_16218 2.685714e-01
R35322 n0_8255_16218 n0_8304_16218 2.800000e-01
R35323 n0_8304_16218 n0_10458_16218 1.230857e+01
R35324 n0_10458_16218 n0_10505_16218 2.685714e-01
R35325 n0_10505_16218 n0_10554_16218 2.800000e-01
R35326 n0_10554_16218 n0_12708_16218 1.230857e+01
R35327 n0_12708_16218 n0_12755_16218 2.685714e-01
R35328 n0_12755_16218 n0_12804_16218 2.800000e-01
R35329 n0_12804_16218 n0_14958_16218 1.230857e+01
R35330 n0_14958_16218 n0_15005_16218 2.685714e-01
R35331 n0_15005_16218 n0_15054_16218 2.800000e-01
R35332 n0_15054_16218 n0_17116_16218 1.178286e+01
R35333 n0_17116_16218 n0_18241_16218 6.428571e+00
R35334 n0_18241_16218 n0_19366_16218 6.428571e+00
R35335 n0_19366_16218 n0_20491_16218 6.428571e+00
R35336 n0_241_16401 n0_429_16401 1.074286e+00
R35337 n0_429_16401 n0_1366_16401 5.354286e+00
R35338 n0_1366_16401 n0_1554_16401 1.074286e+00
R35339 n0_1554_16401 n0_2491_16401 5.354286e+00
R35340 n0_2491_16401 n0_2679_16401 1.074286e+00
R35341 n0_2679_16401 n0_3616_16401 5.354286e+00
R35342 n0_3616_16401 n0_3804_16401 1.074286e+00
R35343 n0_3804_16401 n0_5866_16401 1.178286e+01
R35344 n0_5866_16401 n0_5958_16401 5.257143e-01
R35345 n0_5958_16401 n0_6054_16401 5.485714e-01
R35346 n0_6054_16401 n0_6146_16401 5.257143e-01
R35347 n0_6146_16401 n0_8116_16401 1.125714e+01
R35348 n0_8116_16401 n0_8208_16401 5.257143e-01
R35349 n0_8208_16401 n0_8304_16401 5.485714e-01
R35350 n0_8304_16401 n0_8396_16401 5.257143e-01
R35351 n0_8396_16401 n0_10366_16401 1.125714e+01
R35352 n0_10366_16401 n0_10458_16401 5.257143e-01
R35353 n0_10458_16401 n0_10554_16401 5.485714e-01
R35354 n0_10554_16401 n0_10646_16401 5.257143e-01
R35355 n0_10646_16401 n0_12616_16401 1.125714e+01
R35356 n0_12616_16401 n0_12708_16401 5.257143e-01
R35357 n0_12708_16401 n0_12804_16401 5.485714e-01
R35358 n0_12804_16401 n0_12896_16401 5.257143e-01
R35359 n0_12896_16401 n0_14866_16401 1.125714e+01
R35360 n0_14866_16401 n0_14958_16401 5.257143e-01
R35361 n0_14958_16401 n0_15054_16401 5.485714e-01
R35362 n0_15054_16401 n0_15146_16401 5.257143e-01
R35363 n0_15146_16401 n0_17116_16401 1.125714e+01
R35364 n0_17116_16401 n0_17304_16401 1.074286e+00
R35365 n0_17304_16401 n0_18241_16401 5.354286e+00
R35366 n0_18241_16401 n0_18429_16401 1.074286e+00
R35367 n0_18429_16401 n0_19366_16401 5.354286e+00
R35368 n0_19366_16401 n0_19554_16401 1.074286e+00
R35369 n0_19554_16401 n0_20491_16401 5.354286e+00
R35370 n0_20491_16401 n0_20679_16401 1.074286e+00
R35371 n0_241_16434 n0_429_16434 1.074286e+00
R35372 n0_429_16434 n0_1366_16434 5.354286e+00
R35373 n0_1366_16434 n0_1554_16434 1.074286e+00
R35374 n0_1554_16434 n0_2491_16434 5.354286e+00
R35375 n0_2491_16434 n0_2679_16434 1.074286e+00
R35376 n0_2679_16434 n0_3616_16434 5.354286e+00
R35377 n0_3616_16434 n0_3804_16434 1.074286e+00
R35378 n0_3804_16434 n0_5866_16434 1.178286e+01
R35379 n0_5866_16434 n0_5958_16434 5.257143e-01
R35380 n0_5958_16434 n0_6054_16434 5.485714e-01
R35381 n0_6054_16434 n0_6146_16434 5.257143e-01
R35382 n0_6146_16434 n0_8116_16434 1.125714e+01
R35383 n0_8116_16434 n0_8208_16434 5.257143e-01
R35384 n0_8208_16434 n0_8304_16434 5.485714e-01
R35385 n0_8304_16434 n0_8396_16434 5.257143e-01
R35386 n0_8396_16434 n0_10366_16434 1.125714e+01
R35387 n0_10366_16434 n0_10458_16434 5.257143e-01
R35388 n0_10458_16434 n0_10554_16434 5.485714e-01
R35389 n0_10554_16434 n0_10646_16434 5.257143e-01
R35390 n0_10646_16434 n0_12616_16434 1.125714e+01
R35391 n0_12616_16434 n0_12708_16434 5.257143e-01
R35392 n0_12708_16434 n0_12804_16434 5.485714e-01
R35393 n0_12804_16434 n0_12896_16434 5.257143e-01
R35394 n0_12896_16434 n0_14866_16434 1.125714e+01
R35395 n0_14866_16434 n0_14958_16434 5.257143e-01
R35396 n0_14958_16434 n0_15054_16434 5.485714e-01
R35397 n0_15054_16434 n0_15146_16434 5.257143e-01
R35398 n0_15146_16434 n0_17116_16434 1.125714e+01
R35399 n0_17116_16434 n0_17304_16434 1.074286e+00
R35400 n0_17304_16434 n0_18241_16434 5.354286e+00
R35401 n0_18241_16434 n0_18429_16434 1.074286e+00
R35402 n0_18429_16434 n0_19366_16434 5.354286e+00
R35403 n0_19366_16434 n0_19554_16434 1.074286e+00
R35404 n0_19554_16434 n0_20491_16434 5.354286e+00
R35405 n0_20491_16434 n0_20679_16434 1.074286e+00
R35406 n0_241_16617 n0_429_16617 1.074286e+00
R35407 n0_429_16617 n0_1366_16617 5.354286e+00
R35408 n0_1366_16617 n0_1554_16617 1.074286e+00
R35409 n0_1554_16617 n0_2491_16617 5.354286e+00
R35410 n0_2491_16617 n0_2679_16617 1.074286e+00
R35411 n0_2679_16617 n0_3616_16617 5.354286e+00
R35412 n0_3616_16617 n0_3804_16617 1.074286e+00
R35413 n0_3804_16617 n0_5866_16617 1.178286e+01
R35414 n0_5866_16617 n0_5958_16617 5.257143e-01
R35415 n0_5958_16617 n0_6054_16617 5.485714e-01
R35416 n0_6054_16617 n0_6146_16617 5.257143e-01
R35417 n0_6146_16617 n0_8116_16617 1.125714e+01
R35418 n0_8116_16617 n0_8208_16617 5.257143e-01
R35419 n0_8208_16617 n0_8304_16617 5.485714e-01
R35420 n0_8304_16617 n0_8396_16617 5.257143e-01
R35421 n0_8396_16617 n0_10366_16617 1.125714e+01
R35422 n0_10366_16617 n0_10458_16617 5.257143e-01
R35423 n0_10458_16617 n0_10554_16617 5.485714e-01
R35424 n0_10554_16617 n0_10646_16617 5.257143e-01
R35425 n0_10646_16617 n0_12616_16617 1.125714e+01
R35426 n0_12616_16617 n0_12708_16617 5.257143e-01
R35427 n0_12708_16617 n0_12804_16617 5.485714e-01
R35428 n0_12804_16617 n0_12896_16617 5.257143e-01
R35429 n0_12896_16617 n0_14866_16617 1.125714e+01
R35430 n0_14866_16617 n0_14958_16617 5.257143e-01
R35431 n0_14958_16617 n0_15054_16617 5.485714e-01
R35432 n0_15054_16617 n0_15146_16617 5.257143e-01
R35433 n0_15146_16617 n0_17116_16617 1.125714e+01
R35434 n0_17116_16617 n0_17304_16617 1.074286e+00
R35435 n0_17304_16617 n0_18241_16617 5.354286e+00
R35436 n0_18241_16617 n0_18429_16617 1.074286e+00
R35437 n0_18429_16617 n0_19366_16617 5.354286e+00
R35438 n0_19366_16617 n0_19554_16617 1.074286e+00
R35439 n0_19554_16617 n0_20491_16617 5.354286e+00
R35440 n0_20491_16617 n0_20679_16617 1.074286e+00
R35441 n0_241_16650 n0_429_16650 1.074286e+00
R35442 n0_429_16650 n0_1366_16650 5.354286e+00
R35443 n0_1366_16650 n0_1554_16650 1.074286e+00
R35444 n0_1554_16650 n0_2491_16650 5.354286e+00
R35445 n0_2491_16650 n0_2679_16650 1.074286e+00
R35446 n0_2679_16650 n0_3616_16650 5.354286e+00
R35447 n0_3616_16650 n0_3804_16650 1.074286e+00
R35448 n0_3804_16650 n0_5866_16650 1.178286e+01
R35449 n0_5866_16650 n0_5958_16650 5.257143e-01
R35450 n0_5958_16650 n0_6054_16650 5.485714e-01
R35451 n0_6054_16650 n0_6146_16650 5.257143e-01
R35452 n0_6146_16650 n0_8116_16650 1.125714e+01
R35453 n0_8116_16650 n0_8208_16650 5.257143e-01
R35454 n0_8208_16650 n0_8304_16650 5.485714e-01
R35455 n0_8304_16650 n0_8396_16650 5.257143e-01
R35456 n0_8396_16650 n0_10366_16650 1.125714e+01
R35457 n0_10366_16650 n0_10458_16650 5.257143e-01
R35458 n0_10458_16650 n0_10554_16650 5.485714e-01
R35459 n0_10554_16650 n0_10646_16650 5.257143e-01
R35460 n0_10646_16650 n0_12616_16650 1.125714e+01
R35461 n0_12616_16650 n0_12708_16650 5.257143e-01
R35462 n0_12708_16650 n0_12804_16650 5.485714e-01
R35463 n0_12804_16650 n0_12896_16650 5.257143e-01
R35464 n0_12896_16650 n0_14866_16650 1.125714e+01
R35465 n0_14866_16650 n0_14958_16650 5.257143e-01
R35466 n0_14958_16650 n0_15054_16650 5.485714e-01
R35467 n0_15054_16650 n0_15146_16650 5.257143e-01
R35468 n0_15146_16650 n0_17116_16650 1.125714e+01
R35469 n0_17116_16650 n0_17304_16650 1.074286e+00
R35470 n0_17304_16650 n0_18241_16650 5.354286e+00
R35471 n0_18241_16650 n0_18429_16650 1.074286e+00
R35472 n0_18429_16650 n0_19366_16650 5.354286e+00
R35473 n0_19366_16650 n0_19554_16650 1.074286e+00
R35474 n0_19554_16650 n0_20491_16650 5.354286e+00
R35475 n0_20491_16650 n0_20679_16650 1.074286e+00
R35476 n0_241_16833 n0_429_16833 1.074286e+00
R35477 n0_429_16833 n0_1366_16833 5.354286e+00
R35478 n0_1366_16833 n0_1554_16833 1.074286e+00
R35479 n0_1554_16833 n0_2491_16833 5.354286e+00
R35480 n0_2491_16833 n0_2679_16833 1.074286e+00
R35481 n0_2679_16833 n0_3616_16833 5.354286e+00
R35482 n0_3616_16833 n0_3804_16833 1.074286e+00
R35483 n0_3804_16833 n0_5866_16833 1.178286e+01
R35484 n0_5866_16833 n0_5958_16833 5.257143e-01
R35485 n0_5958_16833 n0_6054_16833 5.485714e-01
R35486 n0_6054_16833 n0_6146_16833 5.257143e-01
R35487 n0_6146_16833 n0_8116_16833 1.125714e+01
R35488 n0_8116_16833 n0_8208_16833 5.257143e-01
R35489 n0_8208_16833 n0_8304_16833 5.485714e-01
R35490 n0_8304_16833 n0_8396_16833 5.257143e-01
R35491 n0_8396_16833 n0_10366_16833 1.125714e+01
R35492 n0_10366_16833 n0_10458_16833 5.257143e-01
R35493 n0_10458_16833 n0_10554_16833 5.485714e-01
R35494 n0_10554_16833 n0_10646_16833 5.257143e-01
R35495 n0_10646_16833 n0_12616_16833 1.125714e+01
R35496 n0_12616_16833 n0_12708_16833 5.257143e-01
R35497 n0_12708_16833 n0_12804_16833 5.485714e-01
R35498 n0_12804_16833 n0_12896_16833 5.257143e-01
R35499 n0_12896_16833 n0_14866_16833 1.125714e+01
R35500 n0_14866_16833 n0_14958_16833 5.257143e-01
R35501 n0_14958_16833 n0_15054_16833 5.485714e-01
R35502 n0_15054_16833 n0_15146_16833 5.257143e-01
R35503 n0_15146_16833 n0_17116_16833 1.125714e+01
R35504 n0_17116_16833 n0_17304_16833 1.074286e+00
R35505 n0_17304_16833 n0_18241_16833 5.354286e+00
R35506 n0_18241_16833 n0_18429_16833 1.074286e+00
R35507 n0_18429_16833 n0_19366_16833 5.354286e+00
R35508 n0_19366_16833 n0_19554_16833 1.074286e+00
R35509 n0_19554_16833 n0_20491_16833 5.354286e+00
R35510 n0_20491_16833 n0_20679_16833 1.074286e+00
R35511 n0_241_16866 n0_429_16866 1.074286e+00
R35512 n0_429_16866 n0_1366_16866 5.354286e+00
R35513 n0_1366_16866 n0_1554_16866 1.074286e+00
R35514 n0_1554_16866 n0_2491_16866 5.354286e+00
R35515 n0_2491_16866 n0_2679_16866 1.074286e+00
R35516 n0_2679_16866 n0_3616_16866 5.354286e+00
R35517 n0_3616_16866 n0_3804_16866 1.074286e+00
R35518 n0_3804_16866 n0_5866_16866 1.178286e+01
R35519 n0_5866_16866 n0_5958_16866 5.257143e-01
R35520 n0_5958_16866 n0_6054_16866 5.485714e-01
R35521 n0_6054_16866 n0_6146_16866 5.257143e-01
R35522 n0_6146_16866 n0_8116_16866 1.125714e+01
R35523 n0_8116_16866 n0_8208_16866 5.257143e-01
R35524 n0_8208_16866 n0_8304_16866 5.485714e-01
R35525 n0_8304_16866 n0_8396_16866 5.257143e-01
R35526 n0_8396_16866 n0_10366_16866 1.125714e+01
R35527 n0_10366_16866 n0_10458_16866 5.257143e-01
R35528 n0_10458_16866 n0_10554_16866 5.485714e-01
R35529 n0_10554_16866 n0_10646_16866 5.257143e-01
R35530 n0_10646_16866 n0_12616_16866 1.125714e+01
R35531 n0_12616_16866 n0_12708_16866 5.257143e-01
R35532 n0_12708_16866 n0_12804_16866 5.485714e-01
R35533 n0_12804_16866 n0_12896_16866 5.257143e-01
R35534 n0_12896_16866 n0_14866_16866 1.125714e+01
R35535 n0_14866_16866 n0_14958_16866 5.257143e-01
R35536 n0_14958_16866 n0_15054_16866 5.485714e-01
R35537 n0_15054_16866 n0_15146_16866 5.257143e-01
R35538 n0_15146_16866 n0_17116_16866 1.125714e+01
R35539 n0_17116_16866 n0_17304_16866 1.074286e+00
R35540 n0_17304_16866 n0_18241_16866 5.354286e+00
R35541 n0_18241_16866 n0_18429_16866 1.074286e+00
R35542 n0_18429_16866 n0_19366_16866 5.354286e+00
R35543 n0_19366_16866 n0_19554_16866 1.074286e+00
R35544 n0_19554_16866 n0_20491_16866 5.354286e+00
R35545 n0_20491_16866 n0_20679_16866 1.074286e+00
R35546 n0_241_17049 n0_429_17049 1.074286e+00
R35547 n0_429_17049 n0_1366_17049 5.354286e+00
R35548 n0_1366_17049 n0_1554_17049 1.074286e+00
R35549 n0_1554_17049 n0_2491_17049 5.354286e+00
R35550 n0_2491_17049 n0_2679_17049 1.074286e+00
R35551 n0_2679_17049 n0_3616_17049 5.354286e+00
R35552 n0_3616_17049 n0_3804_17049 1.074286e+00
R35553 n0_3804_17049 n0_5866_17049 1.178286e+01
R35554 n0_5866_17049 n0_5958_17049 5.257143e-01
R35555 n0_5958_17049 n0_6054_17049 5.485714e-01
R35556 n0_6054_17049 n0_6146_17049 5.257143e-01
R35557 n0_6146_17049 n0_8116_17049 1.125714e+01
R35558 n0_8116_17049 n0_8208_17049 5.257143e-01
R35559 n0_8208_17049 n0_8304_17049 5.485714e-01
R35560 n0_8304_17049 n0_8396_17049 5.257143e-01
R35561 n0_8396_17049 n0_10366_17049 1.125714e+01
R35562 n0_10366_17049 n0_10458_17049 5.257143e-01
R35563 n0_10458_17049 n0_10554_17049 5.485714e-01
R35564 n0_10554_17049 n0_10646_17049 5.257143e-01
R35565 n0_10646_17049 n0_12616_17049 1.125714e+01
R35566 n0_12616_17049 n0_12708_17049 5.257143e-01
R35567 n0_12708_17049 n0_12804_17049 5.485714e-01
R35568 n0_12804_17049 n0_12896_17049 5.257143e-01
R35569 n0_12896_17049 n0_14866_17049 1.125714e+01
R35570 n0_14866_17049 n0_14958_17049 5.257143e-01
R35571 n0_14958_17049 n0_15054_17049 5.485714e-01
R35572 n0_15054_17049 n0_15146_17049 5.257143e-01
R35573 n0_15146_17049 n0_17116_17049 1.125714e+01
R35574 n0_17116_17049 n0_17304_17049 1.074286e+00
R35575 n0_17304_17049 n0_18241_17049 5.354286e+00
R35576 n0_18241_17049 n0_18429_17049 1.074286e+00
R35577 n0_18429_17049 n0_19366_17049 5.354286e+00
R35578 n0_19366_17049 n0_19554_17049 1.074286e+00
R35579 n0_19554_17049 n0_20491_17049 5.354286e+00
R35580 n0_20491_17049 n0_20679_17049 1.074286e+00
R35581 n0_241_17082 n0_429_17082 1.074286e+00
R35582 n0_429_17082 n0_1366_17082 5.354286e+00
R35583 n0_1366_17082 n0_1554_17082 1.074286e+00
R35584 n0_1554_17082 n0_2491_17082 5.354286e+00
R35585 n0_2491_17082 n0_2679_17082 1.074286e+00
R35586 n0_2679_17082 n0_3616_17082 5.354286e+00
R35587 n0_3616_17082 n0_3804_17082 1.074286e+00
R35588 n0_3804_17082 n0_5866_17082 1.178286e+01
R35589 n0_5866_17082 n0_5958_17082 5.257143e-01
R35590 n0_5958_17082 n0_6054_17082 5.485714e-01
R35591 n0_6054_17082 n0_6146_17082 5.257143e-01
R35592 n0_6146_17082 n0_8116_17082 1.125714e+01
R35593 n0_8116_17082 n0_8208_17082 5.257143e-01
R35594 n0_8208_17082 n0_8304_17082 5.485714e-01
R35595 n0_8304_17082 n0_8396_17082 5.257143e-01
R35596 n0_8396_17082 n0_10366_17082 1.125714e+01
R35597 n0_10366_17082 n0_10458_17082 5.257143e-01
R35598 n0_10458_17082 n0_10554_17082 5.485714e-01
R35599 n0_10554_17082 n0_10646_17082 5.257143e-01
R35600 n0_10646_17082 n0_12616_17082 1.125714e+01
R35601 n0_12616_17082 n0_12708_17082 5.257143e-01
R35602 n0_12708_17082 n0_12804_17082 5.485714e-01
R35603 n0_12804_17082 n0_12896_17082 5.257143e-01
R35604 n0_12896_17082 n0_14866_17082 1.125714e+01
R35605 n0_14866_17082 n0_14958_17082 5.257143e-01
R35606 n0_14958_17082 n0_15054_17082 5.485714e-01
R35607 n0_15054_17082 n0_15146_17082 5.257143e-01
R35608 n0_15146_17082 n0_17116_17082 1.125714e+01
R35609 n0_17116_17082 n0_17304_17082 1.074286e+00
R35610 n0_17304_17082 n0_18241_17082 5.354286e+00
R35611 n0_18241_17082 n0_18429_17082 1.074286e+00
R35612 n0_18429_17082 n0_19366_17082 5.354286e+00
R35613 n0_19366_17082 n0_19554_17082 1.074286e+00
R35614 n0_19554_17082 n0_20491_17082 5.354286e+00
R35615 n0_20491_17082 n0_20679_17082 1.074286e+00
R35616 n0_241_17265 n0_429_17265 1.074286e+00
R35617 n0_429_17265 n0_1366_17265 5.354286e+00
R35618 n0_1366_17265 n0_1554_17265 1.074286e+00
R35619 n0_1554_17265 n0_2491_17265 5.354286e+00
R35620 n0_2491_17265 n0_2679_17265 1.074286e+00
R35621 n0_2679_17265 n0_3616_17265 5.354286e+00
R35622 n0_3616_17265 n0_3708_17265 5.257143e-01
R35623 n0_3708_17265 n0_3804_17265 5.485714e-01
R35624 n0_3804_17265 n0_5866_17265 1.178286e+01
R35625 n0_5866_17265 n0_5958_17265 5.257143e-01
R35626 n0_5958_17265 n0_6054_17265 5.485714e-01
R35627 n0_6054_17265 n0_6146_17265 5.257143e-01
R35628 n0_6146_17265 n0_8116_17265 1.125714e+01
R35629 n0_8116_17265 n0_8208_17265 5.257143e-01
R35630 n0_8208_17265 n0_8304_17265 5.485714e-01
R35631 n0_8304_17265 n0_8396_17265 5.257143e-01
R35632 n0_8396_17265 n0_10366_17265 1.125714e+01
R35633 n0_10366_17265 n0_10458_17265 5.257143e-01
R35634 n0_10458_17265 n0_10554_17265 5.485714e-01
R35635 n0_10554_17265 n0_10646_17265 5.257143e-01
R35636 n0_10646_17265 n0_12616_17265 1.125714e+01
R35637 n0_12616_17265 n0_12708_17265 5.257143e-01
R35638 n0_12708_17265 n0_12804_17265 5.485714e-01
R35639 n0_12804_17265 n0_12896_17265 5.257143e-01
R35640 n0_12896_17265 n0_14866_17265 1.125714e+01
R35641 n0_14866_17265 n0_14958_17265 5.257143e-01
R35642 n0_14958_17265 n0_15054_17265 5.485714e-01
R35643 n0_15054_17265 n0_15146_17265 5.257143e-01
R35644 n0_15146_17265 n0_17116_17265 1.125714e+01
R35645 n0_17116_17265 n0_17208_17265 5.257143e-01
R35646 n0_17208_17265 n0_17304_17265 5.485714e-01
R35647 n0_17304_17265 n0_18241_17265 5.354286e+00
R35648 n0_18241_17265 n0_18429_17265 1.074286e+00
R35649 n0_18429_17265 n0_19366_17265 5.354286e+00
R35650 n0_19366_17265 n0_19554_17265 1.074286e+00
R35651 n0_19554_17265 n0_20491_17265 5.354286e+00
R35652 n0_20491_17265 n0_20679_17265 1.074286e+00
R35653 n0_241_17298 n0_380_17298 7.942857e-01
R35654 n0_380_17298 n0_429_17298 2.800000e-01
R35655 n0_429_17298 n0_1366_17298 5.354286e+00
R35656 n0_1366_17298 n0_1505_17298 7.942857e-01
R35657 n0_1505_17298 n0_1554_17298 2.800000e-01
R35658 n0_1554_17298 n0_2491_17298 5.354286e+00
R35659 n0_2491_17298 n0_2630_17298 7.942857e-01
R35660 n0_2630_17298 n0_2679_17298 2.800000e-01
R35661 n0_2679_17298 n0_3616_17298 5.354286e+00
R35662 n0_3616_17298 n0_3708_17298 5.257143e-01
R35663 n0_3708_17298 n0_3755_17298 2.685714e-01
R35664 n0_3755_17298 n0_3804_17298 2.800000e-01
R35665 n0_3804_17298 n0_5866_17298 1.178286e+01
R35666 n0_5866_17298 n0_5958_17298 5.257143e-01
R35667 n0_5958_17298 n0_6005_17298 2.685714e-01
R35668 n0_6005_17298 n0_6054_17298 2.800000e-01
R35669 n0_6054_17298 n0_6146_17298 5.257143e-01
R35670 n0_6146_17298 n0_8116_17298 1.125714e+01
R35671 n0_8116_17298 n0_8208_17298 5.257143e-01
R35672 n0_8208_17298 n0_8255_17298 2.685714e-01
R35673 n0_8255_17298 n0_8304_17298 2.800000e-01
R35674 n0_8304_17298 n0_8396_17298 5.257143e-01
R35675 n0_8396_17298 n0_10366_17298 1.125714e+01
R35676 n0_10366_17298 n0_10458_17298 5.257143e-01
R35677 n0_10458_17298 n0_10505_17298 2.685714e-01
R35678 n0_10505_17298 n0_10554_17298 2.800000e-01
R35679 n0_10554_17298 n0_10646_17298 5.257143e-01
R35680 n0_10646_17298 n0_12616_17298 1.125714e+01
R35681 n0_12616_17298 n0_12708_17298 5.257143e-01
R35682 n0_12708_17298 n0_12755_17298 2.685714e-01
R35683 n0_12755_17298 n0_12804_17298 2.800000e-01
R35684 n0_12804_17298 n0_12896_17298 5.257143e-01
R35685 n0_12896_17298 n0_14866_17298 1.125714e+01
R35686 n0_14866_17298 n0_14958_17298 5.257143e-01
R35687 n0_14958_17298 n0_15005_17298 2.685714e-01
R35688 n0_15005_17298 n0_15054_17298 2.800000e-01
R35689 n0_15054_17298 n0_15146_17298 5.257143e-01
R35690 n0_15146_17298 n0_17116_17298 1.125714e+01
R35691 n0_17116_17298 n0_17208_17298 5.257143e-01
R35692 n0_17208_17298 n0_17255_17298 2.685714e-01
R35693 n0_17255_17298 n0_17304_17298 2.800000e-01
R35694 n0_17304_17298 n0_18241_17298 5.354286e+00
R35695 n0_18241_17298 n0_18380_17298 7.942857e-01
R35696 n0_18380_17298 n0_18429_17298 2.800000e-01
R35697 n0_18429_17298 n0_19366_17298 5.354286e+00
R35698 n0_19366_17298 n0_19505_17298 7.942857e-01
R35699 n0_19505_17298 n0_19554_17298 2.800000e-01
R35700 n0_19554_17298 n0_20491_17298 5.354286e+00
R35701 n0_20491_17298 n0_20630_17298 7.942857e-01
R35702 n0_20630_17298 n0_20679_17298 2.800000e-01
R35703 n0_241_17481 n0_429_17481 1.074286e+00
R35704 n0_429_17481 n0_1366_17481 5.354286e+00
R35705 n0_1366_17481 n0_1554_17481 1.074286e+00
R35706 n0_1554_17481 n0_2491_17481 5.354286e+00
R35707 n0_2491_17481 n0_2679_17481 1.074286e+00
R35708 n0_2679_17481 n0_3616_17481 5.354286e+00
R35709 n0_3616_17481 n0_3708_17481 5.257143e-01
R35710 n0_3708_17481 n0_3804_17481 5.485714e-01
R35711 n0_3804_17481 n0_3896_17481 5.257143e-01
R35712 n0_3896_17481 n0_5866_17481 1.125714e+01
R35713 n0_5866_17481 n0_5958_17481 5.257143e-01
R35714 n0_5958_17481 n0_6054_17481 5.485714e-01
R35715 n0_6054_17481 n0_6146_17481 5.257143e-01
R35716 n0_6146_17481 n0_8116_17481 1.125714e+01
R35717 n0_8116_17481 n0_8208_17481 5.257143e-01
R35718 n0_8208_17481 n0_8304_17481 5.485714e-01
R35719 n0_8304_17481 n0_8396_17481 5.257143e-01
R35720 n0_8396_17481 n0_10366_17481 1.125714e+01
R35721 n0_10366_17481 n0_10458_17481 5.257143e-01
R35722 n0_10458_17481 n0_10554_17481 5.485714e-01
R35723 n0_10554_17481 n0_10646_17481 5.257143e-01
R35724 n0_10646_17481 n0_12616_17481 1.125714e+01
R35725 n0_12616_17481 n0_12708_17481 5.257143e-01
R35726 n0_12708_17481 n0_12804_17481 5.485714e-01
R35727 n0_12804_17481 n0_12896_17481 5.257143e-01
R35728 n0_12896_17481 n0_14866_17481 1.125714e+01
R35729 n0_14866_17481 n0_14958_17481 5.257143e-01
R35730 n0_14958_17481 n0_15054_17481 5.485714e-01
R35731 n0_15054_17481 n0_15146_17481 5.257143e-01
R35732 n0_15146_17481 n0_17116_17481 1.125714e+01
R35733 n0_17116_17481 n0_17208_17481 5.257143e-01
R35734 n0_17208_17481 n0_17304_17481 5.485714e-01
R35735 n0_17304_17481 n0_17396_17481 5.257143e-01
R35736 n0_17396_17481 n0_18241_17481 4.828571e+00
R35737 n0_18241_17481 n0_18429_17481 1.074286e+00
R35738 n0_18429_17481 n0_19366_17481 5.354286e+00
R35739 n0_19366_17481 n0_19554_17481 1.074286e+00
R35740 n0_19554_17481 n0_20491_17481 5.354286e+00
R35741 n0_20491_17481 n0_20679_17481 1.074286e+00
R35742 n0_241_17514 n0_429_17514 1.074286e+00
R35743 n0_429_17514 n0_1366_17514 5.354286e+00
R35744 n0_1366_17514 n0_1554_17514 1.074286e+00
R35745 n0_1554_17514 n0_2491_17514 5.354286e+00
R35746 n0_2491_17514 n0_2679_17514 1.074286e+00
R35747 n0_2679_17514 n0_3616_17514 5.354286e+00
R35748 n0_3616_17514 n0_3708_17514 5.257143e-01
R35749 n0_3708_17514 n0_3804_17514 5.485714e-01
R35750 n0_3804_17514 n0_3896_17514 5.257143e-01
R35751 n0_3896_17514 n0_5866_17514 1.125714e+01
R35752 n0_5866_17514 n0_5958_17514 5.257143e-01
R35753 n0_5958_17514 n0_6054_17514 5.485714e-01
R35754 n0_6054_17514 n0_6146_17514 5.257143e-01
R35755 n0_6146_17514 n0_8116_17514 1.125714e+01
R35756 n0_8116_17514 n0_8208_17514 5.257143e-01
R35757 n0_8208_17514 n0_8304_17514 5.485714e-01
R35758 n0_8304_17514 n0_8396_17514 5.257143e-01
R35759 n0_8396_17514 n0_10366_17514 1.125714e+01
R35760 n0_10366_17514 n0_10458_17514 5.257143e-01
R35761 n0_10458_17514 n0_10554_17514 5.485714e-01
R35762 n0_10554_17514 n0_10646_17514 5.257143e-01
R35763 n0_10646_17514 n0_12616_17514 1.125714e+01
R35764 n0_12616_17514 n0_12708_17514 5.257143e-01
R35765 n0_12708_17514 n0_12804_17514 5.485714e-01
R35766 n0_12804_17514 n0_12896_17514 5.257143e-01
R35767 n0_12896_17514 n0_14866_17514 1.125714e+01
R35768 n0_14866_17514 n0_14958_17514 5.257143e-01
R35769 n0_14958_17514 n0_15054_17514 5.485714e-01
R35770 n0_15054_17514 n0_15146_17514 5.257143e-01
R35771 n0_15146_17514 n0_17116_17514 1.125714e+01
R35772 n0_17116_17514 n0_17208_17514 5.257143e-01
R35773 n0_17208_17514 n0_17304_17514 5.485714e-01
R35774 n0_17304_17514 n0_17396_17514 5.257143e-01
R35775 n0_17396_17514 n0_18241_17514 4.828571e+00
R35776 n0_18241_17514 n0_18429_17514 1.074286e+00
R35777 n0_18429_17514 n0_19366_17514 5.354286e+00
R35778 n0_19366_17514 n0_19554_17514 1.074286e+00
R35779 n0_19554_17514 n0_20491_17514 5.354286e+00
R35780 n0_20491_17514 n0_20679_17514 1.074286e+00
R35781 n0_241_17697 n0_429_17697 1.074286e+00
R35782 n0_429_17697 n0_1366_17697 5.354286e+00
R35783 n0_1366_17697 n0_1554_17697 1.074286e+00
R35784 n0_1554_17697 n0_2491_17697 5.354286e+00
R35785 n0_2491_17697 n0_2679_17697 1.074286e+00
R35786 n0_2679_17697 n0_3616_17697 5.354286e+00
R35787 n0_3616_17697 n0_3708_17697 5.257143e-01
R35788 n0_3708_17697 n0_3804_17697 5.485714e-01
R35789 n0_3804_17697 n0_3896_17697 5.257143e-01
R35790 n0_3896_17697 n0_5866_17697 1.125714e+01
R35791 n0_5866_17697 n0_5958_17697 5.257143e-01
R35792 n0_5958_17697 n0_6054_17697 5.485714e-01
R35793 n0_6054_17697 n0_6146_17697 5.257143e-01
R35794 n0_6146_17697 n0_8116_17697 1.125714e+01
R35795 n0_8116_17697 n0_8208_17697 5.257143e-01
R35796 n0_8208_17697 n0_8304_17697 5.485714e-01
R35797 n0_8304_17697 n0_8396_17697 5.257143e-01
R35798 n0_8396_17697 n0_10366_17697 1.125714e+01
R35799 n0_10366_17697 n0_10458_17697 5.257143e-01
R35800 n0_10458_17697 n0_10554_17697 5.485714e-01
R35801 n0_10554_17697 n0_10646_17697 5.257143e-01
R35802 n0_10646_17697 n0_12616_17697 1.125714e+01
R35803 n0_12616_17697 n0_12708_17697 5.257143e-01
R35804 n0_12708_17697 n0_12804_17697 5.485714e-01
R35805 n0_12804_17697 n0_12896_17697 5.257143e-01
R35806 n0_12896_17697 n0_14866_17697 1.125714e+01
R35807 n0_14866_17697 n0_14958_17697 5.257143e-01
R35808 n0_14958_17697 n0_15054_17697 5.485714e-01
R35809 n0_15054_17697 n0_15146_17697 5.257143e-01
R35810 n0_15146_17697 n0_17116_17697 1.125714e+01
R35811 n0_17116_17697 n0_17208_17697 5.257143e-01
R35812 n0_17208_17697 n0_17304_17697 5.485714e-01
R35813 n0_17304_17697 n0_17396_17697 5.257143e-01
R35814 n0_17396_17697 n0_18241_17697 4.828571e+00
R35815 n0_18241_17697 n0_18429_17697 1.074286e+00
R35816 n0_18429_17697 n0_19366_17697 5.354286e+00
R35817 n0_19366_17697 n0_19554_17697 1.074286e+00
R35818 n0_19554_17697 n0_20491_17697 5.354286e+00
R35819 n0_20491_17697 n0_20679_17697 1.074286e+00
R35820 n0_241_17730 n0_429_17730 1.074286e+00
R35821 n0_429_17730 n0_1366_17730 5.354286e+00
R35822 n0_1366_17730 n0_1554_17730 1.074286e+00
R35823 n0_1554_17730 n0_2491_17730 5.354286e+00
R35824 n0_2491_17730 n0_2679_17730 1.074286e+00
R35825 n0_2679_17730 n0_3616_17730 5.354286e+00
R35826 n0_3616_17730 n0_3708_17730 5.257143e-01
R35827 n0_3708_17730 n0_3804_17730 5.485714e-01
R35828 n0_3804_17730 n0_3896_17730 5.257143e-01
R35829 n0_3896_17730 n0_5866_17730 1.125714e+01
R35830 n0_5866_17730 n0_5958_17730 5.257143e-01
R35831 n0_5958_17730 n0_6054_17730 5.485714e-01
R35832 n0_6054_17730 n0_6146_17730 5.257143e-01
R35833 n0_6146_17730 n0_8116_17730 1.125714e+01
R35834 n0_8116_17730 n0_8208_17730 5.257143e-01
R35835 n0_8208_17730 n0_8304_17730 5.485714e-01
R35836 n0_8304_17730 n0_8396_17730 5.257143e-01
R35837 n0_8396_17730 n0_10366_17730 1.125714e+01
R35838 n0_10366_17730 n0_10458_17730 5.257143e-01
R35839 n0_10458_17730 n0_10554_17730 5.485714e-01
R35840 n0_10554_17730 n0_10646_17730 5.257143e-01
R35841 n0_10646_17730 n0_12616_17730 1.125714e+01
R35842 n0_12616_17730 n0_12708_17730 5.257143e-01
R35843 n0_12708_17730 n0_12804_17730 5.485714e-01
R35844 n0_12804_17730 n0_12896_17730 5.257143e-01
R35845 n0_12896_17730 n0_14866_17730 1.125714e+01
R35846 n0_14866_17730 n0_14958_17730 5.257143e-01
R35847 n0_14958_17730 n0_15054_17730 5.485714e-01
R35848 n0_15054_17730 n0_15146_17730 5.257143e-01
R35849 n0_15146_17730 n0_17116_17730 1.125714e+01
R35850 n0_17116_17730 n0_17208_17730 5.257143e-01
R35851 n0_17208_17730 n0_17304_17730 5.485714e-01
R35852 n0_17304_17730 n0_17396_17730 5.257143e-01
R35853 n0_17396_17730 n0_18241_17730 4.828571e+00
R35854 n0_18241_17730 n0_18429_17730 1.074286e+00
R35855 n0_18429_17730 n0_19366_17730 5.354286e+00
R35856 n0_19366_17730 n0_19554_17730 1.074286e+00
R35857 n0_19554_17730 n0_20491_17730 5.354286e+00
R35858 n0_20491_17730 n0_20679_17730 1.074286e+00
R35859 n0_241_17913 n0_429_17913 1.074286e+00
R35860 n0_429_17913 n0_1366_17913 5.354286e+00
R35861 n0_1366_17913 n0_1554_17913 1.074286e+00
R35862 n0_1554_17913 n0_2491_17913 5.354286e+00
R35863 n0_2491_17913 n0_2679_17913 1.074286e+00
R35864 n0_2679_17913 n0_3616_17913 5.354286e+00
R35865 n0_3616_17913 n0_3708_17913 5.257143e-01
R35866 n0_3708_17913 n0_3804_17913 5.485714e-01
R35867 n0_3804_17913 n0_3896_17913 5.257143e-01
R35868 n0_3896_17913 n0_5866_17913 1.125714e+01
R35869 n0_5866_17913 n0_5958_17913 5.257143e-01
R35870 n0_5958_17913 n0_6054_17913 5.485714e-01
R35871 n0_6054_17913 n0_6146_17913 5.257143e-01
R35872 n0_6146_17913 n0_8116_17913 1.125714e+01
R35873 n0_8116_17913 n0_8208_17913 5.257143e-01
R35874 n0_8208_17913 n0_8304_17913 5.485714e-01
R35875 n0_8304_17913 n0_8396_17913 5.257143e-01
R35876 n0_8396_17913 n0_10366_17913 1.125714e+01
R35877 n0_10366_17913 n0_10458_17913 5.257143e-01
R35878 n0_10458_17913 n0_10554_17913 5.485714e-01
R35879 n0_10554_17913 n0_10646_17913 5.257143e-01
R35880 n0_10646_17913 n0_12616_17913 1.125714e+01
R35881 n0_12616_17913 n0_12708_17913 5.257143e-01
R35882 n0_12708_17913 n0_12804_17913 5.485714e-01
R35883 n0_12804_17913 n0_12896_17913 5.257143e-01
R35884 n0_12896_17913 n0_14866_17913 1.125714e+01
R35885 n0_14866_17913 n0_14958_17913 5.257143e-01
R35886 n0_14958_17913 n0_15054_17913 5.485714e-01
R35887 n0_15054_17913 n0_15146_17913 5.257143e-01
R35888 n0_15146_17913 n0_17116_17913 1.125714e+01
R35889 n0_17116_17913 n0_17208_17913 5.257143e-01
R35890 n0_17208_17913 n0_17304_17913 5.485714e-01
R35891 n0_17304_17913 n0_17396_17913 5.257143e-01
R35892 n0_17396_17913 n0_18241_17913 4.828571e+00
R35893 n0_18241_17913 n0_18429_17913 1.074286e+00
R35894 n0_18429_17913 n0_19366_17913 5.354286e+00
R35895 n0_19366_17913 n0_19554_17913 1.074286e+00
R35896 n0_19554_17913 n0_20491_17913 5.354286e+00
R35897 n0_20491_17913 n0_20679_17913 1.074286e+00
R35898 n0_241_17946 n0_429_17946 1.074286e+00
R35899 n0_429_17946 n0_1366_17946 5.354286e+00
R35900 n0_1366_17946 n0_1554_17946 1.074286e+00
R35901 n0_1554_17946 n0_2491_17946 5.354286e+00
R35902 n0_2491_17946 n0_2679_17946 1.074286e+00
R35903 n0_2679_17946 n0_3616_17946 5.354286e+00
R35904 n0_3616_17946 n0_3708_17946 5.257143e-01
R35905 n0_3708_17946 n0_3804_17946 5.485714e-01
R35906 n0_3804_17946 n0_3896_17946 5.257143e-01
R35907 n0_3896_17946 n0_5866_17946 1.125714e+01
R35908 n0_5866_17946 n0_5958_17946 5.257143e-01
R35909 n0_5958_17946 n0_6054_17946 5.485714e-01
R35910 n0_6054_17946 n0_6146_17946 5.257143e-01
R35911 n0_6146_17946 n0_8116_17946 1.125714e+01
R35912 n0_8116_17946 n0_8208_17946 5.257143e-01
R35913 n0_8208_17946 n0_8304_17946 5.485714e-01
R35914 n0_8304_17946 n0_8396_17946 5.257143e-01
R35915 n0_8396_17946 n0_10366_17946 1.125714e+01
R35916 n0_10366_17946 n0_10458_17946 5.257143e-01
R35917 n0_10458_17946 n0_10554_17946 5.485714e-01
R35918 n0_10554_17946 n0_10646_17946 5.257143e-01
R35919 n0_10646_17946 n0_12616_17946 1.125714e+01
R35920 n0_12616_17946 n0_12708_17946 5.257143e-01
R35921 n0_12708_17946 n0_12804_17946 5.485714e-01
R35922 n0_12804_17946 n0_12896_17946 5.257143e-01
R35923 n0_12896_17946 n0_14866_17946 1.125714e+01
R35924 n0_14866_17946 n0_14958_17946 5.257143e-01
R35925 n0_14958_17946 n0_15054_17946 5.485714e-01
R35926 n0_15054_17946 n0_15146_17946 5.257143e-01
R35927 n0_15146_17946 n0_17116_17946 1.125714e+01
R35928 n0_17116_17946 n0_17208_17946 5.257143e-01
R35929 n0_17208_17946 n0_17304_17946 5.485714e-01
R35930 n0_17304_17946 n0_17396_17946 5.257143e-01
R35931 n0_17396_17946 n0_18241_17946 4.828571e+00
R35932 n0_18241_17946 n0_18429_17946 1.074286e+00
R35933 n0_18429_17946 n0_19366_17946 5.354286e+00
R35934 n0_19366_17946 n0_19554_17946 1.074286e+00
R35935 n0_19554_17946 n0_20491_17946 5.354286e+00
R35936 n0_20491_17946 n0_20679_17946 1.074286e+00
R35937 n0_241_18129 n0_429_18129 1.074286e+00
R35938 n0_429_18129 n0_1366_18129 5.354286e+00
R35939 n0_1366_18129 n0_1554_18129 1.074286e+00
R35940 n0_1554_18129 n0_2491_18129 5.354286e+00
R35941 n0_2491_18129 n0_2679_18129 1.074286e+00
R35942 n0_2679_18129 n0_3616_18129 5.354286e+00
R35943 n0_3616_18129 n0_3708_18129 5.257143e-01
R35944 n0_3708_18129 n0_3804_18129 5.485714e-01
R35945 n0_3804_18129 n0_3896_18129 5.257143e-01
R35946 n0_3896_18129 n0_5866_18129 1.125714e+01
R35947 n0_5866_18129 n0_5958_18129 5.257143e-01
R35948 n0_5958_18129 n0_6054_18129 5.485714e-01
R35949 n0_6054_18129 n0_6146_18129 5.257143e-01
R35950 n0_6146_18129 n0_8116_18129 1.125714e+01
R35951 n0_8116_18129 n0_8208_18129 5.257143e-01
R35952 n0_8208_18129 n0_8304_18129 5.485714e-01
R35953 n0_8304_18129 n0_8396_18129 5.257143e-01
R35954 n0_8396_18129 n0_10366_18129 1.125714e+01
R35955 n0_10366_18129 n0_10458_18129 5.257143e-01
R35956 n0_10458_18129 n0_10554_18129 5.485714e-01
R35957 n0_10554_18129 n0_10646_18129 5.257143e-01
R35958 n0_10646_18129 n0_12616_18129 1.125714e+01
R35959 n0_12616_18129 n0_12708_18129 5.257143e-01
R35960 n0_12708_18129 n0_12804_18129 5.485714e-01
R35961 n0_12804_18129 n0_12896_18129 5.257143e-01
R35962 n0_12896_18129 n0_14866_18129 1.125714e+01
R35963 n0_14866_18129 n0_14958_18129 5.257143e-01
R35964 n0_14958_18129 n0_15054_18129 5.485714e-01
R35965 n0_15054_18129 n0_15146_18129 5.257143e-01
R35966 n0_15146_18129 n0_17116_18129 1.125714e+01
R35967 n0_17116_18129 n0_17208_18129 5.257143e-01
R35968 n0_17208_18129 n0_17304_18129 5.485714e-01
R35969 n0_17304_18129 n0_17396_18129 5.257143e-01
R35970 n0_17396_18129 n0_18241_18129 4.828571e+00
R35971 n0_18241_18129 n0_18429_18129 1.074286e+00
R35972 n0_18429_18129 n0_19366_18129 5.354286e+00
R35973 n0_19366_18129 n0_19554_18129 1.074286e+00
R35974 n0_19554_18129 n0_20491_18129 5.354286e+00
R35975 n0_20491_18129 n0_20679_18129 1.074286e+00
R35976 n0_241_18162 n0_429_18162 1.074286e+00
R35977 n0_429_18162 n0_1366_18162 5.354286e+00
R35978 n0_1366_18162 n0_1554_18162 1.074286e+00
R35979 n0_1554_18162 n0_2491_18162 5.354286e+00
R35980 n0_2491_18162 n0_2679_18162 1.074286e+00
R35981 n0_2679_18162 n0_3616_18162 5.354286e+00
R35982 n0_3616_18162 n0_3708_18162 5.257143e-01
R35983 n0_3708_18162 n0_3804_18162 5.485714e-01
R35984 n0_3804_18162 n0_3896_18162 5.257143e-01
R35985 n0_3896_18162 n0_5866_18162 1.125714e+01
R35986 n0_5866_18162 n0_5958_18162 5.257143e-01
R35987 n0_5958_18162 n0_6054_18162 5.485714e-01
R35988 n0_6054_18162 n0_6146_18162 5.257143e-01
R35989 n0_6146_18162 n0_8116_18162 1.125714e+01
R35990 n0_8116_18162 n0_8208_18162 5.257143e-01
R35991 n0_8208_18162 n0_8304_18162 5.485714e-01
R35992 n0_8304_18162 n0_8396_18162 5.257143e-01
R35993 n0_8396_18162 n0_10366_18162 1.125714e+01
R35994 n0_10366_18162 n0_10458_18162 5.257143e-01
R35995 n0_10458_18162 n0_10554_18162 5.485714e-01
R35996 n0_10554_18162 n0_10646_18162 5.257143e-01
R35997 n0_10646_18162 n0_12616_18162 1.125714e+01
R35998 n0_12616_18162 n0_12708_18162 5.257143e-01
R35999 n0_12708_18162 n0_12804_18162 5.485714e-01
R36000 n0_12804_18162 n0_12896_18162 5.257143e-01
R36001 n0_12896_18162 n0_14866_18162 1.125714e+01
R36002 n0_14866_18162 n0_14958_18162 5.257143e-01
R36003 n0_14958_18162 n0_15054_18162 5.485714e-01
R36004 n0_15054_18162 n0_15146_18162 5.257143e-01
R36005 n0_15146_18162 n0_17116_18162 1.125714e+01
R36006 n0_17116_18162 n0_17208_18162 5.257143e-01
R36007 n0_17208_18162 n0_17304_18162 5.485714e-01
R36008 n0_17304_18162 n0_17396_18162 5.257143e-01
R36009 n0_17396_18162 n0_18241_18162 4.828571e+00
R36010 n0_18241_18162 n0_18429_18162 1.074286e+00
R36011 n0_18429_18162 n0_19366_18162 5.354286e+00
R36012 n0_19366_18162 n0_19554_18162 1.074286e+00
R36013 n0_19554_18162 n0_20491_18162 5.354286e+00
R36014 n0_20491_18162 n0_20679_18162 1.074286e+00
R36015 n0_241_18345 n0_429_18345 1.074286e+00
R36016 n0_429_18345 n0_1366_18345 5.354286e+00
R36017 n0_1366_18345 n0_1554_18345 1.074286e+00
R36018 n0_1554_18345 n0_2491_18345 5.354286e+00
R36019 n0_2491_18345 n0_2679_18345 1.074286e+00
R36020 n0_2679_18345 n0_3616_18345 5.354286e+00
R36021 n0_3616_18345 n0_3708_18345 5.257143e-01
R36022 n0_3708_18345 n0_3804_18345 5.485714e-01
R36023 n0_3804_18345 n0_3896_18345 5.257143e-01
R36024 n0_3896_18345 n0_5866_18345 1.125714e+01
R36025 n0_5866_18345 n0_5958_18345 5.257143e-01
R36026 n0_5958_18345 n0_6054_18345 5.485714e-01
R36027 n0_6054_18345 n0_6146_18345 5.257143e-01
R36028 n0_6146_18345 n0_8116_18345 1.125714e+01
R36029 n0_8116_18345 n0_8208_18345 5.257143e-01
R36030 n0_8208_18345 n0_8304_18345 5.485714e-01
R36031 n0_8304_18345 n0_8396_18345 5.257143e-01
R36032 n0_8396_18345 n0_10366_18345 1.125714e+01
R36033 n0_10366_18345 n0_10458_18345 5.257143e-01
R36034 n0_10458_18345 n0_10554_18345 5.485714e-01
R36035 n0_10554_18345 n0_10646_18345 5.257143e-01
R36036 n0_10646_18345 n0_12616_18345 1.125714e+01
R36037 n0_12616_18345 n0_12708_18345 5.257143e-01
R36038 n0_12708_18345 n0_12804_18345 5.485714e-01
R36039 n0_12804_18345 n0_12896_18345 5.257143e-01
R36040 n0_12896_18345 n0_14866_18345 1.125714e+01
R36041 n0_14866_18345 n0_14958_18345 5.257143e-01
R36042 n0_14958_18345 n0_15054_18345 5.485714e-01
R36043 n0_15054_18345 n0_15146_18345 5.257143e-01
R36044 n0_15146_18345 n0_17116_18345 1.125714e+01
R36045 n0_17116_18345 n0_17208_18345 5.257143e-01
R36046 n0_17208_18345 n0_17304_18345 5.485714e-01
R36047 n0_17304_18345 n0_17396_18345 5.257143e-01
R36048 n0_17396_18345 n0_18241_18345 4.828571e+00
R36049 n0_18241_18345 n0_18429_18345 1.074286e+00
R36050 n0_18429_18345 n0_19366_18345 5.354286e+00
R36051 n0_19366_18345 n0_19554_18345 1.074286e+00
R36052 n0_19554_18345 n0_20491_18345 5.354286e+00
R36053 n0_20491_18345 n0_20679_18345 1.074286e+00
R36054 n0_241_18378 n0_1366_18378 6.428571e+00
R36055 n0_1366_18378 n0_2491_18378 6.428571e+00
R36056 n0_2491_18378 n0_3616_18378 6.428571e+00
R36057 n0_3616_18378 n0_3708_18378 5.257143e-01
R36058 n0_3708_18378 n0_3804_18378 5.485714e-01
R36059 n0_3804_18378 n0_3896_18378 5.257143e-01
R36060 n0_3896_18378 n0_5866_18378 1.125714e+01
R36061 n0_5866_18378 n0_5958_18378 5.257143e-01
R36062 n0_5958_18378 n0_6054_18378 5.485714e-01
R36063 n0_6054_18378 n0_6146_18378 5.257143e-01
R36064 n0_6146_18378 n0_8116_18378 1.125714e+01
R36065 n0_8116_18378 n0_8208_18378 5.257143e-01
R36066 n0_8208_18378 n0_8304_18378 5.485714e-01
R36067 n0_8304_18378 n0_8396_18378 5.257143e-01
R36068 n0_8396_18378 n0_10366_18378 1.125714e+01
R36069 n0_10366_18378 n0_10458_18378 5.257143e-01
R36070 n0_10458_18378 n0_10554_18378 5.485714e-01
R36071 n0_10554_18378 n0_10646_18378 5.257143e-01
R36072 n0_10646_18378 n0_12616_18378 1.125714e+01
R36073 n0_12616_18378 n0_12708_18378 5.257143e-01
R36074 n0_12708_18378 n0_12804_18378 5.485714e-01
R36075 n0_12804_18378 n0_12896_18378 5.257143e-01
R36076 n0_12896_18378 n0_14866_18378 1.125714e+01
R36077 n0_14866_18378 n0_14958_18378 5.257143e-01
R36078 n0_14958_18378 n0_15054_18378 5.485714e-01
R36079 n0_15054_18378 n0_15146_18378 5.257143e-01
R36080 n0_15146_18378 n0_17116_18378 1.125714e+01
R36081 n0_17116_18378 n0_17208_18378 5.257143e-01
R36082 n0_17208_18378 n0_17304_18378 5.485714e-01
R36083 n0_17304_18378 n0_17396_18378 5.257143e-01
R36084 n0_17396_18378 n0_18241_18378 4.828571e+00
R36085 n0_18241_18378 n0_19366_18378 6.428571e+00
R36086 n0_19366_18378 n0_20491_18378 6.428571e+00
R36087 n0_241_18561 n0_1366_18561 6.428571e+00
R36088 n0_1366_18561 n0_3616_18561 1.285714e+01
R36089 n0_3616_18561 n0_3708_18561 5.257143e-01
R36090 n0_3708_18561 n0_3804_18561 5.485714e-01
R36091 n0_3804_18561 n0_3896_18561 5.257143e-01
R36092 n0_3896_18561 n0_5866_18561 1.125714e+01
R36093 n0_5866_18561 n0_5958_18561 5.257143e-01
R36094 n0_5958_18561 n0_6054_18561 5.485714e-01
R36095 n0_6054_18561 n0_6146_18561 5.257143e-01
R36096 n0_6146_18561 n0_8116_18561 1.125714e+01
R36097 n0_8116_18561 n0_8208_18561 5.257143e-01
R36098 n0_8208_18561 n0_8304_18561 5.485714e-01
R36099 n0_8304_18561 n0_8396_18561 5.257143e-01
R36100 n0_8396_18561 n0_10366_18561 1.125714e+01
R36101 n0_10366_18561 n0_10458_18561 5.257143e-01
R36102 n0_10458_18561 n0_10554_18561 5.485714e-01
R36103 n0_10554_18561 n0_10646_18561 5.257143e-01
R36104 n0_10646_18561 n0_12616_18561 1.125714e+01
R36105 n0_12616_18561 n0_12708_18561 5.257143e-01
R36106 n0_12708_18561 n0_12804_18561 5.485714e-01
R36107 n0_12804_18561 n0_12896_18561 5.257143e-01
R36108 n0_12896_18561 n0_14866_18561 1.125714e+01
R36109 n0_14866_18561 n0_14958_18561 5.257143e-01
R36110 n0_14958_18561 n0_15054_18561 5.485714e-01
R36111 n0_15054_18561 n0_15146_18561 5.257143e-01
R36112 n0_15146_18561 n0_17116_18561 1.125714e+01
R36113 n0_17116_18561 n0_17208_18561 5.257143e-01
R36114 n0_17208_18561 n0_17304_18561 5.485714e-01
R36115 n0_17304_18561 n0_17396_18561 5.257143e-01
R36116 n0_17396_18561 n0_19366_18561 1.125714e+01
R36117 n0_19366_18561 n0_20491_18561 6.428571e+00
R36118 n0_241_18594 n0_429_18594 1.074286e+00
R36119 n0_429_18594 n0_1366_18594 5.354286e+00
R36120 n0_1366_18594 n0_1554_18594 1.074286e+00
R36121 n0_1554_18594 n0_3616_18594 1.178286e+01
R36122 n0_3616_18594 n0_3708_18594 5.257143e-01
R36123 n0_3708_18594 n0_3804_18594 5.485714e-01
R36124 n0_3804_18594 n0_3896_18594 5.257143e-01
R36125 n0_3896_18594 n0_5866_18594 1.125714e+01
R36126 n0_5866_18594 n0_5958_18594 5.257143e-01
R36127 n0_5958_18594 n0_6054_18594 5.485714e-01
R36128 n0_6054_18594 n0_6146_18594 5.257143e-01
R36129 n0_6146_18594 n0_8116_18594 1.125714e+01
R36130 n0_8116_18594 n0_8208_18594 5.257143e-01
R36131 n0_8208_18594 n0_8304_18594 5.485714e-01
R36132 n0_8304_18594 n0_8396_18594 5.257143e-01
R36133 n0_8396_18594 n0_10366_18594 1.125714e+01
R36134 n0_10366_18594 n0_10458_18594 5.257143e-01
R36135 n0_10458_18594 n0_10554_18594 5.485714e-01
R36136 n0_10554_18594 n0_10646_18594 5.257143e-01
R36137 n0_10646_18594 n0_12616_18594 1.125714e+01
R36138 n0_12616_18594 n0_12708_18594 5.257143e-01
R36139 n0_12708_18594 n0_12804_18594 5.485714e-01
R36140 n0_12804_18594 n0_12896_18594 5.257143e-01
R36141 n0_12896_18594 n0_14866_18594 1.125714e+01
R36142 n0_14866_18594 n0_14958_18594 5.257143e-01
R36143 n0_14958_18594 n0_15054_18594 5.485714e-01
R36144 n0_15054_18594 n0_15146_18594 5.257143e-01
R36145 n0_15146_18594 n0_17116_18594 1.125714e+01
R36146 n0_17116_18594 n0_17208_18594 5.257143e-01
R36147 n0_17208_18594 n0_17304_18594 5.485714e-01
R36148 n0_17304_18594 n0_17396_18594 5.257143e-01
R36149 n0_17396_18594 n0_19366_18594 1.125714e+01
R36150 n0_19366_18594 n0_19554_18594 1.074286e+00
R36151 n0_19554_18594 n0_20491_18594 5.354286e+00
R36152 n0_20491_18594 n0_20679_18594 1.074286e+00
R36153 n0_241_18777 n0_429_18777 1.074286e+00
R36154 n0_429_18777 n0_1366_18777 5.354286e+00
R36155 n0_1366_18777 n0_1554_18777 1.074286e+00
R36156 n0_1554_18777 n0_3616_18777 1.178286e+01
R36157 n0_3616_18777 n0_3708_18777 5.257143e-01
R36158 n0_3708_18777 n0_3804_18777 5.485714e-01
R36159 n0_3804_18777 n0_3896_18777 5.257143e-01
R36160 n0_3896_18777 n0_5866_18777 1.125714e+01
R36161 n0_5866_18777 n0_5958_18777 5.257143e-01
R36162 n0_5958_18777 n0_6054_18777 5.485714e-01
R36163 n0_6054_18777 n0_6146_18777 5.257143e-01
R36164 n0_6146_18777 n0_8116_18777 1.125714e+01
R36165 n0_8116_18777 n0_8208_18777 5.257143e-01
R36166 n0_8208_18777 n0_8304_18777 5.485714e-01
R36167 n0_8304_18777 n0_8396_18777 5.257143e-01
R36168 n0_8396_18777 n0_10366_18777 1.125714e+01
R36169 n0_10366_18777 n0_10458_18777 5.257143e-01
R36170 n0_10458_18777 n0_10554_18777 5.485714e-01
R36171 n0_10554_18777 n0_10646_18777 5.257143e-01
R36172 n0_10646_18777 n0_12616_18777 1.125714e+01
R36173 n0_12616_18777 n0_12708_18777 5.257143e-01
R36174 n0_12708_18777 n0_12804_18777 5.485714e-01
R36175 n0_12804_18777 n0_12896_18777 5.257143e-01
R36176 n0_12896_18777 n0_14866_18777 1.125714e+01
R36177 n0_14866_18777 n0_14958_18777 5.257143e-01
R36178 n0_14958_18777 n0_15054_18777 5.485714e-01
R36179 n0_15054_18777 n0_15146_18777 5.257143e-01
R36180 n0_15146_18777 n0_17116_18777 1.125714e+01
R36181 n0_17116_18777 n0_17208_18777 5.257143e-01
R36182 n0_17208_18777 n0_17304_18777 5.485714e-01
R36183 n0_17304_18777 n0_17396_18777 5.257143e-01
R36184 n0_17396_18777 n0_19366_18777 1.125714e+01
R36185 n0_19366_18777 n0_19554_18777 1.074286e+00
R36186 n0_19554_18777 n0_20491_18777 5.354286e+00
R36187 n0_20491_18777 n0_20679_18777 1.074286e+00
R36188 n0_241_18810 n0_429_18810 1.074286e+00
R36189 n0_429_18810 n0_1366_18810 5.354286e+00
R36190 n0_1366_18810 n0_1554_18810 1.074286e+00
R36191 n0_1554_18810 n0_3616_18810 1.178286e+01
R36192 n0_3616_18810 n0_3708_18810 5.257143e-01
R36193 n0_3708_18810 n0_3804_18810 5.485714e-01
R36194 n0_3804_18810 n0_3896_18810 5.257143e-01
R36195 n0_3896_18810 n0_5866_18810 1.125714e+01
R36196 n0_5866_18810 n0_5958_18810 5.257143e-01
R36197 n0_5958_18810 n0_6054_18810 5.485714e-01
R36198 n0_6054_18810 n0_6146_18810 5.257143e-01
R36199 n0_6146_18810 n0_8116_18810 1.125714e+01
R36200 n0_8116_18810 n0_8208_18810 5.257143e-01
R36201 n0_8208_18810 n0_8304_18810 5.485714e-01
R36202 n0_8304_18810 n0_8396_18810 5.257143e-01
R36203 n0_8396_18810 n0_10366_18810 1.125714e+01
R36204 n0_10366_18810 n0_10458_18810 5.257143e-01
R36205 n0_10458_18810 n0_10554_18810 5.485714e-01
R36206 n0_10554_18810 n0_10646_18810 5.257143e-01
R36207 n0_10646_18810 n0_12616_18810 1.125714e+01
R36208 n0_12616_18810 n0_12708_18810 5.257143e-01
R36209 n0_12708_18810 n0_12804_18810 5.485714e-01
R36210 n0_12804_18810 n0_12896_18810 5.257143e-01
R36211 n0_12896_18810 n0_14866_18810 1.125714e+01
R36212 n0_14866_18810 n0_14958_18810 5.257143e-01
R36213 n0_14958_18810 n0_15054_18810 5.485714e-01
R36214 n0_15054_18810 n0_15146_18810 5.257143e-01
R36215 n0_15146_18810 n0_17116_18810 1.125714e+01
R36216 n0_17116_18810 n0_17208_18810 5.257143e-01
R36217 n0_17208_18810 n0_17304_18810 5.485714e-01
R36218 n0_17304_18810 n0_17396_18810 5.257143e-01
R36219 n0_17396_18810 n0_19366_18810 1.125714e+01
R36220 n0_19366_18810 n0_19554_18810 1.074286e+00
R36221 n0_19554_18810 n0_20491_18810 5.354286e+00
R36222 n0_20491_18810 n0_20679_18810 1.074286e+00
R36223 n0_241_18993 n0_429_18993 1.074286e+00
R36224 n0_429_18993 n0_1366_18993 5.354286e+00
R36225 n0_1366_18993 n0_1554_18993 1.074286e+00
R36226 n0_1554_18993 n0_3616_18993 1.178286e+01
R36227 n0_3616_18993 n0_3708_18993 5.257143e-01
R36228 n0_3708_18993 n0_3804_18993 5.485714e-01
R36229 n0_3804_18993 n0_3896_18993 5.257143e-01
R36230 n0_3896_18993 n0_5866_18993 1.125714e+01
R36231 n0_5866_18993 n0_5958_18993 5.257143e-01
R36232 n0_5958_18993 n0_6054_18993 5.485714e-01
R36233 n0_6054_18993 n0_6146_18993 5.257143e-01
R36234 n0_6146_18993 n0_8116_18993 1.125714e+01
R36235 n0_8116_18993 n0_8208_18993 5.257143e-01
R36236 n0_8208_18993 n0_8304_18993 5.485714e-01
R36237 n0_8304_18993 n0_8396_18993 5.257143e-01
R36238 n0_8396_18993 n0_10366_18993 1.125714e+01
R36239 n0_10366_18993 n0_10458_18993 5.257143e-01
R36240 n0_10458_18993 n0_10554_18993 5.485714e-01
R36241 n0_10554_18993 n0_10646_18993 5.257143e-01
R36242 n0_10646_18993 n0_12616_18993 1.125714e+01
R36243 n0_12616_18993 n0_12708_18993 5.257143e-01
R36244 n0_12708_18993 n0_12804_18993 5.485714e-01
R36245 n0_12804_18993 n0_12896_18993 5.257143e-01
R36246 n0_12896_18993 n0_14866_18993 1.125714e+01
R36247 n0_14866_18993 n0_14958_18993 5.257143e-01
R36248 n0_14958_18993 n0_15054_18993 5.485714e-01
R36249 n0_15054_18993 n0_15146_18993 5.257143e-01
R36250 n0_15146_18993 n0_17116_18993 1.125714e+01
R36251 n0_17116_18993 n0_17208_18993 5.257143e-01
R36252 n0_17208_18993 n0_17304_18993 5.485714e-01
R36253 n0_17304_18993 n0_17396_18993 5.257143e-01
R36254 n0_17396_18993 n0_19366_18993 1.125714e+01
R36255 n0_19366_18993 n0_19554_18993 1.074286e+00
R36256 n0_19554_18993 n0_20491_18993 5.354286e+00
R36257 n0_20491_18993 n0_20679_18993 1.074286e+00
R36258 n0_241_19026 n0_429_19026 1.074286e+00
R36259 n0_429_19026 n0_1366_19026 5.354286e+00
R36260 n0_1366_19026 n0_1554_19026 1.074286e+00
R36261 n0_1554_19026 n0_3616_19026 1.178286e+01
R36262 n0_3616_19026 n0_3708_19026 5.257143e-01
R36263 n0_3708_19026 n0_3804_19026 5.485714e-01
R36264 n0_3804_19026 n0_3896_19026 5.257143e-01
R36265 n0_3896_19026 n0_5866_19026 1.125714e+01
R36266 n0_5866_19026 n0_5958_19026 5.257143e-01
R36267 n0_5958_19026 n0_6054_19026 5.485714e-01
R36268 n0_6054_19026 n0_6146_19026 5.257143e-01
R36269 n0_6146_19026 n0_8116_19026 1.125714e+01
R36270 n0_8116_19026 n0_8208_19026 5.257143e-01
R36271 n0_8208_19026 n0_8304_19026 5.485714e-01
R36272 n0_8304_19026 n0_8396_19026 5.257143e-01
R36273 n0_8396_19026 n0_10366_19026 1.125714e+01
R36274 n0_10366_19026 n0_10458_19026 5.257143e-01
R36275 n0_10458_19026 n0_10554_19026 5.485714e-01
R36276 n0_10554_19026 n0_10646_19026 5.257143e-01
R36277 n0_10646_19026 n0_12616_19026 1.125714e+01
R36278 n0_12616_19026 n0_12708_19026 5.257143e-01
R36279 n0_12708_19026 n0_12804_19026 5.485714e-01
R36280 n0_12804_19026 n0_12896_19026 5.257143e-01
R36281 n0_12896_19026 n0_14866_19026 1.125714e+01
R36282 n0_14866_19026 n0_14958_19026 5.257143e-01
R36283 n0_14958_19026 n0_15054_19026 5.485714e-01
R36284 n0_15054_19026 n0_15146_19026 5.257143e-01
R36285 n0_15146_19026 n0_17116_19026 1.125714e+01
R36286 n0_17116_19026 n0_17208_19026 5.257143e-01
R36287 n0_17208_19026 n0_17304_19026 5.485714e-01
R36288 n0_17304_19026 n0_17396_19026 5.257143e-01
R36289 n0_17396_19026 n0_19366_19026 1.125714e+01
R36290 n0_19366_19026 n0_19554_19026 1.074286e+00
R36291 n0_19554_19026 n0_20491_19026 5.354286e+00
R36292 n0_20491_19026 n0_20679_19026 1.074286e+00
R36293 n0_241_19209 n0_429_19209 1.074286e+00
R36294 n0_429_19209 n0_1366_19209 5.354286e+00
R36295 n0_1366_19209 n0_1554_19209 1.074286e+00
R36296 n0_1554_19209 n0_3616_19209 1.178286e+01
R36297 n0_3616_19209 n0_3708_19209 5.257143e-01
R36298 n0_3708_19209 n0_3804_19209 5.485714e-01
R36299 n0_3804_19209 n0_3896_19209 5.257143e-01
R36300 n0_3896_19209 n0_5866_19209 1.125714e+01
R36301 n0_5866_19209 n0_5958_19209 5.257143e-01
R36302 n0_5958_19209 n0_6054_19209 5.485714e-01
R36303 n0_6054_19209 n0_6146_19209 5.257143e-01
R36304 n0_6146_19209 n0_8116_19209 1.125714e+01
R36305 n0_8116_19209 n0_8208_19209 5.257143e-01
R36306 n0_8208_19209 n0_8304_19209 5.485714e-01
R36307 n0_8304_19209 n0_8396_19209 5.257143e-01
R36308 n0_8396_19209 n0_10366_19209 1.125714e+01
R36309 n0_10366_19209 n0_10458_19209 5.257143e-01
R36310 n0_10458_19209 n0_10554_19209 5.485714e-01
R36311 n0_10554_19209 n0_10646_19209 5.257143e-01
R36312 n0_10646_19209 n0_12616_19209 1.125714e+01
R36313 n0_12616_19209 n0_12708_19209 5.257143e-01
R36314 n0_12708_19209 n0_12804_19209 5.485714e-01
R36315 n0_12804_19209 n0_12896_19209 5.257143e-01
R36316 n0_12896_19209 n0_14866_19209 1.125714e+01
R36317 n0_14866_19209 n0_14958_19209 5.257143e-01
R36318 n0_14958_19209 n0_15054_19209 5.485714e-01
R36319 n0_15054_19209 n0_15146_19209 5.257143e-01
R36320 n0_15146_19209 n0_17116_19209 1.125714e+01
R36321 n0_17116_19209 n0_17208_19209 5.257143e-01
R36322 n0_17208_19209 n0_17304_19209 5.485714e-01
R36323 n0_17304_19209 n0_17396_19209 5.257143e-01
R36324 n0_17396_19209 n0_19366_19209 1.125714e+01
R36325 n0_19366_19209 n0_19554_19209 1.074286e+00
R36326 n0_19554_19209 n0_20491_19209 5.354286e+00
R36327 n0_20491_19209 n0_20679_19209 1.074286e+00
R36328 n0_241_19242 n0_429_19242 1.074286e+00
R36329 n0_429_19242 n0_1366_19242 5.354286e+00
R36330 n0_1366_19242 n0_1554_19242 1.074286e+00
R36331 n0_1554_19242 n0_3616_19242 1.178286e+01
R36332 n0_3616_19242 n0_3708_19242 5.257143e-01
R36333 n0_3708_19242 n0_3804_19242 5.485714e-01
R36334 n0_3804_19242 n0_3896_19242 5.257143e-01
R36335 n0_3896_19242 n0_5866_19242 1.125714e+01
R36336 n0_5866_19242 n0_5958_19242 5.257143e-01
R36337 n0_5958_19242 n0_6054_19242 5.485714e-01
R36338 n0_6054_19242 n0_6146_19242 5.257143e-01
R36339 n0_6146_19242 n0_8116_19242 1.125714e+01
R36340 n0_8116_19242 n0_8208_19242 5.257143e-01
R36341 n0_8208_19242 n0_8304_19242 5.485714e-01
R36342 n0_8304_19242 n0_8396_19242 5.257143e-01
R36343 n0_8396_19242 n0_10366_19242 1.125714e+01
R36344 n0_10366_19242 n0_10458_19242 5.257143e-01
R36345 n0_10458_19242 n0_10554_19242 5.485714e-01
R36346 n0_10554_19242 n0_10646_19242 5.257143e-01
R36347 n0_10646_19242 n0_12616_19242 1.125714e+01
R36348 n0_12616_19242 n0_12708_19242 5.257143e-01
R36349 n0_12708_19242 n0_12804_19242 5.485714e-01
R36350 n0_12804_19242 n0_12896_19242 5.257143e-01
R36351 n0_12896_19242 n0_14866_19242 1.125714e+01
R36352 n0_14866_19242 n0_14958_19242 5.257143e-01
R36353 n0_14958_19242 n0_15054_19242 5.485714e-01
R36354 n0_15054_19242 n0_15146_19242 5.257143e-01
R36355 n0_15146_19242 n0_17116_19242 1.125714e+01
R36356 n0_17116_19242 n0_17208_19242 5.257143e-01
R36357 n0_17208_19242 n0_17304_19242 5.485714e-01
R36358 n0_17304_19242 n0_17396_19242 5.257143e-01
R36359 n0_17396_19242 n0_19366_19242 1.125714e+01
R36360 n0_19366_19242 n0_19554_19242 1.074286e+00
R36361 n0_19554_19242 n0_20491_19242 5.354286e+00
R36362 n0_20491_19242 n0_20679_19242 1.074286e+00
R36363 n0_241_19425 n0_429_19425 1.074286e+00
R36364 n0_429_19425 n0_1366_19425 5.354286e+00
R36365 n0_1366_19425 n0_1554_19425 1.074286e+00
R36366 n0_1554_19425 n0_3616_19425 1.178286e+01
R36367 n0_3616_19425 n0_3708_19425 5.257143e-01
R36368 n0_3708_19425 n0_3804_19425 5.485714e-01
R36369 n0_3804_19425 n0_3896_19425 5.257143e-01
R36370 n0_3896_19425 n0_5866_19425 1.125714e+01
R36371 n0_5866_19425 n0_5958_19425 5.257143e-01
R36372 n0_5958_19425 n0_6054_19425 5.485714e-01
R36373 n0_6054_19425 n0_6146_19425 5.257143e-01
R36374 n0_6146_19425 n0_8116_19425 1.125714e+01
R36375 n0_8116_19425 n0_8208_19425 5.257143e-01
R36376 n0_8208_19425 n0_8304_19425 5.485714e-01
R36377 n0_8304_19425 n0_8396_19425 5.257143e-01
R36378 n0_8396_19425 n0_10366_19425 1.125714e+01
R36379 n0_10366_19425 n0_10458_19425 5.257143e-01
R36380 n0_10458_19425 n0_10554_19425 5.485714e-01
R36381 n0_10554_19425 n0_10646_19425 5.257143e-01
R36382 n0_10646_19425 n0_12616_19425 1.125714e+01
R36383 n0_12616_19425 n0_12708_19425 5.257143e-01
R36384 n0_12708_19425 n0_12804_19425 5.485714e-01
R36385 n0_12804_19425 n0_12896_19425 5.257143e-01
R36386 n0_12896_19425 n0_14866_19425 1.125714e+01
R36387 n0_14866_19425 n0_14958_19425 5.257143e-01
R36388 n0_14958_19425 n0_15054_19425 5.485714e-01
R36389 n0_15054_19425 n0_15146_19425 5.257143e-01
R36390 n0_15146_19425 n0_17116_19425 1.125714e+01
R36391 n0_17116_19425 n0_17208_19425 5.257143e-01
R36392 n0_17208_19425 n0_17304_19425 5.485714e-01
R36393 n0_17304_19425 n0_17396_19425 5.257143e-01
R36394 n0_17396_19425 n0_19366_19425 1.125714e+01
R36395 n0_19366_19425 n0_19554_19425 1.074286e+00
R36396 n0_19554_19425 n0_20491_19425 5.354286e+00
R36397 n0_20491_19425 n0_20679_19425 1.074286e+00
R36398 n0_241_19458 n0_429_19458 1.074286e+00
R36399 n0_429_19458 n0_1366_19458 5.354286e+00
R36400 n0_1366_19458 n0_1554_19458 1.074286e+00
R36401 n0_1554_19458 n0_3616_19458 1.178286e+01
R36402 n0_3616_19458 n0_3708_19458 5.257143e-01
R36403 n0_3708_19458 n0_3804_19458 5.485714e-01
R36404 n0_3804_19458 n0_3896_19458 5.257143e-01
R36405 n0_3896_19458 n0_5866_19458 1.125714e+01
R36406 n0_5866_19458 n0_5958_19458 5.257143e-01
R36407 n0_5958_19458 n0_6054_19458 5.485714e-01
R36408 n0_6054_19458 n0_6146_19458 5.257143e-01
R36409 n0_6146_19458 n0_8116_19458 1.125714e+01
R36410 n0_8116_19458 n0_8208_19458 5.257143e-01
R36411 n0_8208_19458 n0_8304_19458 5.485714e-01
R36412 n0_8304_19458 n0_8396_19458 5.257143e-01
R36413 n0_8396_19458 n0_10366_19458 1.125714e+01
R36414 n0_10366_19458 n0_10458_19458 5.257143e-01
R36415 n0_10458_19458 n0_10554_19458 5.485714e-01
R36416 n0_10554_19458 n0_10646_19458 5.257143e-01
R36417 n0_10646_19458 n0_12616_19458 1.125714e+01
R36418 n0_12616_19458 n0_12708_19458 5.257143e-01
R36419 n0_12708_19458 n0_12804_19458 5.485714e-01
R36420 n0_12804_19458 n0_12896_19458 5.257143e-01
R36421 n0_12896_19458 n0_14866_19458 1.125714e+01
R36422 n0_14866_19458 n0_14958_19458 5.257143e-01
R36423 n0_14958_19458 n0_15054_19458 5.485714e-01
R36424 n0_15054_19458 n0_15146_19458 5.257143e-01
R36425 n0_15146_19458 n0_17116_19458 1.125714e+01
R36426 n0_17116_19458 n0_17208_19458 5.257143e-01
R36427 n0_17208_19458 n0_17304_19458 5.485714e-01
R36428 n0_17304_19458 n0_17396_19458 5.257143e-01
R36429 n0_17396_19458 n0_19366_19458 1.125714e+01
R36430 n0_19366_19458 n0_19554_19458 1.074286e+00
R36431 n0_19554_19458 n0_20491_19458 5.354286e+00
R36432 n0_20491_19458 n0_20679_19458 1.074286e+00
R36433 n0_241_19641 n0_380_19641 7.942857e-01
R36434 n0_380_19641 n0_429_19641 2.800000e-01
R36435 n0_429_19641 n0_1366_19641 5.354286e+00
R36436 n0_1366_19641 n0_1646_19641 1.600000e+00
R36437 n0_1646_19641 n0_3616_19641 1.125714e+01
R36438 n0_3616_19641 n0_3708_19641 5.257143e-01
R36439 n0_3708_19641 n0_3755_19641 2.685714e-01
R36440 n0_3755_19641 n0_3804_19641 2.800000e-01
R36441 n0_3804_19641 n0_3896_19641 5.257143e-01
R36442 n0_3896_19641 n0_5866_19641 1.125714e+01
R36443 n0_5866_19641 n0_5958_19641 5.257143e-01
R36444 n0_5958_19641 n0_6005_19641 2.685714e-01
R36445 n0_6005_19641 n0_6054_19641 2.800000e-01
R36446 n0_6054_19641 n0_6146_19641 5.257143e-01
R36447 n0_6146_19641 n0_8116_19641 1.125714e+01
R36448 n0_8116_19641 n0_8208_19641 5.257143e-01
R36449 n0_8208_19641 n0_8255_19641 2.685714e-01
R36450 n0_8255_19641 n0_8304_19641 2.800000e-01
R36451 n0_8304_19641 n0_8396_19641 5.257143e-01
R36452 n0_8396_19641 n0_10366_19641 1.125714e+01
R36453 n0_10366_19641 n0_10458_19641 5.257143e-01
R36454 n0_10458_19641 n0_10505_19641 2.685714e-01
R36455 n0_10505_19641 n0_10554_19641 2.800000e-01
R36456 n0_10554_19641 n0_10646_19641 5.257143e-01
R36457 n0_10646_19641 n0_12616_19641 1.125714e+01
R36458 n0_12616_19641 n0_12708_19641 5.257143e-01
R36459 n0_12708_19641 n0_12755_19641 2.685714e-01
R36460 n0_12755_19641 n0_12804_19641 2.800000e-01
R36461 n0_12804_19641 n0_12896_19641 5.257143e-01
R36462 n0_12896_19641 n0_14866_19641 1.125714e+01
R36463 n0_14866_19641 n0_14958_19641 5.257143e-01
R36464 n0_14958_19641 n0_15005_19641 2.685714e-01
R36465 n0_15005_19641 n0_15054_19641 2.800000e-01
R36466 n0_15054_19641 n0_15146_19641 5.257143e-01
R36467 n0_15146_19641 n0_17116_19641 1.125714e+01
R36468 n0_17116_19641 n0_17208_19641 5.257143e-01
R36469 n0_17208_19641 n0_17255_19641 2.685714e-01
R36470 n0_17255_19641 n0_17304_19641 2.800000e-01
R36471 n0_17304_19641 n0_17396_19641 5.257143e-01
R36472 n0_17396_19641 n0_19366_19641 1.125714e+01
R36473 n0_19366_19641 n0_19646_19641 1.600000e+00
R36474 n0_19646_19641 n0_20491_19641 4.828571e+00
R36475 n0_20491_19641 n0_20630_19641 7.942857e-01
R36476 n0_20630_19641 n0_20679_19641 2.800000e-01
R36477 n0_241_19674 n0_380_19674 7.942857e-01
R36478 n0_380_19674 n0_429_19674 2.800000e-01
R36479 n0_429_19674 n0_1366_19674 5.354286e+00
R36480 n0_1366_19674 n0_1646_19674 1.600000e+00
R36481 n0_1646_19674 n0_3616_19674 1.125714e+01
R36482 n0_3616_19674 n0_3708_19674 5.257143e-01
R36483 n0_3708_19674 n0_3755_19674 2.685714e-01
R36484 n0_3755_19674 n0_3804_19674 2.800000e-01
R36485 n0_3804_19674 n0_3896_19674 5.257143e-01
R36486 n0_3896_19674 n0_5866_19674 1.125714e+01
R36487 n0_5866_19674 n0_5958_19674 5.257143e-01
R36488 n0_5958_19674 n0_6005_19674 2.685714e-01
R36489 n0_6005_19674 n0_6054_19674 2.800000e-01
R36490 n0_6054_19674 n0_6146_19674 5.257143e-01
R36491 n0_6146_19674 n0_8116_19674 1.125714e+01
R36492 n0_8116_19674 n0_8208_19674 5.257143e-01
R36493 n0_8208_19674 n0_8255_19674 2.685714e-01
R36494 n0_8255_19674 n0_8304_19674 2.800000e-01
R36495 n0_8304_19674 n0_8396_19674 5.257143e-01
R36496 n0_8396_19674 n0_10366_19674 1.125714e+01
R36497 n0_10366_19674 n0_10458_19674 5.257143e-01
R36498 n0_10458_19674 n0_10505_19674 2.685714e-01
R36499 n0_10505_19674 n0_10554_19674 2.800000e-01
R36500 n0_10554_19674 n0_10646_19674 5.257143e-01
R36501 n0_10646_19674 n0_12616_19674 1.125714e+01
R36502 n0_12616_19674 n0_12708_19674 5.257143e-01
R36503 n0_12708_19674 n0_12755_19674 2.685714e-01
R36504 n0_12755_19674 n0_12804_19674 2.800000e-01
R36505 n0_12804_19674 n0_12896_19674 5.257143e-01
R36506 n0_12896_19674 n0_14866_19674 1.125714e+01
R36507 n0_14866_19674 n0_14958_19674 5.257143e-01
R36508 n0_14958_19674 n0_15005_19674 2.685714e-01
R36509 n0_15005_19674 n0_15054_19674 2.800000e-01
R36510 n0_15054_19674 n0_15146_19674 5.257143e-01
R36511 n0_15146_19674 n0_17116_19674 1.125714e+01
R36512 n0_17116_19674 n0_17208_19674 5.257143e-01
R36513 n0_17208_19674 n0_17255_19674 2.685714e-01
R36514 n0_17255_19674 n0_17304_19674 2.800000e-01
R36515 n0_17304_19674 n0_17396_19674 5.257143e-01
R36516 n0_17396_19674 n0_19366_19674 1.125714e+01
R36517 n0_19366_19674 n0_19646_19674 1.600000e+00
R36518 n0_19646_19674 n0_20491_19674 4.828571e+00
R36519 n0_20491_19674 n0_20630_19674 7.942857e-01
R36520 n0_20630_19674 n0_20679_19674 2.800000e-01
R36521 n0_241_19857 n0_429_19857 1.074286e+00
R36522 n0_429_19857 n0_1366_19857 5.354286e+00
R36523 n0_1366_19857 n0_1458_19857 5.257143e-01
R36524 n0_1458_19857 n0_1554_19857 5.485714e-01
R36525 n0_1554_19857 n0_1646_19857 5.257143e-01
R36526 n0_1646_19857 n0_3616_19857 1.125714e+01
R36527 n0_3616_19857 n0_3708_19857 5.257143e-01
R36528 n0_3708_19857 n0_3804_19857 5.485714e-01
R36529 n0_3804_19857 n0_3896_19857 5.257143e-01
R36530 n0_3896_19857 n0_5866_19857 1.125714e+01
R36531 n0_5866_19857 n0_5958_19857 5.257143e-01
R36532 n0_5958_19857 n0_6054_19857 5.485714e-01
R36533 n0_6054_19857 n0_6146_19857 5.257143e-01
R36534 n0_6146_19857 n0_8116_19857 1.125714e+01
R36535 n0_8116_19857 n0_8208_19857 5.257143e-01
R36536 n0_8208_19857 n0_8304_19857 5.485714e-01
R36537 n0_8304_19857 n0_8396_19857 5.257143e-01
R36538 n0_8396_19857 n0_10366_19857 1.125714e+01
R36539 n0_10366_19857 n0_10458_19857 5.257143e-01
R36540 n0_10458_19857 n0_10554_19857 5.485714e-01
R36541 n0_10554_19857 n0_10646_19857 5.257143e-01
R36542 n0_10646_19857 n0_12616_19857 1.125714e+01
R36543 n0_12616_19857 n0_12708_19857 5.257143e-01
R36544 n0_12708_19857 n0_12804_19857 5.485714e-01
R36545 n0_12804_19857 n0_12896_19857 5.257143e-01
R36546 n0_12896_19857 n0_14866_19857 1.125714e+01
R36547 n0_14866_19857 n0_14958_19857 5.257143e-01
R36548 n0_14958_19857 n0_15054_19857 5.485714e-01
R36549 n0_15054_19857 n0_15146_19857 5.257143e-01
R36550 n0_15146_19857 n0_17116_19857 1.125714e+01
R36551 n0_17116_19857 n0_17208_19857 5.257143e-01
R36552 n0_17208_19857 n0_17304_19857 5.485714e-01
R36553 n0_17304_19857 n0_17396_19857 5.257143e-01
R36554 n0_17396_19857 n0_19366_19857 1.125714e+01
R36555 n0_19366_19857 n0_19458_19857 5.257143e-01
R36556 n0_19458_19857 n0_19554_19857 5.485714e-01
R36557 n0_19554_19857 n0_19646_19857 5.257143e-01
R36558 n0_19646_19857 n0_20491_19857 4.828571e+00
R36559 n0_20491_19857 n0_20679_19857 1.074286e+00
R36560 n0_241_19890 n0_429_19890 1.074286e+00
R36561 n0_429_19890 n0_1366_19890 5.354286e+00
R36562 n0_1366_19890 n0_1458_19890 5.257143e-01
R36563 n0_1458_19890 n0_1554_19890 5.485714e-01
R36564 n0_1554_19890 n0_1646_19890 5.257143e-01
R36565 n0_1646_19890 n0_3616_19890 1.125714e+01
R36566 n0_3616_19890 n0_3708_19890 5.257143e-01
R36567 n0_3708_19890 n0_3804_19890 5.485714e-01
R36568 n0_3804_19890 n0_3896_19890 5.257143e-01
R36569 n0_3896_19890 n0_5866_19890 1.125714e+01
R36570 n0_5866_19890 n0_5958_19890 5.257143e-01
R36571 n0_5958_19890 n0_6054_19890 5.485714e-01
R36572 n0_6054_19890 n0_6146_19890 5.257143e-01
R36573 n0_6146_19890 n0_8116_19890 1.125714e+01
R36574 n0_8116_19890 n0_8208_19890 5.257143e-01
R36575 n0_8208_19890 n0_8304_19890 5.485714e-01
R36576 n0_8304_19890 n0_8396_19890 5.257143e-01
R36577 n0_8396_19890 n0_10366_19890 1.125714e+01
R36578 n0_10366_19890 n0_10458_19890 5.257143e-01
R36579 n0_10458_19890 n0_10554_19890 5.485714e-01
R36580 n0_10554_19890 n0_10646_19890 5.257143e-01
R36581 n0_10646_19890 n0_12616_19890 1.125714e+01
R36582 n0_12616_19890 n0_12708_19890 5.257143e-01
R36583 n0_12708_19890 n0_12804_19890 5.485714e-01
R36584 n0_12804_19890 n0_12896_19890 5.257143e-01
R36585 n0_12896_19890 n0_14866_19890 1.125714e+01
R36586 n0_14866_19890 n0_14958_19890 5.257143e-01
R36587 n0_14958_19890 n0_15054_19890 5.485714e-01
R36588 n0_15054_19890 n0_15146_19890 5.257143e-01
R36589 n0_15146_19890 n0_17116_19890 1.125714e+01
R36590 n0_17116_19890 n0_17208_19890 5.257143e-01
R36591 n0_17208_19890 n0_17304_19890 5.485714e-01
R36592 n0_17304_19890 n0_17396_19890 5.257143e-01
R36593 n0_17396_19890 n0_19366_19890 1.125714e+01
R36594 n0_19366_19890 n0_19458_19890 5.257143e-01
R36595 n0_19458_19890 n0_19554_19890 5.485714e-01
R36596 n0_19554_19890 n0_19646_19890 5.257143e-01
R36597 n0_19646_19890 n0_20491_19890 4.828571e+00
R36598 n0_20491_19890 n0_20679_19890 1.074286e+00
R36599 n0_241_20073 n0_429_20073 1.074286e+00
R36600 n0_429_20073 n0_1366_20073 5.354286e+00
R36601 n0_1366_20073 n0_1458_20073 5.257143e-01
R36602 n0_1458_20073 n0_1554_20073 5.485714e-01
R36603 n0_1554_20073 n0_1646_20073 5.257143e-01
R36604 n0_1646_20073 n0_3616_20073 1.125714e+01
R36605 n0_3616_20073 n0_3708_20073 5.257143e-01
R36606 n0_3708_20073 n0_3804_20073 5.485714e-01
R36607 n0_3804_20073 n0_3896_20073 5.257143e-01
R36608 n0_3896_20073 n0_5866_20073 1.125714e+01
R36609 n0_5866_20073 n0_5958_20073 5.257143e-01
R36610 n0_5958_20073 n0_6054_20073 5.485714e-01
R36611 n0_6054_20073 n0_6146_20073 5.257143e-01
R36612 n0_6146_20073 n0_8116_20073 1.125714e+01
R36613 n0_8116_20073 n0_8208_20073 5.257143e-01
R36614 n0_8208_20073 n0_8304_20073 5.485714e-01
R36615 n0_8304_20073 n0_8396_20073 5.257143e-01
R36616 n0_8396_20073 n0_10366_20073 1.125714e+01
R36617 n0_10366_20073 n0_10458_20073 5.257143e-01
R36618 n0_10458_20073 n0_10554_20073 5.485714e-01
R36619 n0_10554_20073 n0_10646_20073 5.257143e-01
R36620 n0_10646_20073 n0_12616_20073 1.125714e+01
R36621 n0_12616_20073 n0_12708_20073 5.257143e-01
R36622 n0_12708_20073 n0_12804_20073 5.485714e-01
R36623 n0_12804_20073 n0_12896_20073 5.257143e-01
R36624 n0_12896_20073 n0_14866_20073 1.125714e+01
R36625 n0_14866_20073 n0_14958_20073 5.257143e-01
R36626 n0_14958_20073 n0_15054_20073 5.485714e-01
R36627 n0_15054_20073 n0_15146_20073 5.257143e-01
R36628 n0_15146_20073 n0_17116_20073 1.125714e+01
R36629 n0_17116_20073 n0_17208_20073 5.257143e-01
R36630 n0_17208_20073 n0_17304_20073 5.485714e-01
R36631 n0_17304_20073 n0_17396_20073 5.257143e-01
R36632 n0_17396_20073 n0_19366_20073 1.125714e+01
R36633 n0_19366_20073 n0_19458_20073 5.257143e-01
R36634 n0_19458_20073 n0_19554_20073 5.485714e-01
R36635 n0_19554_20073 n0_19646_20073 5.257143e-01
R36636 n0_19646_20073 n0_20491_20073 4.828571e+00
R36637 n0_20491_20073 n0_20679_20073 1.074286e+00
R36638 n0_241_20106 n0_429_20106 1.074286e+00
R36639 n0_429_20106 n0_1366_20106 5.354286e+00
R36640 n0_1366_20106 n0_1458_20106 5.257143e-01
R36641 n0_1458_20106 n0_1554_20106 5.485714e-01
R36642 n0_1554_20106 n0_1646_20106 5.257143e-01
R36643 n0_1646_20106 n0_3616_20106 1.125714e+01
R36644 n0_3616_20106 n0_3708_20106 5.257143e-01
R36645 n0_3708_20106 n0_3804_20106 5.485714e-01
R36646 n0_3804_20106 n0_3896_20106 5.257143e-01
R36647 n0_3896_20106 n0_5866_20106 1.125714e+01
R36648 n0_5866_20106 n0_5958_20106 5.257143e-01
R36649 n0_5958_20106 n0_6054_20106 5.485714e-01
R36650 n0_6054_20106 n0_6146_20106 5.257143e-01
R36651 n0_6146_20106 n0_8116_20106 1.125714e+01
R36652 n0_8116_20106 n0_8208_20106 5.257143e-01
R36653 n0_8208_20106 n0_8304_20106 5.485714e-01
R36654 n0_8304_20106 n0_8396_20106 5.257143e-01
R36655 n0_8396_20106 n0_10366_20106 1.125714e+01
R36656 n0_10366_20106 n0_10458_20106 5.257143e-01
R36657 n0_10458_20106 n0_10554_20106 5.485714e-01
R36658 n0_10554_20106 n0_10646_20106 5.257143e-01
R36659 n0_10646_20106 n0_12616_20106 1.125714e+01
R36660 n0_12616_20106 n0_12708_20106 5.257143e-01
R36661 n0_12708_20106 n0_12804_20106 5.485714e-01
R36662 n0_12804_20106 n0_12896_20106 5.257143e-01
R36663 n0_12896_20106 n0_14866_20106 1.125714e+01
R36664 n0_14866_20106 n0_14958_20106 5.257143e-01
R36665 n0_14958_20106 n0_15054_20106 5.485714e-01
R36666 n0_15054_20106 n0_15146_20106 5.257143e-01
R36667 n0_15146_20106 n0_17116_20106 1.125714e+01
R36668 n0_17116_20106 n0_17208_20106 5.257143e-01
R36669 n0_17208_20106 n0_17304_20106 5.485714e-01
R36670 n0_17304_20106 n0_17396_20106 5.257143e-01
R36671 n0_17396_20106 n0_19366_20106 1.125714e+01
R36672 n0_19366_20106 n0_19458_20106 5.257143e-01
R36673 n0_19458_20106 n0_19554_20106 5.485714e-01
R36674 n0_19554_20106 n0_19646_20106 5.257143e-01
R36675 n0_19646_20106 n0_20491_20106 4.828571e+00
R36676 n0_20491_20106 n0_20679_20106 1.074286e+00
R36677 n0_241_20289 n0_429_20289 1.074286e+00
R36678 n0_429_20289 n0_1366_20289 5.354286e+00
R36679 n0_1366_20289 n0_1458_20289 5.257143e-01
R36680 n0_1458_20289 n0_1554_20289 5.485714e-01
R36681 n0_1554_20289 n0_1646_20289 5.257143e-01
R36682 n0_1646_20289 n0_3616_20289 1.125714e+01
R36683 n0_3616_20289 n0_3708_20289 5.257143e-01
R36684 n0_3708_20289 n0_3804_20289 5.485714e-01
R36685 n0_3804_20289 n0_3896_20289 5.257143e-01
R36686 n0_3896_20289 n0_5866_20289 1.125714e+01
R36687 n0_5866_20289 n0_5958_20289 5.257143e-01
R36688 n0_5958_20289 n0_6054_20289 5.485714e-01
R36689 n0_6054_20289 n0_6146_20289 5.257143e-01
R36690 n0_6146_20289 n0_8116_20289 1.125714e+01
R36691 n0_8116_20289 n0_8208_20289 5.257143e-01
R36692 n0_8208_20289 n0_8304_20289 5.485714e-01
R36693 n0_8304_20289 n0_8396_20289 5.257143e-01
R36694 n0_8396_20289 n0_10366_20289 1.125714e+01
R36695 n0_10366_20289 n0_10458_20289 5.257143e-01
R36696 n0_10458_20289 n0_10554_20289 5.485714e-01
R36697 n0_10554_20289 n0_10646_20289 5.257143e-01
R36698 n0_10646_20289 n0_12616_20289 1.125714e+01
R36699 n0_12616_20289 n0_12708_20289 5.257143e-01
R36700 n0_12708_20289 n0_12804_20289 5.485714e-01
R36701 n0_12804_20289 n0_12896_20289 5.257143e-01
R36702 n0_12896_20289 n0_14866_20289 1.125714e+01
R36703 n0_14866_20289 n0_14958_20289 5.257143e-01
R36704 n0_14958_20289 n0_15054_20289 5.485714e-01
R36705 n0_15054_20289 n0_15146_20289 5.257143e-01
R36706 n0_15146_20289 n0_17116_20289 1.125714e+01
R36707 n0_17116_20289 n0_17208_20289 5.257143e-01
R36708 n0_17208_20289 n0_17304_20289 5.485714e-01
R36709 n0_17304_20289 n0_17396_20289 5.257143e-01
R36710 n0_17396_20289 n0_19366_20289 1.125714e+01
R36711 n0_19366_20289 n0_19458_20289 5.257143e-01
R36712 n0_19458_20289 n0_19554_20289 5.485714e-01
R36713 n0_19554_20289 n0_19646_20289 5.257143e-01
R36714 n0_19646_20289 n0_20491_20289 4.828571e+00
R36715 n0_20491_20289 n0_20679_20289 1.074286e+00
R36716 n0_241_20322 n0_429_20322 1.074286e+00
R36717 n0_429_20322 n0_1366_20322 5.354286e+00
R36718 n0_1366_20322 n0_1458_20322 5.257143e-01
R36719 n0_1458_20322 n0_1554_20322 5.485714e-01
R36720 n0_1554_20322 n0_1646_20322 5.257143e-01
R36721 n0_1646_20322 n0_3616_20322 1.125714e+01
R36722 n0_3616_20322 n0_3708_20322 5.257143e-01
R36723 n0_3708_20322 n0_3804_20322 5.485714e-01
R36724 n0_3804_20322 n0_3896_20322 5.257143e-01
R36725 n0_3896_20322 n0_5866_20322 1.125714e+01
R36726 n0_5866_20322 n0_5958_20322 5.257143e-01
R36727 n0_5958_20322 n0_6054_20322 5.485714e-01
R36728 n0_6054_20322 n0_6146_20322 5.257143e-01
R36729 n0_6146_20322 n0_8116_20322 1.125714e+01
R36730 n0_8116_20322 n0_8208_20322 5.257143e-01
R36731 n0_8208_20322 n0_8304_20322 5.485714e-01
R36732 n0_8304_20322 n0_8396_20322 5.257143e-01
R36733 n0_8396_20322 n0_10366_20322 1.125714e+01
R36734 n0_10366_20322 n0_10458_20322 5.257143e-01
R36735 n0_10458_20322 n0_10554_20322 5.485714e-01
R36736 n0_10554_20322 n0_10646_20322 5.257143e-01
R36737 n0_10646_20322 n0_12616_20322 1.125714e+01
R36738 n0_12616_20322 n0_12708_20322 5.257143e-01
R36739 n0_12708_20322 n0_12804_20322 5.485714e-01
R36740 n0_12804_20322 n0_12896_20322 5.257143e-01
R36741 n0_12896_20322 n0_14866_20322 1.125714e+01
R36742 n0_14866_20322 n0_14958_20322 5.257143e-01
R36743 n0_14958_20322 n0_15054_20322 5.485714e-01
R36744 n0_15054_20322 n0_15146_20322 5.257143e-01
R36745 n0_15146_20322 n0_17116_20322 1.125714e+01
R36746 n0_17116_20322 n0_17208_20322 5.257143e-01
R36747 n0_17208_20322 n0_17304_20322 5.485714e-01
R36748 n0_17304_20322 n0_17396_20322 5.257143e-01
R36749 n0_17396_20322 n0_19366_20322 1.125714e+01
R36750 n0_19366_20322 n0_19458_20322 5.257143e-01
R36751 n0_19458_20322 n0_19554_20322 5.485714e-01
R36752 n0_19554_20322 n0_19646_20322 5.257143e-01
R36753 n0_19646_20322 n0_20491_20322 4.828571e+00
R36754 n0_20491_20322 n0_20679_20322 1.074286e+00
R36755 n0_241_20505 n0_429_20505 1.074286e+00
R36756 n0_429_20505 n0_1366_20505 5.354286e+00
R36757 n0_1366_20505 n0_1458_20505 5.257143e-01
R36758 n0_1458_20505 n0_1554_20505 5.485714e-01
R36759 n0_1554_20505 n0_1646_20505 5.257143e-01
R36760 n0_1646_20505 n0_3616_20505 1.125714e+01
R36761 n0_3616_20505 n0_3708_20505 5.257143e-01
R36762 n0_3708_20505 n0_3804_20505 5.485714e-01
R36763 n0_3804_20505 n0_3896_20505 5.257143e-01
R36764 n0_3896_20505 n0_5866_20505 1.125714e+01
R36765 n0_5866_20505 n0_5958_20505 5.257143e-01
R36766 n0_5958_20505 n0_6054_20505 5.485714e-01
R36767 n0_6054_20505 n0_6146_20505 5.257143e-01
R36768 n0_6146_20505 n0_8116_20505 1.125714e+01
R36769 n0_8116_20505 n0_8208_20505 5.257143e-01
R36770 n0_8208_20505 n0_8304_20505 5.485714e-01
R36771 n0_8304_20505 n0_8396_20505 5.257143e-01
R36772 n0_8396_20505 n0_10366_20505 1.125714e+01
R36773 n0_10366_20505 n0_10458_20505 5.257143e-01
R36774 n0_10458_20505 n0_10554_20505 5.485714e-01
R36775 n0_10554_20505 n0_10646_20505 5.257143e-01
R36776 n0_10646_20505 n0_12616_20505 1.125714e+01
R36777 n0_12616_20505 n0_12708_20505 5.257143e-01
R36778 n0_12708_20505 n0_12804_20505 5.485714e-01
R36779 n0_12804_20505 n0_12896_20505 5.257143e-01
R36780 n0_12896_20505 n0_14866_20505 1.125714e+01
R36781 n0_14866_20505 n0_14958_20505 5.257143e-01
R36782 n0_14958_20505 n0_15054_20505 5.485714e-01
R36783 n0_15054_20505 n0_15146_20505 5.257143e-01
R36784 n0_15146_20505 n0_17116_20505 1.125714e+01
R36785 n0_17116_20505 n0_17208_20505 5.257143e-01
R36786 n0_17208_20505 n0_17304_20505 5.485714e-01
R36787 n0_17304_20505 n0_17396_20505 5.257143e-01
R36788 n0_17396_20505 n0_19366_20505 1.125714e+01
R36789 n0_19366_20505 n0_19458_20505 5.257143e-01
R36790 n0_19458_20505 n0_19554_20505 5.485714e-01
R36791 n0_19554_20505 n0_19646_20505 5.257143e-01
R36792 n0_19646_20505 n0_20491_20505 4.828571e+00
R36793 n0_20491_20505 n0_20679_20505 1.074286e+00
R36794 n0_241_20538 n0_429_20538 1.074286e+00
R36795 n0_429_20538 n0_1366_20538 5.354286e+00
R36796 n0_1366_20538 n0_1458_20538 5.257143e-01
R36797 n0_1458_20538 n0_1554_20538 5.485714e-01
R36798 n0_1554_20538 n0_1646_20538 5.257143e-01
R36799 n0_1646_20538 n0_3616_20538 1.125714e+01
R36800 n0_3616_20538 n0_3708_20538 5.257143e-01
R36801 n0_3708_20538 n0_3804_20538 5.485714e-01
R36802 n0_3804_20538 n0_3896_20538 5.257143e-01
R36803 n0_3896_20538 n0_5866_20538 1.125714e+01
R36804 n0_5866_20538 n0_5958_20538 5.257143e-01
R36805 n0_5958_20538 n0_6054_20538 5.485714e-01
R36806 n0_6054_20538 n0_6146_20538 5.257143e-01
R36807 n0_6146_20538 n0_8116_20538 1.125714e+01
R36808 n0_8116_20538 n0_8208_20538 5.257143e-01
R36809 n0_8208_20538 n0_8304_20538 5.485714e-01
R36810 n0_8304_20538 n0_8396_20538 5.257143e-01
R36811 n0_8396_20538 n0_10366_20538 1.125714e+01
R36812 n0_10366_20538 n0_10458_20538 5.257143e-01
R36813 n0_10458_20538 n0_10554_20538 5.485714e-01
R36814 n0_10554_20538 n0_10646_20538 5.257143e-01
R36815 n0_10646_20538 n0_12616_20538 1.125714e+01
R36816 n0_12616_20538 n0_12708_20538 5.257143e-01
R36817 n0_12708_20538 n0_12804_20538 5.485714e-01
R36818 n0_12804_20538 n0_12896_20538 5.257143e-01
R36819 n0_12896_20538 n0_14866_20538 1.125714e+01
R36820 n0_14866_20538 n0_14958_20538 5.257143e-01
R36821 n0_14958_20538 n0_15054_20538 5.485714e-01
R36822 n0_15054_20538 n0_15146_20538 5.257143e-01
R36823 n0_15146_20538 n0_17116_20538 1.125714e+01
R36824 n0_17116_20538 n0_17208_20538 5.257143e-01
R36825 n0_17208_20538 n0_17304_20538 5.485714e-01
R36826 n0_17304_20538 n0_17396_20538 5.257143e-01
R36827 n0_17396_20538 n0_19366_20538 1.125714e+01
R36828 n0_19366_20538 n0_19458_20538 5.257143e-01
R36829 n0_19458_20538 n0_19554_20538 5.485714e-01
R36830 n0_19554_20538 n0_19646_20538 5.257143e-01
R36831 n0_19646_20538 n0_20491_20538 4.828571e+00
R36832 n0_20491_20538 n0_20679_20538 1.074286e+00
R36833 n0_1458_20721 n0_1505_20721 2.685714e-01
R36834 n0_1505_20721 n0_1554_20721 2.800000e-01
R36835 n0_1554_20721 n0_3708_20721 1.230857e+01
R36836 n0_3708_20721 n0_3755_20721 2.685714e-01
R36837 n0_3755_20721 n0_3804_20721 2.800000e-01
R36838 n0_3804_20721 n0_5958_20721 1.230857e+01
R36839 n0_5958_20721 n0_6005_20721 2.685714e-01
R36840 n0_6005_20721 n0_6054_20721 2.800000e-01
R36841 n0_6054_20721 n0_8208_20721 1.230857e+01
R36842 n0_8208_20721 n0_8255_20721 2.685714e-01
R36843 n0_8255_20721 n0_8304_20721 2.800000e-01
R36844 n0_8304_20721 n0_10458_20721 1.230857e+01
R36845 n0_10458_20721 n0_10505_20721 2.685714e-01
R36846 n0_10505_20721 n0_10554_20721 2.800000e-01
R36847 n0_10554_20721 n0_12708_20721 1.230857e+01
R36848 n0_12708_20721 n0_12755_20721 2.685714e-01
R36849 n0_12755_20721 n0_12804_20721 2.800000e-01
R36850 n0_12804_20721 n0_14958_20721 1.230857e+01
R36851 n0_14958_20721 n0_15005_20721 2.685714e-01
R36852 n0_15005_20721 n0_15054_20721 2.800000e-01
R36853 n0_15054_20721 n0_17208_20721 1.230857e+01
R36854 n0_17208_20721 n0_17255_20721 2.685714e-01
R36855 n0_17255_20721 n0_17304_20721 2.800000e-01
R36856 n0_17304_20721 n0_19458_20721 1.230857e+01
R36857 n0_19458_20721 n0_19505_20721 2.685714e-01
R36858 n0_19505_20721 n0_19554_20721 2.800000e-01
R36859 n0_1366_20754 n0_1458_20754 5.257143e-01
R36860 n0_1458_20754 n0_1505_20754 2.685714e-01
R36861 n0_1505_20754 n0_1554_20754 2.800000e-01
R36862 n0_1554_20754 n0_1646_20754 5.257143e-01
R36863 n0_1646_20754 n0_3616_20754 1.125714e+01
R36864 n0_3616_20754 n0_3708_20754 5.257143e-01
R36865 n0_3708_20754 n0_3755_20754 2.685714e-01
R36866 n0_3755_20754 n0_3804_20754 2.800000e-01
R36867 n0_3804_20754 n0_3896_20754 5.257143e-01
R36868 n0_3896_20754 n0_5866_20754 1.125714e+01
R36869 n0_5866_20754 n0_5958_20754 5.257143e-01
R36870 n0_5958_20754 n0_6005_20754 2.685714e-01
R36871 n0_6005_20754 n0_6054_20754 2.800000e-01
R36872 n0_6054_20754 n0_6146_20754 5.257143e-01
R36873 n0_6146_20754 n0_8116_20754 1.125714e+01
R36874 n0_8116_20754 n0_8208_20754 5.257143e-01
R36875 n0_8208_20754 n0_8255_20754 2.685714e-01
R36876 n0_8255_20754 n0_8304_20754 2.800000e-01
R36877 n0_8304_20754 n0_8396_20754 5.257143e-01
R36878 n0_8396_20754 n0_10366_20754 1.125714e+01
R36879 n0_10366_20754 n0_10458_20754 5.257143e-01
R36880 n0_10458_20754 n0_10505_20754 2.685714e-01
R36881 n0_10505_20754 n0_10554_20754 2.800000e-01
R36882 n0_10554_20754 n0_10646_20754 5.257143e-01
R36883 n0_10646_20754 n0_12616_20754 1.125714e+01
R36884 n0_12616_20754 n0_12708_20754 5.257143e-01
R36885 n0_12708_20754 n0_12755_20754 2.685714e-01
R36886 n0_12755_20754 n0_12804_20754 2.800000e-01
R36887 n0_12804_20754 n0_12896_20754 5.257143e-01
R36888 n0_12896_20754 n0_14866_20754 1.125714e+01
R36889 n0_14866_20754 n0_14958_20754 5.257143e-01
R36890 n0_14958_20754 n0_15005_20754 2.685714e-01
R36891 n0_15005_20754 n0_15054_20754 2.800000e-01
R36892 n0_15054_20754 n0_15146_20754 5.257143e-01
R36893 n0_15146_20754 n0_17116_20754 1.125714e+01
R36894 n0_17116_20754 n0_17208_20754 5.257143e-01
R36895 n0_17208_20754 n0_17255_20754 2.685714e-01
R36896 n0_17255_20754 n0_17304_20754 2.800000e-01
R36897 n0_17304_20754 n0_17396_20754 5.257143e-01
R36898 n0_17396_20754 n0_19366_20754 1.125714e+01
R36899 n0_19366_20754 n0_19458_20754 5.257143e-01
R36900 n0_19458_20754 n0_19505_20754 2.685714e-01
R36901 n0_19505_20754 n0_19554_20754 2.800000e-01
R36902 n0_19554_20754 n0_19646_20754 5.257143e-01
R36903 n0_241_13663 n0_429_13663 1.342857e-01
R36904 n0_429_13663 n0_1366_13663 6.692857e-01
R36905 n0_1366_13663 n0_1554_13663 1.342857e-01
R36906 n0_241_4375 n0_429_4375 1.342857e-01
R36907 n0_429_4375 n0_1366_4375 6.692857e-01
R36908 n0_1366_4375 n0_1554_4375 1.342857e-01
R36909 n0_241_19040 n0_429_19040 4.700000e-01
R36910 n0_429_19040 n0_1366_19040 2.342500e+00
R36911 n0_1366_19040 n0_1554_19040 4.700000e-01
R36912 n0_241_19256 n0_429_19256 4.700000e-01
R36913 n0_429_19256 n0_1366_19256 2.342500e+00
R36914 n0_1366_19256 n0_1554_19256 4.700000e-01
R36915 n0_241_19472 n0_429_19472 4.700000e-01
R36916 n0_429_19472 n0_1366_19472 2.342500e+00
R36917 n0_1366_19472 n0_1554_19472 4.700000e-01
R36918 n0_241_17960 n0_429_17960 4.700000e-01
R36919 n0_429_17960 n0_1366_17960 2.342500e+00
R36920 n0_1366_17960 n0_1554_17960 4.700000e-01
R36921 n0_1554_17960 n0_2491_17960 2.342500e+00
R36922 n0_2491_17960 n0_2679_17960 4.700000e-01
R36923 n0_1366_201 n0_1458_201 5.257143e-01
R36924 n0_1458_201 n0_1554_201 5.485714e-01
R36925 n0_1554_201 n0_1646_201 5.257143e-01
R36926 n0_1646_201 n0_3616_201 1.125714e+01
R36927 n0_3616_201 n0_3708_201 5.257143e-01
R36928 n0_3708_201 n0_3804_201 5.485714e-01
R36929 n0_3804_201 n0_3896_201 5.257143e-01
R36930 n0_3896_201 n0_5866_201 1.125714e+01
R36931 n0_5866_201 n0_5958_201 5.257143e-01
R36932 n0_5958_201 n0_6054_201 5.485714e-01
R36933 n0_6054_201 n0_6146_201 5.257143e-01
R36934 n0_6146_201 n0_8116_201 1.125714e+01
R36935 n0_8116_201 n0_8208_201 5.257143e-01
R36936 n0_8208_201 n0_8304_201 5.485714e-01
R36937 n0_8304_201 n0_8396_201 5.257143e-01
R36938 n0_1366_234 n0_1458_234 5.257143e-01
R36939 n0_1458_234 n0_1554_234 5.485714e-01
R36940 n0_1554_234 n0_1646_234 5.257143e-01
R36941 n0_1646_234 n0_3616_234 1.125714e+01
R36942 n0_3616_234 n0_3708_234 5.257143e-01
R36943 n0_3708_234 n0_3804_234 5.485714e-01
R36944 n0_3804_234 n0_3896_234 5.257143e-01
R36945 n0_3896_234 n0_5866_234 1.125714e+01
R36946 n0_5866_234 n0_5958_234 5.257143e-01
R36947 n0_5958_234 n0_6054_234 5.485714e-01
R36948 n0_6054_234 n0_6146_234 5.257143e-01
R36949 n0_6146_234 n0_8116_234 1.125714e+01
R36950 n0_8116_234 n0_8208_234 5.257143e-01
R36951 n0_8208_234 n0_8304_234 5.485714e-01
R36952 n0_8304_234 n0_8396_234 5.257143e-01
R36953 n0_1366_20937 n0_1458_20937 5.257143e-01
R36954 n0_1458_20937 n0_1554_20937 5.485714e-01
R36955 n0_1554_20937 n0_1646_20937 5.257143e-01
R36956 n0_1646_20937 n0_3616_20937 1.125714e+01
R36957 n0_3616_20937 n0_3708_20937 5.257143e-01
R36958 n0_3708_20937 n0_3804_20937 5.485714e-01
R36959 n0_3804_20937 n0_3896_20937 5.257143e-01
R36960 n0_3896_20937 n0_5866_20937 1.125714e+01
R36961 n0_5866_20937 n0_5958_20937 5.257143e-01
R36962 n0_5958_20937 n0_6054_20937 5.485714e-01
R36963 n0_6054_20937 n0_6146_20937 5.257143e-01
R36964 n0_6146_20937 n0_8116_20937 1.125714e+01
R36965 n0_8116_20937 n0_8208_20937 5.257143e-01
R36966 n0_8208_20937 n0_8304_20937 5.485714e-01
R36967 n0_8304_20937 n0_8396_20937 5.257143e-01
R36968 n0_8396_20937 n0_10366_20937 1.125714e+01
R36969 n0_10366_20937 n0_10458_20937 5.257143e-01
R36970 n0_10458_20937 n0_10554_20937 5.485714e-01
R36971 n0_10554_20937 n0_10646_20937 5.257143e-01
R36972 n0_10646_20937 n0_12616_20937 1.125714e+01
R36973 n0_12616_20937 n0_12708_20937 5.257143e-01
R36974 n0_12708_20937 n0_12804_20937 5.485714e-01
R36975 n0_12804_20937 n0_12896_20937 5.257143e-01
R36976 n0_12896_20937 n0_14866_20937 1.125714e+01
R36977 n0_14866_20937 n0_14958_20937 5.257143e-01
R36978 n0_14958_20937 n0_15054_20937 5.485714e-01
R36979 n0_15054_20937 n0_15146_20937 5.257143e-01
R36980 n0_15146_20937 n0_17116_20937 1.125714e+01
R36981 n0_17116_20937 n0_17208_20937 5.257143e-01
R36982 n0_17208_20937 n0_17304_20937 5.485714e-01
R36983 n0_17304_20937 n0_17396_20937 5.257143e-01
R36984 n0_17396_20937 n0_19366_20937 1.125714e+01
R36985 n0_19366_20937 n0_19458_20937 5.257143e-01
R36986 n0_19458_20937 n0_19554_20937 5.485714e-01
R36987 n0_19554_20937 n0_19646_20937 5.257143e-01
R36988 n0_1366_20970 n0_1458_20970 5.257143e-01
R36989 n0_1458_20970 n0_1554_20970 5.485714e-01
R36990 n0_1554_20970 n0_1646_20970 5.257143e-01
R36991 n0_1646_20970 n0_3616_20970 1.125714e+01
R36992 n0_3616_20970 n0_3708_20970 5.257143e-01
R36993 n0_3708_20970 n0_3804_20970 5.485714e-01
R36994 n0_3804_20970 n0_3896_20970 5.257143e-01
R36995 n0_3896_20970 n0_5866_20970 1.125714e+01
R36996 n0_5866_20970 n0_5958_20970 5.257143e-01
R36997 n0_5958_20970 n0_6054_20970 5.485714e-01
R36998 n0_6054_20970 n0_6146_20970 5.257143e-01
R36999 n0_6146_20970 n0_8116_20970 1.125714e+01
R37000 n0_8116_20970 n0_8208_20970 5.257143e-01
R37001 n0_8208_20970 n0_8304_20970 5.485714e-01
R37002 n0_8304_20970 n0_8396_20970 5.257143e-01
R37003 n0_8396_20970 n0_10366_20970 1.125714e+01
R37004 n0_10366_20970 n0_10458_20970 5.257143e-01
R37005 n0_10458_20970 n0_10554_20970 5.485714e-01
R37006 n0_10554_20970 n0_10646_20970 5.257143e-01
R37007 n0_10646_20970 n0_12616_20970 1.125714e+01
R37008 n0_12616_20970 n0_12708_20970 5.257143e-01
R37009 n0_12708_20970 n0_12804_20970 5.485714e-01
R37010 n0_12804_20970 n0_12896_20970 5.257143e-01
R37011 n0_12896_20970 n0_14866_20970 1.125714e+01
R37012 n0_14866_20970 n0_14958_20970 5.257143e-01
R37013 n0_14958_20970 n0_15054_20970 5.485714e-01
R37014 n0_15054_20970 n0_15146_20970 5.257143e-01
R37015 n0_15146_20970 n0_17116_20970 1.125714e+01
R37016 n0_17116_20970 n0_17208_20970 5.257143e-01
R37017 n0_17208_20970 n0_17304_20970 5.485714e-01
R37018 n0_17304_20970 n0_17396_20970 5.257143e-01
R37019 n0_17396_20970 n0_19366_20970 1.125714e+01
R37020 n0_19366_20970 n0_19458_20970 5.257143e-01
R37021 n0_19458_20970 n0_19554_20970 5.485714e-01
R37022 n0_19554_20970 n0_19646_20970 5.257143e-01
R37023 n0_1366_1760 n0_1554_1760 4.700000e-01
R37024 n0_1366_3272 n0_1554_3272 4.700000e-01
R37025 n0_1554_3272 n0_2491_3272 2.342500e+00
R37026 n0_2491_3272 n0_2679_3272 4.700000e-01
R37027 n0_1366_11071 n0_1554_11071 1.342857e-01
R37028 n0_1554_11071 n0_2491_11071 6.692857e-01
R37029 n0_2491_11071 n0_2679_11071 1.342857e-01
R37030 n0_1366_13447 n0_1554_13447 1.342857e-01
R37031 n0_1554_13447 n0_2491_13447 6.692857e-01
R37032 n0_2491_13447 n0_2679_13447 1.342857e-01
R37033 n0_1366_14504 n0_1554_14504 4.700000e-01
R37034 n0_1554_14504 n0_2491_14504 2.342500e+00
R37035 n0_2491_14504 n0_2679_14504 4.700000e-01
R37036 n0_1366_16687 n0_1554_16687 1.342857e-01
R37037 n0_1554_16687 n0_2491_16687 6.692857e-01
R37038 n0_2491_16687 n0_2679_16687 1.342857e-01
R37039 n0_1366_4159 n0_1554_4159 1.342857e-01
R37040 n0_1554_4159 n0_2491_4159 6.692857e-01
R37041 n0_2491_4159 n0_2679_4159 1.342857e-01
R37042 n0_2679_4159 n0_3616_4159 6.692857e-01
R37043 n0_3616_4159 n0_3804_4159 1.342857e-01
R37044 n0_1366_8911 n0_1554_8911 1.342857e-01
R37045 n0_1554_8911 n0_2491_8911 6.692857e-01
R37046 n0_2491_8911 n0_2679_8911 1.342857e-01
R37047 n0_2679_8911 n0_3616_8911 6.692857e-01
R37048 n0_3616_8911 n0_3804_8911 1.342857e-01
R37049 n0_1366_16471 n0_1554_16471 1.342857e-01
R37050 n0_1554_16471 n0_2491_16471 6.692857e-01
R37051 n0_2491_16471 n0_2679_16471 1.342857e-01
R37052 n0_2679_16471 n0_3616_16471 6.692857e-01
R37053 n0_3616_16471 n0_3804_16471 1.342857e-01
R37054 n0_1366_3920 n0_1505_3920 3.475000e-01
R37055 n0_1505_3920 n0_1554_3920 1.225000e-01
R37056 n0_1554_3920 n0_2491_3920 2.342500e+00
R37057 n0_2491_3920 n0_2630_3920 3.475000e-01
R37058 n0_2630_3920 n0_2679_3920 1.225000e-01
R37059 n0_2679_3920 n0_3616_3920 2.342500e+00
R37060 n0_3616_3920 n0_3708_3920 2.300000e-01
R37061 n0_3708_3920 n0_3755_3920 1.175000e-01
R37062 n0_3755_3920 n0_3804_3920 1.225000e-01
R37063 n0_1366_3704 n0_1554_3704 4.700000e-01
R37064 n0_1554_3704 n0_2491_3704 2.342500e+00
R37065 n0_2491_3704 n0_2679_3704 4.700000e-01
R37066 n0_2679_3704 n0_3616_3704 2.342500e+00
R37067 n0_3616_3704 n0_3708_3704 2.300000e-01
R37068 n0_3708_3704 n0_3804_3704 2.400000e-01
R37069 n0_3804_3704 n0_3896_3704 2.300000e-01
R37070 n0_1366_4352 n0_1554_4352 4.700000e-01
R37071 n0_1554_4352 n0_2491_4352 2.342500e+00
R37072 n0_2491_4352 n0_2679_4352 4.700000e-01
R37073 n0_2679_4352 n0_3616_4352 2.342500e+00
R37074 n0_3616_4352 n0_3804_4352 4.700000e-01
R37075 n0_1366_16880 n0_1554_16880 4.700000e-01
R37076 n0_1554_16880 n0_2491_16880 2.342500e+00
R37077 n0_2491_16880 n0_2679_16880 4.700000e-01
R37078 n0_2679_16880 n0_3616_16880 2.342500e+00
R37079 n0_3616_16880 n0_3804_16880 4.700000e-01
R37080 n0_1366_15368 n0_1554_15368 4.700000e-01
R37081 n0_1554_15368 n0_2491_15368 2.342500e+00
R37082 n0_2491_15368 n0_2679_15368 4.700000e-01
R37083 n0_2679_15368 n0_3616_15368 2.342500e+00
R37084 n0_3616_15368 n0_3804_15368 4.700000e-01
R37085 n0_3804_15368 n0_4741_15368 2.342500e+00
R37086 n0_4741_15368 n0_4929_15368 4.700000e-01
R37087 n0_1366_17528 n0_1554_17528 4.700000e-01
R37088 n0_1554_17528 n0_2491_17528 2.342500e+00
R37089 n0_2491_17528 n0_2679_17528 4.700000e-01
R37090 n0_2679_17528 n0_3616_17528 2.342500e+00
R37091 n0_3616_17528 n0_3708_17528 2.300000e-01
R37092 n0_3708_17528 n0_3804_17528 2.400000e-01
R37093 n0_3804_17528 n0_3896_17528 2.300000e-01
R37094 n0_3896_17528 n0_5866_17528 4.925000e+00
R37095 n0_5866_17528 n0_5958_17528 2.300000e-01
R37096 n0_5958_17528 n0_6054_17528 2.400000e-01
R37097 n0_6054_17528 n0_6146_17528 2.300000e-01
R37098 n0_1366_5432 n0_1554_5432 4.700000e-01
R37099 n0_1554_5432 n0_2491_5432 2.342500e+00
R37100 n0_2491_5432 n0_2679_5432 4.700000e-01
R37101 n0_2679_5432 n0_3616_5432 2.342500e+00
R37102 n0_3616_5432 n0_3804_5432 4.700000e-01
R37103 n0_3804_5432 n0_4741_5432 2.342500e+00
R37104 n0_4741_5432 n0_4929_5432 4.700000e-01
R37105 n0_4929_5432 n0_5866_5432 2.342500e+00
R37106 n0_5866_5432 n0_5958_5432 2.300000e-01
R37107 n0_5958_5432 n0_6054_5432 2.400000e-01
R37108 n0_6054_5432 n0_6146_5432 2.300000e-01
R37109 n0_1366_6535 n0_1554_6535 1.342857e-01
R37110 n0_1554_6535 n0_2491_6535 6.692857e-01
R37111 n0_2491_6535 n0_2679_6535 1.342857e-01
R37112 n0_2679_6535 n0_3616_6535 6.692857e-01
R37113 n0_3616_6535 n0_3804_6535 1.342857e-01
R37114 n0_3804_6535 n0_4741_6535 6.692857e-01
R37115 n0_4741_6535 n0_4929_6535 1.342857e-01
R37116 n0_4929_6535 n0_5866_6535 6.692857e-01
R37117 n0_5866_6535 n0_6054_6535 1.342857e-01
R37118 n0_1366_8888 n0_1554_8888 4.700000e-01
R37119 n0_1554_8888 n0_2491_8888 2.342500e+00
R37120 n0_2491_8888 n0_2679_8888 4.700000e-01
R37121 n0_2679_8888 n0_3616_8888 2.342500e+00
R37122 n0_3616_8888 n0_3804_8888 4.700000e-01
R37123 n0_3804_8888 n0_4741_8888 2.342500e+00
R37124 n0_4741_8888 n0_4929_8888 4.700000e-01
R37125 n0_4929_8888 n0_5866_8888 2.342500e+00
R37126 n0_5866_8888 n0_6054_8888 4.700000e-01
R37127 n0_6054_8888 n0_6991_8888 2.342500e+00
R37128 n0_6991_8888 n0_7179_8888 4.700000e-01
R37129 n0_7179_8888 n0_8116_8888 2.342500e+00
R37130 n0_8116_8888 n0_8304_8888 4.700000e-01
R37131 n0_1366_9968 n0_1554_9968 4.700000e-01
R37132 n0_1554_9968 n0_2491_9968 2.342500e+00
R37133 n0_2491_9968 n0_2679_9968 4.700000e-01
R37134 n0_2679_9968 n0_3616_9968 2.342500e+00
R37135 n0_3616_9968 n0_3804_9968 4.700000e-01
R37136 n0_3804_9968 n0_4741_9968 2.342500e+00
R37137 n0_4741_9968 n0_4929_9968 4.700000e-01
R37138 n0_4929_9968 n0_5866_9968 2.342500e+00
R37139 n0_5866_9968 n0_6054_9968 4.700000e-01
R37140 n0_6054_9968 n0_6991_9968 2.342500e+00
R37141 n0_6991_9968 n0_7179_9968 4.700000e-01
R37142 n0_7179_9968 n0_8116_9968 2.342500e+00
R37143 n0_8116_9968 n0_8304_9968 4.700000e-01
R37144 n0_1366_11048 n0_1554_11048 4.700000e-01
R37145 n0_1554_11048 n0_2491_11048 2.342500e+00
R37146 n0_2491_11048 n0_2679_11048 4.700000e-01
R37147 n0_2679_11048 n0_3616_11048 2.342500e+00
R37148 n0_3616_11048 n0_3804_11048 4.700000e-01
R37149 n0_3804_11048 n0_4741_11048 2.342500e+00
R37150 n0_4741_11048 n0_4929_11048 4.700000e-01
R37151 n0_4929_11048 n0_5866_11048 2.342500e+00
R37152 n0_5866_11048 n0_6054_11048 4.700000e-01
R37153 n0_6054_11048 n0_6991_11048 2.342500e+00
R37154 n0_6991_11048 n0_7179_11048 4.700000e-01
R37155 n0_7179_11048 n0_8116_11048 2.342500e+00
R37156 n0_8116_11048 n0_8304_11048 4.700000e-01
R37157 n0_1366_12128 n0_1554_12128 4.700000e-01
R37158 n0_1554_12128 n0_2491_12128 2.342500e+00
R37159 n0_2491_12128 n0_2679_12128 4.700000e-01
R37160 n0_2679_12128 n0_3616_12128 2.342500e+00
R37161 n0_3616_12128 n0_3804_12128 4.700000e-01
R37162 n0_3804_12128 n0_4741_12128 2.342500e+00
R37163 n0_4741_12128 n0_4929_12128 4.700000e-01
R37164 n0_4929_12128 n0_5866_12128 2.342500e+00
R37165 n0_5866_12128 n0_6054_12128 4.700000e-01
R37166 n0_6054_12128 n0_6991_12128 2.342500e+00
R37167 n0_6991_12128 n0_7179_12128 4.700000e-01
R37168 n0_7179_12128 n0_8116_12128 2.342500e+00
R37169 n0_8116_12128 n0_8304_12128 4.700000e-01
R37170 n0_1366_7808 n0_1554_7808 4.700000e-01
R37171 n0_1554_7808 n0_2491_7808 2.342500e+00
R37172 n0_2491_7808 n0_2679_7808 4.700000e-01
R37173 n0_2679_7808 n0_3616_7808 2.342500e+00
R37174 n0_3616_7808 n0_3804_7808 4.700000e-01
R37175 n0_3804_7808 n0_4741_7808 2.342500e+00
R37176 n0_4741_7808 n0_4929_7808 4.700000e-01
R37177 n0_4929_7808 n0_5866_7808 2.342500e+00
R37178 n0_5866_7808 n0_6054_7808 4.700000e-01
R37179 n0_6054_7808 n0_6991_7808 2.342500e+00
R37180 n0_6991_7808 n0_7179_7808 4.700000e-01
R37181 n0_7179_7808 n0_8116_7808 2.342500e+00
R37182 n0_8116_7808 n0_8208_7808 2.300000e-01
R37183 n0_8208_7808 n0_8304_7808 2.400000e-01
R37184 n0_8304_7808 n0_8396_7808 2.300000e-01
R37185 n0_2491_12151 n0_2679_12151 1.342857e-01
R37186 n0_2679_12151 n0_3616_12151 6.692857e-01
R37187 n0_3616_12151 n0_3804_12151 1.342857e-01
R37188 n0_2491_13640 n0_2679_13640 4.700000e-01
R37189 n0_2679_13640 n0_3616_13640 2.342500e+00
R37190 n0_3616_13640 n0_3804_13640 4.700000e-01
R37191 n0_2491_16664 n0_2679_16664 4.700000e-01
R37192 n0_2679_16664 n0_3616_16664 2.342500e+00
R37193 n0_3616_16664 n0_3804_16664 4.700000e-01
R37194 n0_2491_17551 n0_2679_17551 1.342857e-01
R37195 n0_2679_17551 n0_3616_17551 6.692857e-01
R37196 n0_3616_17551 n0_3708_17551 6.571429e-02
R37197 n0_3708_17551 n0_3804_17551 6.857143e-02
R37198 n0_3804_17551 n0_3896_17551 6.571429e-02
R37199 n0_2491_14100 n0_2679_14100 1.342857e-01
R37200 n0_2679_14100 n0_3616_14100 6.692857e-01
R37201 n0_3616_14100 n0_3804_14100 1.342857e-01
R37202 n0_3804_14100 n0_4741_14100 6.692857e-01
R37203 n0_4741_14100 n0_4929_14100 1.342857e-01
R37204 n0_2491_13879 n0_3616_13879 8.035714e-01
R37205 n0_3616_13879 n0_4741_13879 8.035714e-01
R37206 n0_4741_13879 n0_5866_13879 8.035714e-01
R37207 n0_2491_15584 n0_2679_15584 4.700000e-01
R37208 n0_2679_15584 n0_3616_15584 2.342500e+00
R37209 n0_3616_15584 n0_3804_15584 4.700000e-01
R37210 n0_3804_15584 n0_4741_15584 2.342500e+00
R37211 n0_4741_15584 n0_4929_15584 4.700000e-01
R37212 n0_4929_15584 n0_5866_15584 2.342500e+00
R37213 n0_5866_15584 n0_5958_15584 2.300000e-01
R37214 n0_5958_15584 n0_6054_15584 2.400000e-01
R37215 n0_6054_15584 n0_6146_15584 2.300000e-01
R37216 n0_2491_13424 n0_2679_13424 4.700000e-01
R37217 n0_2679_13424 n0_3616_13424 2.342500e+00
R37218 n0_3616_13424 n0_3804_13424 4.700000e-01
R37219 n0_3804_13424 n0_4741_13424 2.342500e+00
R37220 n0_4741_13424 n0_4929_13424 4.700000e-01
R37221 n0_4929_13424 n0_5866_13424 2.342500e+00
R37222 n0_5866_13424 n0_6054_13424 4.700000e-01
R37223 n0_6054_13424 n0_6991_13424 2.342500e+00
R37224 n0_6991_13424 n0_7179_13424 4.700000e-01
R37225 n0_7179_13424 n0_8116_13424 2.342500e+00
R37226 n0_8116_13424 n0_8208_13424 2.300000e-01
R37227 n0_8208_13424 n0_8304_13424 2.400000e-01
R37228 n0_8304_13424 n0_8396_13424 2.300000e-01
R37229 n0_3616_1652 n0_3708_1652 2.300000e-01
R37230 n0_3708_1652 n0_3755_1652 1.175000e-01
R37231 n0_3755_1652 n0_3804_1652 1.225000e-01
R37232 n0_3804_1652 n0_3896_1652 2.300000e-01
R37233 n0_3616_1976 n0_3708_1976 2.300000e-01
R37234 n0_3708_1976 n0_3804_1976 2.400000e-01
R37235 n0_3804_1976 n0_3896_1976 2.300000e-01
R37236 n0_3616_4136 n0_3804_4136 4.700000e-01
R37237 n0_3616_356 n0_3708_356 2.300000e-01
R37238 n0_3708_356 n0_3804_356 2.400000e-01
R37239 n0_3804_356 n0_3896_356 2.300000e-01
R37240 n0_3896_356 n0_5866_356 4.925000e+00
R37241 n0_5866_356 n0_5958_356 2.300000e-01
R37242 n0_5958_356 n0_6054_356 2.400000e-01
R37243 n0_6054_356 n0_6146_356 2.300000e-01
R37244 n0_3616_788 n0_3708_788 2.300000e-01
R37245 n0_3708_788 n0_3804_788 2.400000e-01
R37246 n0_3804_788 n0_3896_788 2.300000e-01
R37247 n0_3896_788 n0_5866_788 4.925000e+00
R37248 n0_5866_788 n0_5958_788 2.300000e-01
R37249 n0_5958_788 n0_6054_788 2.400000e-01
R37250 n0_6054_788 n0_6146_788 2.300000e-01
R37251 n0_3616_4375 n0_3804_4375 1.342857e-01
R37252 n0_3804_4375 n0_5866_4375 1.472857e+00
R37253 n0_5866_4375 n0_5958_4375 6.571429e-02
R37254 n0_5958_4375 n0_6054_4375 6.857143e-02
R37255 n0_6054_4375 n0_6146_4375 6.571429e-02
R37256 n0_3708_17335 n0_3755_17335 3.357143e-02
R37257 n0_3755_17335 n0_3804_17335 3.500000e-02
R37258 n0_4741_8911 n0_4929_8911 1.342857e-01
R37259 n0_4929_8911 n0_5866_8911 6.692857e-01
R37260 n0_5866_8911 n0_6054_8911 1.342857e-01
R37261 n0_4741_11071 n0_4929_11071 1.342857e-01
R37262 n0_4929_11071 n0_5866_11071 6.692857e-01
R37263 n0_5866_11071 n0_6054_11071 1.342857e-01
R37264 n0_4741_16016 n0_4929_16016 4.700000e-01
R37265 n0_4929_16016 n0_5866_16016 2.342500e+00
R37266 n0_5866_16016 n0_5958_16016 2.300000e-01
R37267 n0_5958_16016 n0_6054_16016 2.400000e-01
R37268 n0_6054_16016 n0_6146_16016 2.300000e-01
R37269 n0_5958_17335 n0_6005_17335 3.357143e-02
R37270 n0_6005_17335 n0_6054_17335 3.500000e-02
R37271 n0_5866_3056 n0_5958_3056 2.300000e-01
R37272 n0_5958_3056 n0_6054_3056 2.400000e-01
R37273 n0_6054_3056 n0_6146_3056 2.300000e-01
R37274 n0_5866_4352 n0_5958_4352 2.300000e-01
R37275 n0_5958_4352 n0_6054_4352 2.400000e-01
R37276 n0_6054_4352 n0_6146_4352 2.300000e-01
R37277 n0_5866_1760 n0_5958_1760 2.300000e-01
R37278 n0_5958_1760 n0_6054_1760 2.400000e-01
R37279 n0_6054_1760 n0_6146_1760 2.300000e-01
R37280 n0_5866_2408 n0_5958_2408 2.300000e-01
R37281 n0_5958_2408 n0_6054_2408 2.400000e-01
R37282 n0_6054_2408 n0_6146_2408 2.300000e-01
R37283 n0_5866_2840 n0_5958_2840 2.300000e-01
R37284 n0_5958_2840 n0_6054_2840 2.400000e-01
R37285 n0_6054_2840 n0_6146_2840 2.300000e-01
R37286 n0_5866_3488 n0_5958_3488 2.300000e-01
R37287 n0_5958_3488 n0_6054_3488 2.400000e-01
R37288 n0_6054_3488 n0_6146_3488 2.300000e-01
R37289 n0_5866_4136 n0_5958_4136 2.300000e-01
R37290 n0_5958_4136 n0_6054_4136 2.400000e-01
R37291 n0_6054_4136 n0_6146_4136 2.300000e-01
R37292 n0_5866_18824 n0_5958_18824 2.300000e-01
R37293 n0_5958_18824 n0_6054_18824 2.400000e-01
R37294 n0_6054_18824 n0_6146_18824 2.300000e-01
R37295 n0_5866_19472 n0_5958_19472 2.300000e-01
R37296 n0_5958_19472 n0_6054_19472 2.400000e-01
R37297 n0_6054_19472 n0_6146_19472 2.300000e-01
R37298 n0_5866_17096 n0_5958_17096 2.300000e-01
R37299 n0_5958_17096 n0_6054_17096 2.400000e-01
R37300 n0_6054_17096 n0_6146_17096 2.300000e-01
R37301 n0_5866_17312 n0_5958_17312 2.300000e-01
R37302 n0_5958_17312 n0_6005_17312 1.175000e-01
R37303 n0_6005_17312 n0_6054_17312 1.225000e-01
R37304 n0_6054_17312 n0_6146_17312 2.300000e-01
R37305 n0_5866_18392 n0_5958_18392 2.300000e-01
R37306 n0_5958_18392 n0_6005_18392 1.175000e-01
R37307 n0_6005_18392 n0_6054_18392 1.225000e-01
R37308 n0_6054_18392 n0_6146_18392 2.300000e-01
R37309 n0_5866_18608 n0_5958_18608 2.300000e-01
R37310 n0_5958_18608 n0_6054_18608 2.400000e-01
R37311 n0_6054_18608 n0_6146_18608 2.300000e-01
R37312 n0_5866_19040 n0_5958_19040 2.300000e-01
R37313 n0_5958_19040 n0_6054_19040 2.400000e-01
R37314 n0_6054_19040 n0_6146_19040 2.300000e-01
R37315 n0_5866_4568 n0_5958_4568 2.300000e-01
R37316 n0_5958_4568 n0_6054_4568 2.400000e-01
R37317 n0_6054_4568 n0_6146_4568 2.300000e-01
R37318 n0_5866_5216 n0_5958_5216 2.300000e-01
R37319 n0_5958_5216 n0_6054_5216 2.400000e-01
R37320 n0_6054_5216 n0_6146_5216 2.300000e-01
R37321 n0_5866_15800 n0_5958_15800 2.300000e-01
R37322 n0_5958_15800 n0_6054_15800 2.400000e-01
R37323 n0_6054_15800 n0_6146_15800 2.300000e-01
R37324 n0_5866_5455 n0_5958_5455 6.571429e-02
R37325 n0_5958_5455 n0_6054_5455 6.857143e-02
R37326 n0_6054_5455 n0_6146_5455 6.571429e-02
R37327 n0_6146_5455 n0_8116_5455 1.407143e+00
R37328 n0_8116_5455 n0_8208_5455 6.571429e-02
R37329 n0_8208_5455 n0_8304_5455 6.857143e-02
R37330 n0_8304_5455 n0_8396_5455 6.571429e-02
R37331 n0_5866_17119 n0_5958_17119 6.571429e-02
R37332 n0_5958_17119 n0_6054_17119 6.857143e-02
R37333 n0_6054_17119 n0_6146_17119 6.571429e-02
R37334 n0_6146_17119 n0_8116_17119 1.407143e+00
R37335 n0_8116_17119 n0_8208_17119 6.571429e-02
R37336 n0_8208_17119 n0_8304_17119 6.857143e-02
R37337 n0_8304_17119 n0_8396_17119 6.571429e-02
R37338 n0_8396_17119 n0_10366_17119 1.407143e+00
R37339 n0_10366_17119 n0_10458_17119 6.571429e-02
R37340 n0_10458_17119 n0_10554_17119 6.857143e-02
R37341 n0_10554_17119 n0_10646_17119 6.571429e-02
R37342 n0_8116_1760 n0_8208_1760 2.300000e-01
R37343 n0_8208_1760 n0_8304_1760 2.400000e-01
R37344 n0_8304_1760 n0_8396_1760 2.300000e-01
R37345 n0_8116_2863 n0_8208_2863 6.571429e-02
R37346 n0_8208_2863 n0_8304_2863 6.857143e-02
R37347 n0_8304_2863 n0_8396_2863 6.571429e-02
R37348 n0_8116_18421 n0_8208_18421 6.571429e-02
R37349 n0_8208_18421 n0_8255_18421 3.357143e-02
R37350 n0_8255_18421 n0_8304_18421 3.500000e-02
R37351 n0_8304_18421 n0_8396_18421 6.571429e-02
R37352 n0_8116_19279 n0_8208_19279 6.571429e-02
R37353 n0_8208_19279 n0_8304_19279 6.857143e-02
R37354 n0_8304_19279 n0_8396_19279 6.571429e-02
R37355 n0_8116_6535 n0_8208_6535 6.571429e-02
R37356 n0_8208_6535 n0_8304_6535 6.857143e-02
R37357 n0_8304_6535 n0_8396_6535 6.571429e-02
R37358 n0_8116_3488 n0_8208_3488 2.300000e-01
R37359 n0_8208_3488 n0_8304_3488 2.400000e-01
R37360 n0_8304_3488 n0_8396_3488 2.300000e-01
R37361 n0_8116_4568 n0_8208_4568 2.300000e-01
R37362 n0_8208_4568 n0_8304_4568 2.400000e-01
R37363 n0_8304_4568 n0_8396_4568 2.300000e-01
R37364 n0_8116_2408 n0_8208_2408 2.300000e-01
R37365 n0_8208_2408 n0_8304_2408 2.400000e-01
R37366 n0_8304_2408 n0_8396_2408 2.300000e-01
R37367 n0_8116_4136 n0_8208_4136 2.300000e-01
R37368 n0_8208_4136 n0_8304_4136 2.400000e-01
R37369 n0_8304_4136 n0_8396_4136 2.300000e-01
R37370 n0_8116_5216 n0_8208_5216 2.300000e-01
R37371 n0_8208_5216 n0_8304_5216 2.400000e-01
R37372 n0_8304_5216 n0_8396_5216 2.300000e-01
R37373 n0_8116_5432 n0_8208_5432 2.300000e-01
R37374 n0_8208_5432 n0_8304_5432 2.400000e-01
R37375 n0_8304_5432 n0_8396_5432 2.300000e-01
R37376 n0_8116_15584 n0_8208_15584 2.300000e-01
R37377 n0_8208_15584 n0_8304_15584 2.400000e-01
R37378 n0_8304_15584 n0_8396_15584 2.300000e-01
R37379 n0_8116_15800 n0_8208_15800 2.300000e-01
R37380 n0_8208_15800 n0_8304_15800 2.400000e-01
R37381 n0_8304_15800 n0_8396_15800 2.300000e-01
R37382 n0_8116_16016 n0_8208_16016 2.300000e-01
R37383 n0_8208_16016 n0_8304_16016 2.400000e-01
R37384 n0_8304_16016 n0_8396_16016 2.300000e-01
R37385 n0_8116_17096 n0_8208_17096 2.300000e-01
R37386 n0_8208_17096 n0_8304_17096 2.400000e-01
R37387 n0_8304_17096 n0_8396_17096 2.300000e-01
R37388 n0_8116_17312 n0_8208_17312 2.300000e-01
R37389 n0_8208_17312 n0_8255_17312 1.175000e-01
R37390 n0_8255_17312 n0_8304_17312 1.225000e-01
R37391 n0_8304_17312 n0_8396_17312 2.300000e-01
R37392 n0_8116_18608 n0_8208_18608 2.300000e-01
R37393 n0_8208_18608 n0_8304_18608 2.400000e-01
R37394 n0_8304_18608 n0_8396_18608 2.300000e-01
R37395 n0_8116_14396 n0_8208_14396 2.300000e-01
R37396 n0_8208_14396 n0_8304_14396 2.400000e-01
R37397 n0_8304_14396 n0_8396_14396 2.300000e-01
R37398 n0_8116_1783 n0_8208_1783 6.571429e-02
R37399 n0_8208_1783 n0_8304_1783 6.857143e-02
R37400 n0_8304_1783 n0_8396_1783 6.571429e-02
R37401 n0_8116_2840 n0_8208_2840 2.300000e-01
R37402 n0_8208_2840 n0_8304_2840 2.400000e-01
R37403 n0_8304_2840 n0_8396_2840 2.300000e-01
R37404 n0_8116_6512 n0_8208_6512 2.300000e-01
R37405 n0_8208_6512 n0_8304_6512 2.400000e-01
R37406 n0_8304_6512 n0_8396_6512 2.300000e-01
R37407 n0_8116_6944 n0_8208_6944 2.300000e-01
R37408 n0_8208_6944 n0_8304_6944 2.400000e-01
R37409 n0_8304_6944 n0_8396_6944 2.300000e-01
R37410 n0_8116_7160 n0_8208_7160 2.300000e-01
R37411 n0_8208_7160 n0_8255_7160 1.175000e-01
R37412 n0_8255_7160 n0_8304_7160 1.225000e-01
R37413 n0_8304_7160 n0_8396_7160 2.300000e-01
R37414 n0_8116_7376 n0_8208_7376 2.300000e-01
R37415 n0_8208_7376 n0_8304_7376 2.400000e-01
R37416 n0_8304_7376 n0_8396_7376 2.300000e-01
R37417 n0_8116_13640 n0_8208_13640 2.300000e-01
R37418 n0_8208_13640 n0_8304_13640 2.400000e-01
R37419 n0_8304_13640 n0_8396_13640 2.300000e-01
R37420 n0_8116_13856 n0_8208_13856 2.300000e-01
R37421 n0_8208_13856 n0_8304_13856 2.400000e-01
R37422 n0_8304_13856 n0_8396_13856 2.300000e-01
R37423 n0_8116_14072 n0_8208_14072 2.300000e-01
R37424 n0_8208_14072 n0_8304_14072 2.400000e-01
R37425 n0_8304_14072 n0_8396_14072 2.300000e-01
R37426 n0_8116_14504 n0_8208_14504 2.300000e-01
R37427 n0_8208_14504 n0_8304_14504 2.400000e-01
R37428 n0_8304_14504 n0_8396_14504 2.300000e-01
R37429 n0_8116_18392 n0_8208_18392 2.300000e-01
R37430 n0_8208_18392 n0_8255_18392 1.175000e-01
R37431 n0_8255_18392 n0_8304_18392 1.225000e-01
R37432 n0_8304_18392 n0_8396_18392 2.300000e-01
R37433 n0_8116_19256 n0_8208_19256 2.300000e-01
R37434 n0_8208_19256 n0_8304_19256 2.400000e-01
R37435 n0_8304_19256 n0_8396_19256 2.300000e-01
R37436 n0_8116_5239 n0_8208_5239 6.571429e-02
R37437 n0_8208_5239 n0_8304_5239 6.857143e-02
R37438 n0_8304_5239 n0_8396_5239 6.571429e-02
R37439 n0_8396_5239 n0_10366_5239 1.407143e+00
R37440 n0_10366_5239 n0_10458_5239 6.571429e-02
R37441 n0_10458_5239 n0_10554_5239 6.857143e-02
R37442 n0_10554_5239 n0_10646_5239 6.571429e-02
R37443 n0_10366_1760 n0_10458_1760 2.300000e-01
R37444 n0_10458_1760 n0_10554_1760 2.400000e-01
R37445 n0_10554_1760 n0_10646_1760 2.300000e-01
R37446 n0_10366_2408 n0_10458_2408 2.300000e-01
R37447 n0_10458_2408 n0_10554_2408 2.400000e-01
R37448 n0_10554_2408 n0_10646_2408 2.300000e-01
R37449 n0_10366_2840 n0_10458_2840 2.300000e-01
R37450 n0_10458_2840 n0_10554_2840 2.400000e-01
R37451 n0_10554_2840 n0_10646_2840 2.300000e-01
R37452 n0_10366_3488 n0_10458_3488 2.300000e-01
R37453 n0_10458_3488 n0_10554_3488 2.400000e-01
R37454 n0_10554_3488 n0_10646_3488 2.300000e-01
R37455 n0_10366_4136 n0_10458_4136 2.300000e-01
R37456 n0_10458_4136 n0_10554_4136 2.400000e-01
R37457 n0_10554_4136 n0_10646_4136 2.300000e-01
R37458 n0_10366_4568 n0_10458_4568 2.300000e-01
R37459 n0_10458_4568 n0_10554_4568 2.400000e-01
R37460 n0_10554_4568 n0_10646_4568 2.300000e-01
R37461 n0_10366_5432 n0_10458_5432 2.300000e-01
R37462 n0_10458_5432 n0_10554_5432 2.400000e-01
R37463 n0_10554_5432 n0_10646_5432 2.300000e-01
R37464 n0_10366_6512 n0_10458_6512 2.300000e-01
R37465 n0_10458_6512 n0_10554_6512 2.400000e-01
R37466 n0_10554_6512 n0_10646_6512 2.300000e-01
R37467 n0_10366_6944 n0_10458_6944 2.300000e-01
R37468 n0_10458_6944 n0_10554_6944 2.400000e-01
R37469 n0_10554_6944 n0_10646_6944 2.300000e-01
R37470 n0_10366_7160 n0_10458_7160 2.300000e-01
R37471 n0_10458_7160 n0_10505_7160 1.175000e-01
R37472 n0_10505_7160 n0_10554_7160 1.225000e-01
R37473 n0_10554_7160 n0_10646_7160 2.300000e-01
R37474 n0_10366_7376 n0_10458_7376 2.300000e-01
R37475 n0_10458_7376 n0_10554_7376 2.400000e-01
R37476 n0_10554_7376 n0_10646_7376 2.300000e-01
R37477 n0_10366_13879 n0_10458_13879 6.571429e-02
R37478 n0_10458_13879 n0_10554_13879 6.857143e-02
R37479 n0_10554_13879 n0_10646_13879 6.571429e-02
R37480 n0_10366_14072 n0_10458_14072 2.300000e-01
R37481 n0_10458_14072 n0_10554_14072 2.400000e-01
R37482 n0_10554_14072 n0_10646_14072 2.300000e-01
R37483 n0_10366_15823 n0_10458_15823 6.571429e-02
R37484 n0_10458_15823 n0_10554_15823 6.857143e-02
R37485 n0_10554_15823 n0_10646_15823 6.571429e-02
R37486 n0_10366_17096 n0_10458_17096 2.300000e-01
R37487 n0_10458_17096 n0_10554_17096 2.400000e-01
R37488 n0_10554_17096 n0_10646_17096 2.300000e-01
R37489 n0_10366_13640 n0_10458_13640 2.300000e-01
R37490 n0_10458_13640 n0_10554_13640 2.400000e-01
R37491 n0_10554_13640 n0_10646_13640 2.300000e-01
R37492 n0_10366_14504 n0_10458_14504 2.300000e-01
R37493 n0_10458_14504 n0_10554_14504 2.400000e-01
R37494 n0_10554_14504 n0_10646_14504 2.300000e-01
R37495 n0_10366_15584 n0_10458_15584 2.300000e-01
R37496 n0_10458_15584 n0_10554_15584 2.400000e-01
R37497 n0_10554_15584 n0_10646_15584 2.300000e-01
R37498 n0_10366_16016 n0_10458_16016 2.300000e-01
R37499 n0_10458_16016 n0_10554_16016 2.400000e-01
R37500 n0_10554_16016 n0_10646_16016 2.300000e-01
R37501 n0_10366_17312 n0_10458_17312 2.300000e-01
R37502 n0_10458_17312 n0_10505_17312 1.175000e-01
R37503 n0_10505_17312 n0_10554_17312 1.225000e-01
R37504 n0_10554_17312 n0_10646_17312 2.300000e-01
R37505 n0_10366_18392 n0_10458_18392 2.300000e-01
R37506 n0_10458_18392 n0_10505_18392 1.175000e-01
R37507 n0_10505_18392 n0_10554_18392 1.225000e-01
R37508 n0_10554_18392 n0_10646_18392 2.300000e-01
R37509 n0_10366_18608 n0_10458_18608 2.300000e-01
R37510 n0_10458_18608 n0_10554_18608 2.400000e-01
R37511 n0_10554_18608 n0_10646_18608 2.300000e-01
R37512 n0_10366_19256 n0_10458_19256 2.300000e-01
R37513 n0_10458_19256 n0_10554_19256 2.400000e-01
R37514 n0_10554_19256 n0_10646_19256 2.300000e-01
R37515 n0_10366_201 n0_10458_201 5.257143e-01
R37516 n0_10458_201 n0_10554_201 5.485714e-01
R37517 n0_10554_201 n0_10646_201 5.257143e-01
R37518 n0_10646_201 n0_12616_201 1.125714e+01
R37519 n0_12616_201 n0_12708_201 5.257143e-01
R37520 n0_12708_201 n0_12804_201 5.485714e-01
R37521 n0_12804_201 n0_12896_201 5.257143e-01
R37522 n0_12896_201 n0_14866_201 1.125714e+01
R37523 n0_14866_201 n0_14958_201 5.257143e-01
R37524 n0_14958_201 n0_15054_201 5.485714e-01
R37525 n0_15054_201 n0_15146_201 5.257143e-01
R37526 n0_15146_201 n0_17116_201 1.125714e+01
R37527 n0_17116_201 n0_17208_201 5.257143e-01
R37528 n0_17208_201 n0_17304_201 5.485714e-01
R37529 n0_17304_201 n0_17396_201 5.257143e-01
R37530 n0_17396_201 n0_19366_201 1.125714e+01
R37531 n0_19366_201 n0_19458_201 5.257143e-01
R37532 n0_19458_201 n0_19554_201 5.485714e-01
R37533 n0_19554_201 n0_19646_201 5.257143e-01
R37534 n0_10366_234 n0_10458_234 5.257143e-01
R37535 n0_10458_234 n0_10554_234 5.485714e-01
R37536 n0_10554_234 n0_10646_234 5.257143e-01
R37537 n0_10646_234 n0_12616_234 1.125714e+01
R37538 n0_12616_234 n0_12708_234 5.257143e-01
R37539 n0_12708_234 n0_12804_234 5.485714e-01
R37540 n0_12804_234 n0_12896_234 5.257143e-01
R37541 n0_12896_234 n0_14866_234 1.125714e+01
R37542 n0_14866_234 n0_14958_234 5.257143e-01
R37543 n0_14958_234 n0_15054_234 5.485714e-01
R37544 n0_15054_234 n0_15146_234 5.257143e-01
R37545 n0_15146_234 n0_17116_234 1.125714e+01
R37546 n0_17116_234 n0_17208_234 5.257143e-01
R37547 n0_17208_234 n0_17304_234 5.485714e-01
R37548 n0_17304_234 n0_17396_234 5.257143e-01
R37549 n0_17396_234 n0_19366_234 1.125714e+01
R37550 n0_19366_234 n0_19458_234 5.257143e-01
R37551 n0_19458_234 n0_19554_234 5.485714e-01
R37552 n0_19554_234 n0_19646_234 5.257143e-01
R37553 n0_10366_417 n0_10458_417 5.257143e-01
R37554 n0_10458_417 n0_10505_417 2.685714e-01
R37555 n0_10505_417 n0_10554_417 2.800000e-01
R37556 n0_10554_417 n0_10646_417 5.257143e-01
R37557 n0_10646_417 n0_12616_417 1.125714e+01
R37558 n0_12616_417 n0_12708_417 5.257143e-01
R37559 n0_12708_417 n0_12755_417 2.685714e-01
R37560 n0_12755_417 n0_12804_417 2.800000e-01
R37561 n0_12804_417 n0_12896_417 5.257143e-01
R37562 n0_12896_417 n0_14866_417 1.125714e+01
R37563 n0_14866_417 n0_14958_417 5.257143e-01
R37564 n0_14958_417 n0_15005_417 2.685714e-01
R37565 n0_15005_417 n0_15054_417 2.800000e-01
R37566 n0_15054_417 n0_15146_417 5.257143e-01
R37567 n0_15146_417 n0_17116_417 1.125714e+01
R37568 n0_17116_417 n0_17208_417 5.257143e-01
R37569 n0_17208_417 n0_17255_417 2.685714e-01
R37570 n0_17255_417 n0_17304_417 2.800000e-01
R37571 n0_17304_417 n0_17396_417 5.257143e-01
R37572 n0_17396_417 n0_19366_417 1.125714e+01
R37573 n0_19366_417 n0_19458_417 5.257143e-01
R37574 n0_19458_417 n0_19505_417 2.685714e-01
R37575 n0_19505_417 n0_19554_417 2.800000e-01
R37576 n0_19554_417 n0_19646_417 5.257143e-01
R37577 n0_10366_450 n0_10458_450 5.257143e-01
R37578 n0_10458_450 n0_10505_450 2.685714e-01
R37579 n0_10505_450 n0_10554_450 2.800000e-01
R37580 n0_10554_450 n0_10646_450 5.257143e-01
R37581 n0_10646_450 n0_12616_450 1.125714e+01
R37582 n0_12616_450 n0_12708_450 5.257143e-01
R37583 n0_12708_450 n0_12755_450 2.685714e-01
R37584 n0_12755_450 n0_12804_450 2.800000e-01
R37585 n0_12804_450 n0_12896_450 5.257143e-01
R37586 n0_12896_450 n0_14866_450 1.125714e+01
R37587 n0_14866_450 n0_14958_450 5.257143e-01
R37588 n0_14958_450 n0_15005_450 2.685714e-01
R37589 n0_15005_450 n0_15054_450 2.800000e-01
R37590 n0_15054_450 n0_15146_450 5.257143e-01
R37591 n0_15146_450 n0_17116_450 1.125714e+01
R37592 n0_17116_450 n0_17208_450 5.257143e-01
R37593 n0_17208_450 n0_17255_450 2.685714e-01
R37594 n0_17255_450 n0_17304_450 2.800000e-01
R37595 n0_17304_450 n0_17396_450 5.257143e-01
R37596 n0_17396_450 n0_19366_450 1.125714e+01
R37597 n0_19366_450 n0_19458_450 5.257143e-01
R37598 n0_19458_450 n0_19505_450 2.685714e-01
R37599 n0_19505_450 n0_19554_450 2.800000e-01
R37600 n0_19554_450 n0_19646_450 5.257143e-01
R37601 n0_10366_633 n0_10458_633 5.257143e-01
R37602 n0_10458_633 n0_10554_633 5.485714e-01
R37603 n0_10554_633 n0_10646_633 5.257143e-01
R37604 n0_10646_633 n0_12616_633 1.125714e+01
R37605 n0_12616_633 n0_12708_633 5.257143e-01
R37606 n0_12708_633 n0_12804_633 5.485714e-01
R37607 n0_12804_633 n0_12896_633 5.257143e-01
R37608 n0_12896_633 n0_14866_633 1.125714e+01
R37609 n0_14866_633 n0_14958_633 5.257143e-01
R37610 n0_14958_633 n0_15054_633 5.485714e-01
R37611 n0_15054_633 n0_15146_633 5.257143e-01
R37612 n0_15146_633 n0_17116_633 1.125714e+01
R37613 n0_17116_633 n0_17208_633 5.257143e-01
R37614 n0_17208_633 n0_17304_633 5.485714e-01
R37615 n0_17304_633 n0_17396_633 5.257143e-01
R37616 n0_17396_633 n0_19366_633 1.125714e+01
R37617 n0_19366_633 n0_19458_633 5.257143e-01
R37618 n0_19458_633 n0_19554_633 5.485714e-01
R37619 n0_19554_633 n0_19646_633 5.257143e-01
R37620 n0_19646_633 n0_20491_633 4.828571e+00
R37621 n0_20491_633 n0_20679_633 1.074286e+00
R37622 n0_10366_666 n0_10458_666 5.257143e-01
R37623 n0_10458_666 n0_10554_666 5.485714e-01
R37624 n0_10554_666 n0_10646_666 5.257143e-01
R37625 n0_10646_666 n0_12616_666 1.125714e+01
R37626 n0_12616_666 n0_12708_666 5.257143e-01
R37627 n0_12708_666 n0_12804_666 5.485714e-01
R37628 n0_12804_666 n0_12896_666 5.257143e-01
R37629 n0_12896_666 n0_14866_666 1.125714e+01
R37630 n0_14866_666 n0_14958_666 5.257143e-01
R37631 n0_14958_666 n0_15054_666 5.485714e-01
R37632 n0_15054_666 n0_15146_666 5.257143e-01
R37633 n0_15146_666 n0_17116_666 1.125714e+01
R37634 n0_17116_666 n0_17208_666 5.257143e-01
R37635 n0_17208_666 n0_17304_666 5.485714e-01
R37636 n0_17304_666 n0_17396_666 5.257143e-01
R37637 n0_17396_666 n0_19366_666 1.125714e+01
R37638 n0_19366_666 n0_19458_666 5.257143e-01
R37639 n0_19458_666 n0_19554_666 5.485714e-01
R37640 n0_19554_666 n0_19646_666 5.257143e-01
R37641 n0_19646_666 n0_20491_666 4.828571e+00
R37642 n0_20491_666 n0_20679_666 1.074286e+00
R37643 n0_10366_849 n0_10458_849 5.257143e-01
R37644 n0_10458_849 n0_10554_849 5.485714e-01
R37645 n0_10554_849 n0_10646_849 5.257143e-01
R37646 n0_10646_849 n0_12616_849 1.125714e+01
R37647 n0_12616_849 n0_12708_849 5.257143e-01
R37648 n0_12708_849 n0_12804_849 5.485714e-01
R37649 n0_12804_849 n0_12896_849 5.257143e-01
R37650 n0_12896_849 n0_14866_849 1.125714e+01
R37651 n0_14866_849 n0_14958_849 5.257143e-01
R37652 n0_14958_849 n0_15054_849 5.485714e-01
R37653 n0_15054_849 n0_15146_849 5.257143e-01
R37654 n0_15146_849 n0_17116_849 1.125714e+01
R37655 n0_17116_849 n0_17208_849 5.257143e-01
R37656 n0_17208_849 n0_17304_849 5.485714e-01
R37657 n0_17304_849 n0_17396_849 5.257143e-01
R37658 n0_17396_849 n0_19366_849 1.125714e+01
R37659 n0_19366_849 n0_19458_849 5.257143e-01
R37660 n0_19458_849 n0_19554_849 5.485714e-01
R37661 n0_19554_849 n0_19646_849 5.257143e-01
R37662 n0_19646_849 n0_20491_849 4.828571e+00
R37663 n0_20491_849 n0_20679_849 1.074286e+00
R37664 n0_10366_882 n0_10458_882 5.257143e-01
R37665 n0_10458_882 n0_10554_882 5.485714e-01
R37666 n0_10554_882 n0_10646_882 5.257143e-01
R37667 n0_10646_882 n0_12616_882 1.125714e+01
R37668 n0_12616_882 n0_12708_882 5.257143e-01
R37669 n0_12708_882 n0_12804_882 5.485714e-01
R37670 n0_12804_882 n0_12896_882 5.257143e-01
R37671 n0_12896_882 n0_14866_882 1.125714e+01
R37672 n0_14866_882 n0_14958_882 5.257143e-01
R37673 n0_14958_882 n0_15054_882 5.485714e-01
R37674 n0_15054_882 n0_15146_882 5.257143e-01
R37675 n0_15146_882 n0_17116_882 1.125714e+01
R37676 n0_17116_882 n0_17208_882 5.257143e-01
R37677 n0_17208_882 n0_17304_882 5.485714e-01
R37678 n0_17304_882 n0_17396_882 5.257143e-01
R37679 n0_17396_882 n0_19366_882 1.125714e+01
R37680 n0_19366_882 n0_19458_882 5.257143e-01
R37681 n0_19458_882 n0_19554_882 5.485714e-01
R37682 n0_19554_882 n0_19646_882 5.257143e-01
R37683 n0_19646_882 n0_20491_882 4.828571e+00
R37684 n0_20491_882 n0_20679_882 1.074286e+00
R37685 n0_10366_1065 n0_10458_1065 5.257143e-01
R37686 n0_10458_1065 n0_10554_1065 5.485714e-01
R37687 n0_10554_1065 n0_10646_1065 5.257143e-01
R37688 n0_10646_1065 n0_12616_1065 1.125714e+01
R37689 n0_12616_1065 n0_12708_1065 5.257143e-01
R37690 n0_12708_1065 n0_12804_1065 5.485714e-01
R37691 n0_12804_1065 n0_12896_1065 5.257143e-01
R37692 n0_12896_1065 n0_14866_1065 1.125714e+01
R37693 n0_14866_1065 n0_14958_1065 5.257143e-01
R37694 n0_14958_1065 n0_15054_1065 5.485714e-01
R37695 n0_15054_1065 n0_15146_1065 5.257143e-01
R37696 n0_15146_1065 n0_17116_1065 1.125714e+01
R37697 n0_17116_1065 n0_17208_1065 5.257143e-01
R37698 n0_17208_1065 n0_17304_1065 5.485714e-01
R37699 n0_17304_1065 n0_17396_1065 5.257143e-01
R37700 n0_17396_1065 n0_19366_1065 1.125714e+01
R37701 n0_19366_1065 n0_19458_1065 5.257143e-01
R37702 n0_19458_1065 n0_19554_1065 5.485714e-01
R37703 n0_19554_1065 n0_19646_1065 5.257143e-01
R37704 n0_19646_1065 n0_20491_1065 4.828571e+00
R37705 n0_20491_1065 n0_20679_1065 1.074286e+00
R37706 n0_10366_1783 n0_10458_1783 6.571429e-02
R37707 n0_10458_1783 n0_10554_1783 6.857143e-02
R37708 n0_10554_1783 n0_10646_1783 6.571429e-02
R37709 n0_10366_2647 n0_10458_2647 6.571429e-02
R37710 n0_10458_2647 n0_10505_2647 3.357143e-02
R37711 n0_10505_2647 n0_10554_2647 3.500000e-02
R37712 n0_10554_2647 n0_10646_2647 6.571429e-02
R37713 n0_10366_2863 n0_10458_2863 6.571429e-02
R37714 n0_10458_2863 n0_10554_2863 6.857143e-02
R37715 n0_10554_2863 n0_10646_2863 6.571429e-02
R37716 n0_10366_3511 n0_10458_3511 6.571429e-02
R37717 n0_10458_3511 n0_10554_3511 6.857143e-02
R37718 n0_10554_3511 n0_10646_3511 6.571429e-02
R37719 n0_10366_4159 n0_10458_4159 6.571429e-02
R37720 n0_10458_4159 n0_10554_4159 6.857143e-02
R37721 n0_10554_4159 n0_10646_4159 6.571429e-02
R37722 n0_10366_4591 n0_10458_4591 6.571429e-02
R37723 n0_10458_4591 n0_10554_4591 6.857143e-02
R37724 n0_10554_4591 n0_10646_4591 6.571429e-02
R37725 n0_10366_5455 n0_10458_5455 6.571429e-02
R37726 n0_10458_5455 n0_10554_5455 6.857143e-02
R37727 n0_10554_5455 n0_10646_5455 6.571429e-02
R37728 n0_10366_6535 n0_10458_6535 6.571429e-02
R37729 n0_10458_6535 n0_10554_6535 6.857143e-02
R37730 n0_10554_6535 n0_10646_6535 6.571429e-02
R37731 n0_10366_6967 n0_10458_6967 6.571429e-02
R37732 n0_10458_6967 n0_10554_6967 6.857143e-02
R37733 n0_10554_6967 n0_10646_6967 6.571429e-02
R37734 n0_10366_7178 n0_10458_7178 6.571429e-02
R37735 n0_10458_7178 n0_10505_7178 3.357143e-02
R37736 n0_10505_7178 n0_10554_7178 3.500000e-02
R37737 n0_10554_7178 n0_10646_7178 6.571429e-02
R37738 n0_10366_7399 n0_10458_7399 6.571429e-02
R37739 n0_10458_7399 n0_10554_7399 6.857143e-02
R37740 n0_10554_7399 n0_10646_7399 6.571429e-02
R37741 n0_10366_13856 n0_10458_13856 2.300000e-01
R37742 n0_10458_13856 n0_10554_13856 2.400000e-01
R37743 n0_10554_13856 n0_10646_13856 2.300000e-01
R37744 n0_10366_14079 n0_10458_14079 1.187097e-01
R37745 n0_10458_14079 n0_10554_14079 1.238710e-01
R37746 n0_10554_14079 n0_10646_14079 1.187097e-01
R37747 n0_10366_15800 n0_10458_15800 2.300000e-01
R37748 n0_10458_15800 n0_10554_15800 2.400000e-01
R37749 n0_10554_15800 n0_10646_15800 2.300000e-01
R37750 n0_10366_17103 n0_10458_17103 1.187097e-01
R37751 n0_10458_17103 n0_10554_17103 1.238710e-01
R37752 n0_10554_17103 n0_10646_17103 1.187097e-01
R37753 n0_10366_6751 n0_10458_6751 6.571429e-02
R37754 n0_10458_6751 n0_10554_6751 6.857143e-02
R37755 n0_10554_6751 n0_10646_6751 6.571429e-02
R37756 n0_10646_6751 n0_12616_6751 1.407143e+00
R37757 n0_12616_6751 n0_12708_6751 6.571429e-02
R37758 n0_12708_6751 n0_12804_6751 6.857143e-02
R37759 n0_12804_6751 n0_12896_6751 6.571429e-02
R37760 n0_10366_13663 n0_10458_13663 6.571429e-02
R37761 n0_10458_13663 n0_10554_13663 6.857143e-02
R37762 n0_10554_13663 n0_10646_13663 6.571429e-02
R37763 n0_10646_13663 n0_12616_13663 1.407143e+00
R37764 n0_12616_13663 n0_12708_13663 6.571429e-02
R37765 n0_12708_13663 n0_12804_13663 6.857143e-02
R37766 n0_12804_13663 n0_12896_13663 6.571429e-02
R37767 n0_12616_6967 n0_12708_6967 6.571429e-02
R37768 n0_12708_6967 n0_12804_6967 6.857143e-02
R37769 n0_12804_6967 n0_12896_6967 6.571429e-02
R37770 n0_12616_5239 n0_12708_5239 6.571429e-02
R37771 n0_12708_5239 n0_12804_5239 6.857143e-02
R37772 n0_12804_5239 n0_12896_5239 6.571429e-02
R37773 n0_12616_7178 n0_12708_7178 6.571429e-02
R37774 n0_12708_7178 n0_12755_7178 3.357143e-02
R37775 n0_12755_7178 n0_12804_7178 3.500000e-02
R37776 n0_12804_7178 n0_12896_7178 6.571429e-02
R37777 n0_12616_7399 n0_12708_7399 6.571429e-02
R37778 n0_12708_7399 n0_12804_7399 6.857143e-02
R37779 n0_12804_7399 n0_12896_7399 6.571429e-02
R37780 n0_12616_15807 n0_12708_15807 1.187097e-01
R37781 n0_12708_15807 n0_12804_15807 1.238710e-01
R37782 n0_12804_15807 n0_12896_15807 1.187097e-01
R37783 n0_12616_17103 n0_12708_17103 1.187097e-01
R37784 n0_12708_17103 n0_12804_17103 1.238710e-01
R37785 n0_12804_17103 n0_12896_17103 1.187097e-01
R37786 n0_12616_19263 n0_12708_19263 1.187097e-01
R37787 n0_12708_19263 n0_12804_19263 1.238710e-01
R37788 n0_12804_19263 n0_12896_19263 1.187097e-01
R37789 n0_12616_5671 n0_12708_5671 6.571429e-02
R37790 n0_12708_5671 n0_12804_5671 6.857143e-02
R37791 n0_12804_5671 n0_12896_5671 6.571429e-02
R37792 n0_12616_6319 n0_12708_6319 6.571429e-02
R37793 n0_12708_6319 n0_12804_6319 6.857143e-02
R37794 n0_12804_6319 n0_12896_6319 6.571429e-02
R37795 n0_12616_3511 n0_12708_3511 6.571429e-02
R37796 n0_12708_3511 n0_12804_3511 6.857143e-02
R37797 n0_12804_3511 n0_12896_3511 6.571429e-02
R37798 n0_12616_4159 n0_12708_4159 6.571429e-02
R37799 n0_12708_4159 n0_12804_4159 6.857143e-02
R37800 n0_12804_4159 n0_12896_4159 6.571429e-02
R37801 n0_12616_4591 n0_12708_4591 6.571429e-02
R37802 n0_12708_4591 n0_12804_4591 6.857143e-02
R37803 n0_12804_4591 n0_12896_4591 6.571429e-02
R37804 n0_12616_15368 n0_12708_15368 2.300000e-01
R37805 n0_12708_15368 n0_12804_15368 2.400000e-01
R37806 n0_12804_15368 n0_12896_15368 2.300000e-01
R37807 n0_12616_18608 n0_12708_18608 2.300000e-01
R37808 n0_12708_18608 n0_12804_18608 2.400000e-01
R37809 n0_12804_18608 n0_12896_18608 2.300000e-01
R37810 n0_12616_1783 n0_12708_1783 6.571429e-02
R37811 n0_12708_1783 n0_12804_1783 6.857143e-02
R37812 n0_12804_1783 n0_12896_1783 6.571429e-02
R37813 n0_12616_16448 n0_12708_16448 2.300000e-01
R37814 n0_12708_16448 n0_12804_16448 2.400000e-01
R37815 n0_12804_16448 n0_12896_16448 2.300000e-01
R37816 n0_12896_16448 n0_14866_16448 4.925000e+00
R37817 n0_14866_16448 n0_14958_16448 2.300000e-01
R37818 n0_14958_16448 n0_15054_16448 2.400000e-01
R37819 n0_15054_16448 n0_15146_16448 2.300000e-01
R37820 n0_12616_17528 n0_12708_17528 2.300000e-01
R37821 n0_12708_17528 n0_12804_17528 2.400000e-01
R37822 n0_12804_17528 n0_12896_17528 2.300000e-01
R37823 n0_12896_17528 n0_14866_17528 4.925000e+00
R37824 n0_14866_17528 n0_14958_17528 2.300000e-01
R37825 n0_14958_17528 n0_15054_17528 2.400000e-01
R37826 n0_15054_17528 n0_15146_17528 2.300000e-01
R37827 n0_12616_18176 n0_12708_18176 2.300000e-01
R37828 n0_12708_18176 n0_12804_18176 2.400000e-01
R37829 n0_12804_18176 n0_12896_18176 2.300000e-01
R37830 n0_12896_18176 n0_14866_18176 4.925000e+00
R37831 n0_14866_18176 n0_14958_18176 2.300000e-01
R37832 n0_14958_18176 n0_15054_18176 2.400000e-01
R37833 n0_15054_18176 n0_15146_18176 2.300000e-01
R37834 n0_12616_2863 n0_12708_2863 6.571429e-02
R37835 n0_12708_2863 n0_12804_2863 6.857143e-02
R37836 n0_12804_2863 n0_12896_2863 6.571429e-02
R37837 n0_12896_2863 n0_14866_2863 1.407143e+00
R37838 n0_14866_2863 n0_14958_2863 6.571429e-02
R37839 n0_14958_2863 n0_15054_2863 6.857143e-02
R37840 n0_15054_2863 n0_15146_2863 6.571429e-02
R37841 n0_15146_2863 n0_17116_2863 1.407143e+00
R37842 n0_17116_2863 n0_17208_2863 6.571429e-02
R37843 n0_17208_2863 n0_17304_2863 6.857143e-02
R37844 n0_17304_2863 n0_17396_2863 6.571429e-02
R37845 n0_12616_2431 n0_12708_2431 6.571429e-02
R37846 n0_12708_2431 n0_12804_2431 6.857143e-02
R37847 n0_12804_2431 n0_12896_2431 6.571429e-02
R37848 n0_12896_2431 n0_14866_2431 1.407143e+00
R37849 n0_14866_2431 n0_14958_2431 6.571429e-02
R37850 n0_14958_2431 n0_15054_2431 6.857143e-02
R37851 n0_15054_2431 n0_15146_2431 6.571429e-02
R37852 n0_15146_2431 n0_17116_2431 1.407143e+00
R37853 n0_17116_2431 n0_17208_2431 6.571429e-02
R37854 n0_17208_2431 n0_17304_2431 6.857143e-02
R37855 n0_17304_2431 n0_17396_2431 6.571429e-02
R37856 n0_12616_5023 n0_12708_5023 6.571429e-02
R37857 n0_12708_5023 n0_12755_5023 3.357143e-02
R37858 n0_12755_5023 n0_12804_5023 3.500000e-02
R37859 n0_12804_5023 n0_12896_5023 6.571429e-02
R37860 n0_12616_14079 n0_12708_14079 1.187097e-01
R37861 n0_12708_14079 n0_12804_14079 1.238710e-01
R37862 n0_12804_14079 n0_12896_14079 1.187097e-01
R37863 n0_12616_14727 n0_12708_14727 1.187097e-01
R37864 n0_12708_14727 n0_12804_14727 1.238710e-01
R37865 n0_12804_14727 n0_12896_14727 1.187097e-01
R37866 n0_12616_15800 n0_12708_15800 2.300000e-01
R37867 n0_12708_15800 n0_12804_15800 2.400000e-01
R37868 n0_12804_15800 n0_12896_15800 2.300000e-01
R37869 n0_12616_18183 n0_12708_18183 1.187097e-01
R37870 n0_12708_18183 n0_12804_18183 1.238710e-01
R37871 n0_12804_18183 n0_12896_18183 1.187097e-01
R37872 n0_12616_19256 n0_12708_19256 2.300000e-01
R37873 n0_12708_19256 n0_12804_19256 2.400000e-01
R37874 n0_12804_19256 n0_12896_19256 2.300000e-01
R37875 n0_12616_8695 n0_12804_8695 1.342857e-01
R37876 n0_12804_8695 n0_13741_8695 6.692857e-01
R37877 n0_13741_8695 n0_13929_8695 1.342857e-01
R37878 n0_12616_9775 n0_12804_9775 1.342857e-01
R37879 n0_12804_9775 n0_13741_9775 6.692857e-01
R37880 n0_13741_9775 n0_13929_9775 1.342857e-01
R37881 n0_12616_10832 n0_12804_10832 4.700000e-01
R37882 n0_12804_10832 n0_13741_10832 2.342500e+00
R37883 n0_13741_10832 n0_13929_10832 4.700000e-01
R37884 n0_12616_11912 n0_12804_11912 4.700000e-01
R37885 n0_12804_11912 n0_13741_11912 2.342500e+00
R37886 n0_13741_11912 n0_13929_11912 4.700000e-01
R37887 n0_12616_3943 n0_12708_3943 6.571429e-02
R37888 n0_12708_3943 n0_12804_3943 6.857143e-02
R37889 n0_12804_3943 n0_12896_3943 6.571429e-02
R37890 n0_12896_3943 n0_14866_3943 1.407143e+00
R37891 n0_14866_3943 n0_14958_3943 6.571429e-02
R37892 n0_14958_3943 n0_15054_3943 6.857143e-02
R37893 n0_15054_3943 n0_15146_3943 6.571429e-02
R37894 n0_12616_17983 n0_12708_17983 6.571429e-02
R37895 n0_12708_17983 n0_12804_17983 6.857143e-02
R37896 n0_12804_17983 n0_12896_17983 6.571429e-02
R37897 n0_12896_17983 n0_14866_17983 1.407143e+00
R37898 n0_14866_17983 n0_14958_17983 6.571429e-02
R37899 n0_14958_17983 n0_15054_17983 6.857143e-02
R37900 n0_15054_17983 n0_15146_17983 6.571429e-02
R37901 n0_12616_17096 n0_12708_17096 2.300000e-01
R37902 n0_12708_17096 n0_12804_17096 2.400000e-01
R37903 n0_12804_17096 n0_12896_17096 2.300000e-01
R37904 n0_12896_17096 n0_14866_17096 4.925000e+00
R37905 n0_14866_17096 n0_14958_17096 2.300000e-01
R37906 n0_14958_17096 n0_15054_17096 2.400000e-01
R37907 n0_15054_17096 n0_15146_17096 2.300000e-01
R37908 n0_12616_11048 n0_12804_11048 4.700000e-01
R37909 n0_12804_11048 n0_13741_11048 2.342500e+00
R37910 n0_13741_11048 n0_13929_11048 4.700000e-01
R37911 n0_13929_11048 n0_14866_11048 2.342500e+00
R37912 n0_14866_11048 n0_15054_11048 4.700000e-01
R37913 n0_15054_11048 n0_15991_11048 2.342500e+00
R37914 n0_15991_11048 n0_16179_11048 4.700000e-01
R37915 n0_16179_11048 n0_17116_11048 2.342500e+00
R37916 n0_17116_11048 n0_17304_11048 4.700000e-01
R37917 n0_12616_7831 n0_12708_7831 6.571429e-02
R37918 n0_12708_7831 n0_12804_7831 6.857143e-02
R37919 n0_12804_7831 n0_12896_7831 6.571429e-02
R37920 n0_12896_7831 n0_13741_7831 6.035714e-01
R37921 n0_13741_7831 n0_13929_7831 1.342857e-01
R37922 n0_13929_7831 n0_14866_7831 6.692857e-01
R37923 n0_14866_7831 n0_15054_7831 1.342857e-01
R37924 n0_15054_7831 n0_15991_7831 6.692857e-01
R37925 n0_15991_7831 n0_16179_7831 1.342857e-01
R37926 n0_16179_7831 n0_17116_7831 6.692857e-01
R37927 n0_17116_7831 n0_17304_7831 1.342857e-01
R37928 n0_17304_7831 n0_18241_7831 6.692857e-01
R37929 n0_18241_7831 n0_18429_7831 1.342857e-01
R37930 n0_18429_7831 n0_19366_7831 6.692857e-01
R37931 n0_19366_7831 n0_19554_7831 1.342857e-01
R37932 n0_12616_8911 n0_12804_8911 1.342857e-01
R37933 n0_12804_8911 n0_13741_8911 6.692857e-01
R37934 n0_13741_8911 n0_13929_8911 1.342857e-01
R37935 n0_13929_8911 n0_14866_8911 6.692857e-01
R37936 n0_14866_8911 n0_15054_8911 1.342857e-01
R37937 n0_15054_8911 n0_15991_8911 6.692857e-01
R37938 n0_15991_8911 n0_16179_8911 1.342857e-01
R37939 n0_16179_8911 n0_17116_8911 6.692857e-01
R37940 n0_17116_8911 n0_17304_8911 1.342857e-01
R37941 n0_17304_8911 n0_18241_8911 6.692857e-01
R37942 n0_18241_8911 n0_18429_8911 1.342857e-01
R37943 n0_18429_8911 n0_19366_8911 6.692857e-01
R37944 n0_19366_8911 n0_19554_8911 1.342857e-01
R37945 n0_12616_9991 n0_12804_9991 1.342857e-01
R37946 n0_12804_9991 n0_13741_9991 6.692857e-01
R37947 n0_13741_9991 n0_13929_9991 1.342857e-01
R37948 n0_13929_9991 n0_14866_9991 6.692857e-01
R37949 n0_14866_9991 n0_15054_9991 1.342857e-01
R37950 n0_15054_9991 n0_15991_9991 6.692857e-01
R37951 n0_15991_9991 n0_16179_9991 1.342857e-01
R37952 n0_16179_9991 n0_17116_9991 6.692857e-01
R37953 n0_17116_9991 n0_17304_9991 1.342857e-01
R37954 n0_17304_9991 n0_18241_9991 6.692857e-01
R37955 n0_18241_9991 n0_18429_9991 1.342857e-01
R37956 n0_18429_9991 n0_19366_9991 6.692857e-01
R37957 n0_19366_9991 n0_19554_9991 1.342857e-01
R37958 n0_12616_12128 n0_12804_12128 4.700000e-01
R37959 n0_12804_12128 n0_13741_12128 2.342500e+00
R37960 n0_13741_12128 n0_13929_12128 4.700000e-01
R37961 n0_13929_12128 n0_14866_12128 2.342500e+00
R37962 n0_14866_12128 n0_15054_12128 4.700000e-01
R37963 n0_15054_12128 n0_15991_12128 2.342500e+00
R37964 n0_15991_12128 n0_16179_12128 4.700000e-01
R37965 n0_16179_12128 n0_17116_12128 2.342500e+00
R37966 n0_17116_12128 n0_17304_12128 4.700000e-01
R37967 n0_17304_12128 n0_18241_12128 2.342500e+00
R37968 n0_18241_12128 n0_18429_12128 4.700000e-01
R37969 n0_18429_12128 n0_19366_12128 2.342500e+00
R37970 n0_19366_12128 n0_19554_12128 4.700000e-01
R37971 n0_13741_12992 n0_13929_12992 4.700000e-01
R37972 n0_13929_12992 n0_14866_12992 2.342500e+00
R37973 n0_14866_12992 n0_15054_12992 4.700000e-01
R37974 n0_15054_12992 n0_15991_12992 2.342500e+00
R37975 n0_15991_12992 n0_16179_12992 4.700000e-01
R37976 n0_13741_12776 n0_13880_12776 3.475000e-01
R37977 n0_13880_12776 n0_13929_12776 1.225000e-01
R37978 n0_13929_12776 n0_14866_12776 2.342500e+00
R37979 n0_14866_12776 n0_15005_12776 3.475000e-01
R37980 n0_15005_12776 n0_15054_12776 1.225000e-01
R37981 n0_15054_12776 n0_15991_12776 2.342500e+00
R37982 n0_15991_12776 n0_16130_12776 3.475000e-01
R37983 n0_16130_12776 n0_16179_12776 1.225000e-01
R37984 n0_14866_3511 n0_14958_3511 6.571429e-02
R37985 n0_14958_3511 n0_15054_3511 6.857143e-02
R37986 n0_15054_3511 n0_15146_3511 6.571429e-02
R37987 n0_14866_15368 n0_14958_15368 2.300000e-01
R37988 n0_14958_15368 n0_15054_15368 2.400000e-01
R37989 n0_15054_15368 n0_15146_15368 2.300000e-01
R37990 n0_14866_15800 n0_14958_15800 2.300000e-01
R37991 n0_14958_15800 n0_15054_15800 2.400000e-01
R37992 n0_15054_15800 n0_15146_15800 2.300000e-01
R37993 n0_14866_19263 n0_14958_19263 1.187097e-01
R37994 n0_14958_19263 n0_15054_19263 1.238710e-01
R37995 n0_15054_19263 n0_15146_19263 1.187097e-01
R37996 n0_14866_1783 n0_14958_1783 6.571429e-02
R37997 n0_14958_1783 n0_15054_1783 6.857143e-02
R37998 n0_15054_1783 n0_15146_1783 6.571429e-02
R37999 n0_14866_18608 n0_14958_18608 2.300000e-01
R38000 n0_14958_18608 n0_15054_18608 2.400000e-01
R38001 n0_15054_18608 n0_15146_18608 2.300000e-01
R38002 n0_14866_14511 n0_15054_14511 2.425806e-01
R38003 n0_15054_14511 n0_15991_14511 1.209032e+00
R38004 n0_15991_14511 n0_16179_14511 2.425806e-01
R38005 n0_16179_14511 n0_17116_14511 1.209032e+00
R38006 n0_17116_14511 n0_17304_14511 2.425806e-01
R38007 n0_17304_14511 n0_18241_14511 1.209032e+00
R38008 n0_18241_14511 n0_18429_14511 2.425806e-01
R38009 n0_18429_14511 n0_19366_14511 1.209032e+00
R38010 n0_19366_14511 n0_19554_14511 2.425806e-01
R38011 n0_14866_5671 n0_14958_5671 6.571429e-02
R38012 n0_14958_5671 n0_15054_5671 6.857143e-02
R38013 n0_15054_5671 n0_15146_5671 6.571429e-02
R38014 n0_14866_6535 n0_15054_6535 1.342857e-01
R38015 n0_14866_4159 n0_14958_4159 6.571429e-02
R38016 n0_14958_4159 n0_15054_4159 6.857143e-02
R38017 n0_15054_4159 n0_15146_4159 6.571429e-02
R38018 n0_14866_4591 n0_14958_4591 6.571429e-02
R38019 n0_14958_4591 n0_15054_4591 6.857143e-02
R38020 n0_15054_4591 n0_15146_4591 6.571429e-02
R38021 n0_14866_5239 n0_14958_5239 6.571429e-02
R38022 n0_14958_5239 n0_15054_5239 6.857143e-02
R38023 n0_15054_5239 n0_15146_5239 6.571429e-02
R38024 n0_15146_5239 n0_15991_5239 6.035714e-01
R38025 n0_15991_5239 n0_16179_5239 1.342857e-01
R38026 n0_16179_5239 n0_17116_5239 6.692857e-01
R38027 n0_17116_5239 n0_17304_5239 1.342857e-01
R38028 n0_17304_5239 n0_18241_5239 6.692857e-01
R38029 n0_18241_5239 n0_18429_5239 1.342857e-01
R38030 n0_18429_5239 n0_19366_5239 6.692857e-01
R38031 n0_19366_5239 n0_19554_5239 1.342857e-01
R38032 n0_14866_3295 n0_14958_3295 6.571429e-02
R38033 n0_14958_3295 n0_15054_3295 6.857143e-02
R38034 n0_15054_3295 n0_15146_3295 6.571429e-02
R38035 n0_14866_4375 n0_14958_4375 6.571429e-02
R38036 n0_14958_4375 n0_15054_4375 6.857143e-02
R38037 n0_15054_4375 n0_15146_4375 6.571429e-02
R38038 n0_14866_19256 n0_14958_19256 2.300000e-01
R38039 n0_14958_19256 n0_15054_19256 2.400000e-01
R38040 n0_15054_19256 n0_15146_19256 2.300000e-01
R38041 n0_14866_12135 n0_15054_12135 2.425806e-01
R38042 n0_15054_12135 n0_15991_12135 1.209032e+00
R38043 n0_15991_12135 n0_16179_12135 2.425806e-01
R38044 n0_16179_12135 n0_17116_12135 1.209032e+00
R38045 n0_17116_12135 n0_17304_12135 2.425806e-01
R38046 n0_14866_14943 n0_15054_14943 2.425806e-01
R38047 n0_15054_14943 n0_15991_14943 1.209032e+00
R38048 n0_15991_14943 n0_16179_14943 2.425806e-01
R38049 n0_16179_14943 n0_17116_14943 1.209032e+00
R38050 n0_17116_14943 n0_17304_14943 2.425806e-01
R38051 n0_14866_16687 n0_14958_16687 6.571429e-02
R38052 n0_14958_16687 n0_15054_16687 6.857143e-02
R38053 n0_15054_16687 n0_15146_16687 6.571429e-02
R38054 n0_15146_16687 n0_17116_16687 1.407143e+00
R38055 n0_17116_16687 n0_17304_16687 1.342857e-01
R38056 n0_14866_15159 n0_14958_15159 1.187097e-01
R38057 n0_14958_15159 n0_15005_15159 6.064516e-02
R38058 n0_15005_15159 n0_15054_15159 6.322581e-02
R38059 n0_15054_15159 n0_15146_15159 1.187097e-01
R38060 n0_15146_15159 n0_15991_15159 1.090323e+00
R38061 n0_15991_15159 n0_16130_15159 1.793548e-01
R38062 n0_16130_15159 n0_16179_15159 6.322581e-02
R38063 n0_16179_15159 n0_17116_15159 1.209032e+00
R38064 n0_17116_15159 n0_17255_15159 1.793548e-01
R38065 n0_17255_15159 n0_17304_15159 6.322581e-02
R38066 n0_14866_4807 n0_14958_4807 6.571429e-02
R38067 n0_14958_4807 n0_15054_4807 6.857143e-02
R38068 n0_15054_4807 n0_15146_4807 6.571429e-02
R38069 n0_15146_4807 n0_17116_4807 1.407143e+00
R38070 n0_17116_4807 n0_17304_4807 1.342857e-01
R38071 n0_17304_4807 n0_18241_4807 6.692857e-01
R38072 n0_18241_4807 n0_18429_4807 1.342857e-01
R38073 n0_14866_5455 n0_14958_5455 6.571429e-02
R38074 n0_14958_5455 n0_15054_5455 6.857143e-02
R38075 n0_15054_5455 n0_15146_5455 6.571429e-02
R38076 n0_15146_5455 n0_15991_5455 6.035714e-01
R38077 n0_15991_5455 n0_16179_5455 1.342857e-01
R38078 n0_16179_5455 n0_17116_5455 6.692857e-01
R38079 n0_17116_5455 n0_17304_5455 1.342857e-01
R38080 n0_17304_5455 n0_18241_5455 6.692857e-01
R38081 n0_18241_5455 n0_18429_5455 1.342857e-01
R38082 n0_18429_5455 n0_19366_5455 6.692857e-01
R38083 n0_19366_5455 n0_19554_5455 1.342857e-01
R38084 n0_14866_15584 n0_14958_15584 2.300000e-01
R38085 n0_14958_15584 n0_15054_15584 2.400000e-01
R38086 n0_15054_15584 n0_15146_15584 2.300000e-01
R38087 n0_15146_15584 n0_15991_15584 2.112500e+00
R38088 n0_15991_15584 n0_16179_15584 4.700000e-01
R38089 n0_16179_15584 n0_17116_15584 2.342500e+00
R38090 n0_17116_15584 n0_17304_15584 4.700000e-01
R38091 n0_17304_15584 n0_18241_15584 2.342500e+00
R38092 n0_18241_15584 n0_18429_15584 4.700000e-01
R38093 n0_18429_15584 n0_19366_15584 2.342500e+00
R38094 n0_19366_15584 n0_19554_15584 4.700000e-01
R38095 n0_14866_6319 n0_15054_6319 1.342857e-01
R38096 n0_15054_6319 n0_15991_6319 6.692857e-01
R38097 n0_15991_6319 n0_16179_6319 1.342857e-01
R38098 n0_16179_6319 n0_17116_6319 6.692857e-01
R38099 n0_17116_6319 n0_17304_6319 1.342857e-01
R38100 n0_17304_6319 n0_18241_6319 6.692857e-01
R38101 n0_18241_6319 n0_18429_6319 1.342857e-01
R38102 n0_18429_6319 n0_19366_6319 6.692857e-01
R38103 n0_19366_6319 n0_19554_6319 1.342857e-01
R38104 n0_19554_6319 n0_20491_6319 6.692857e-01
R38105 n0_20491_6319 n0_20679_6319 1.342857e-01
R38106 n0_15991_13647 n0_16179_13647 2.425806e-01
R38107 n0_16179_13647 n0_17116_13647 1.209032e+00
R38108 n0_17116_13647 n0_17304_13647 2.425806e-01
R38109 n0_15991_5023 n0_17116_5023 8.035714e-01
R38110 n0_17116_5023 n0_18241_5023 8.035714e-01
R38111 n0_17116_17535 n0_17208_17535 1.187097e-01
R38112 n0_17208_17535 n0_17304_17535 1.238710e-01
R38113 n0_17304_17535 n0_17396_17535 1.187097e-01
R38114 n0_17116_18176 n0_17208_18176 2.300000e-01
R38115 n0_17208_18176 n0_17304_18176 2.400000e-01
R38116 n0_17304_18176 n0_17396_18176 2.300000e-01
R38117 n0_17116_19040 n0_17208_19040 2.300000e-01
R38118 n0_17208_19040 n0_17304_19040 2.400000e-01
R38119 n0_17304_19040 n0_17396_19040 2.300000e-01
R38120 n0_17116_1783 n0_17208_1783 6.571429e-02
R38121 n0_17208_1783 n0_17304_1783 6.857143e-02
R38122 n0_17304_1783 n0_17396_1783 6.571429e-02
R38123 n0_17116_3295 n0_17208_3295 6.571429e-02
R38124 n0_17208_3295 n0_17304_3295 6.857143e-02
R38125 n0_17304_3295 n0_17396_3295 6.571429e-02
R38126 n0_17396_3295 n0_18241_3295 6.035714e-01
R38127 n0_18241_3295 n0_18429_3295 1.342857e-01
R38128 n0_18429_3295 n0_19366_3295 6.692857e-01
R38129 n0_19366_3295 n0_19554_3295 1.342857e-01
R38130 n0_17116_4375 n0_17304_4375 1.342857e-01
R38131 n0_17304_4375 n0_18241_4375 6.692857e-01
R38132 n0_18241_4375 n0_18429_4375 1.342857e-01
R38133 n0_18429_4375 n0_19366_4375 6.692857e-01
R38134 n0_19366_4375 n0_19554_4375 1.342857e-01
R38135 n0_17116_16664 n0_17304_16664 4.700000e-01
R38136 n0_17304_16664 n0_18241_16664 2.342500e+00
R38137 n0_18241_16664 n0_18429_16664 4.700000e-01
R38138 n0_18429_16664 n0_19366_16664 2.342500e+00
R38139 n0_19366_16664 n0_19554_16664 4.700000e-01
R38140 n0_17116_4591 n0_17304_4591 1.342857e-01
R38141 n0_17304_4591 n0_18241_4591 6.692857e-01
R38142 n0_18241_4591 n0_18429_4591 1.342857e-01
R38143 n0_17116_13640 n0_17304_13640 4.700000e-01
R38144 n0_17304_13640 n0_18241_13640 2.342500e+00
R38145 n0_18241_13640 n0_18429_13640 4.700000e-01
R38146 n0_17116_11055 n0_17304_11055 2.425806e-01
R38147 n0_17304_11055 n0_18241_11055 1.209032e+00
R38148 n0_18241_11055 n0_18429_11055 2.425806e-01
R38149 n0_18429_11055 n0_19366_11055 1.209032e+00
R38150 n0_19366_11055 n0_19554_11055 2.425806e-01
R38151 n0_17116_17119 n0_17304_17119 1.342857e-01
R38152 n0_17304_17119 n0_18241_17119 6.692857e-01
R38153 n0_18241_17119 n0_18429_17119 1.342857e-01
R38154 n0_18429_17119 n0_19366_17119 6.692857e-01
R38155 n0_19366_17119 n0_19554_17119 1.342857e-01
R38156 n0_17116_14936 n0_17304_14936 4.700000e-01
R38157 n0_17304_14936 n0_18241_14936 2.342500e+00
R38158 n0_18241_14936 n0_18429_14936 4.700000e-01
R38159 n0_18429_14936 n0_19366_14936 2.342500e+00
R38160 n0_19366_14936 n0_19554_14936 4.700000e-01
R38161 n0_19554_14936 n0_20491_14936 2.342500e+00
R38162 n0_20491_14936 n0_20679_14936 4.700000e-01
R38163 n0_17116_15152 n0_17255_15152 3.475000e-01
R38164 n0_17255_15152 n0_17304_15152 1.225000e-01
R38165 n0_17304_15152 n0_18241_15152 2.342500e+00
R38166 n0_18241_15152 n0_18380_15152 3.475000e-01
R38167 n0_18380_15152 n0_18429_15152 1.225000e-01
R38168 n0_18429_15152 n0_19366_15152 2.342500e+00
R38169 n0_19366_15152 n0_19505_15152 3.475000e-01
R38170 n0_19505_15152 n0_19554_15152 1.225000e-01
R38171 n0_19554_15152 n0_20491_15152 2.342500e+00
R38172 n0_20491_15152 n0_20630_15152 3.475000e-01
R38173 n0_20630_15152 n0_20679_15152 1.225000e-01
R38174 n0_18241_13647 n0_18429_13647 2.425806e-01
R38175 n0_18429_13647 n0_19366_13647 1.209032e+00
R38176 n0_19366_13647 n0_19554_13647 2.425806e-01
R38177 n0_18241_14504 n0_18429_14504 4.700000e-01
R38178 n0_18429_14504 n0_19366_14504 2.342500e+00
R38179 n0_19366_14504 n0_19554_14504 4.700000e-01
R38180 n0_18241_16671 n0_18429_16671 2.425806e-01
R38181 n0_18429_16671 n0_19366_16671 1.209032e+00
R38182 n0_19366_16671 n0_19554_16671 2.425806e-01
R38183 n0_18241_17744 n0_18429_17744 4.700000e-01
R38184 n0_18429_17744 n0_19366_17744 2.342500e+00
R38185 n0_19366_17744 n0_19554_17744 4.700000e-01
R38186 n0_19366_1999 n0_19554_1999 1.342857e-01
R38187 n0_19366_18932 n0_19554_18932 4.700000e-01
R38188 n0_19366_1976 n0_19554_1976 4.700000e-01
R38189 n0_19554_1976 n0_20491_1976 2.342500e+00
R38190 n0_20491_1976 n0_20679_1976 4.700000e-01
R38191 n0_19366_19040 n0_19554_19040 4.700000e-01
R38192 n0_19554_19040 n0_20491_19040 2.342500e+00
R38193 n0_20491_19040 n0_20679_19040 4.700000e-01
R38194 n0_19366_5671 n0_19554_5671 1.342857e-01
R38195 n0_19554_5671 n0_20491_5671 6.692857e-01
R38196 n0_20491_5671 n0_20679_5671 1.342857e-01
R38197 n0_19366_16687 n0_19554_16687 1.342857e-01
R38198 n0_19554_16687 n0_20491_16687 6.692857e-01
R38199 n0_20491_16687 n0_20679_16687 1.342857e-01
R38200 n0_20491_9213 n0_20679_9213 1.074286e+00
R38201 n0_20491_11956 n0_20679_11956 1.074286e+00
rrcc n2_17255_2721 _X_n2_17255_2721 2.500000e-01
va1 _X_n2_1505_10596 0 0
rr1f8 n3_20630_11721 _X_n3_20630_11721 2.500000e-01
rr1ae n3_9380_7221 _X_n3_9380_7221 2.500000e-01
rrce n2_19505_471 _X_n2_19505_471 2.500000e-01
va3 _X_n2_2630_10596 0 0
v21b _X_n3_13880_18471 0 1.8
va5 _X_n2_3755_10596 0 0
v21d _X_n3_13880_16221 0 1.8
* layer: M6,VDD net: 3
R38202 n3_333_383 n3_333_424 2.603175e-02
R38203 n3_333_424 n3_333_431 4.444444e-03
R38204 n3_333_431 n3_333_464 2.095238e-02
R38205 n3_333_464 n3_333_520 3.555556e-02
R38206 n3_333_520 n3_333_647 8.063492e-02
R38207 n3_333_647 n3_333_680 2.095238e-02
R38208 n3_333_680 n3_333_863 1.161905e-01
R38209 n3_333_863 n3_333_896 2.095238e-02
R38210 n3_333_896 n3_333_1079 1.161905e-01
R38211 n3_333_1079 n3_333_1112 2.095238e-02
R38212 n3_333_1112 n3_333_1295 1.161905e-01
R38213 n3_333_1295 n3_333_1328 2.095238e-02
R38214 n3_333_424 n3_380_424 2.984127e-02
R38215 n3_380_424 n3_521_424 8.952381e-02
R38216 n3_333_520 n3_380_520 2.984127e-02
R38217 n3_380_520 n3_521_520 8.952381e-02
R38218 n3_333_2674 n3_380_2674 2.984127e-02
R38219 n3_380_2674 n3_521_2674 8.952381e-02
R38220 n3_333_2770 n3_380_2770 2.984127e-02
R38221 n3_380_2770 n3_521_2770 8.952381e-02
R38222 n3_333_4924 n3_380_4924 2.984127e-02
R38223 n3_380_4924 n3_521_4924 8.952381e-02
R38224 n3_333_5020 n3_380_5020 2.984127e-02
R38225 n3_380_5020 n3_521_5020 8.952381e-02
R38226 n3_333_7174 n3_380_7174 2.984127e-02
R38227 n3_380_7174 n3_521_7174 8.952381e-02
R38228 n3_333_7270 n3_380_7270 2.984127e-02
R38229 n3_380_7270 n3_521_7270 8.952381e-02
R38230 n3_333_9424 n3_380_9424 2.984127e-02
R38231 n3_380_9424 n3_521_9424 8.952381e-02
R38232 n3_333_9520 n3_380_9520 2.984127e-02
R38233 n3_380_9520 n3_521_9520 8.952381e-02
R38234 n3_333_11674 n3_380_11674 2.984127e-02
R38235 n3_380_11674 n3_521_11674 8.952381e-02
R38236 n3_333_11770 n3_380_11770 2.984127e-02
R38237 n3_380_11770 n3_521_11770 8.952381e-02
R38238 n3_333_13924 n3_380_13924 2.984127e-02
R38239 n3_380_13924 n3_521_13924 8.952381e-02
R38240 n3_333_14020 n3_380_14020 2.984127e-02
R38241 n3_380_14020 n3_521_14020 8.952381e-02
R38242 n3_333_16174 n3_380_16174 2.984127e-02
R38243 n3_380_16174 n3_521_16174 8.952381e-02
R38244 n3_333_16270 n3_380_16270 2.984127e-02
R38245 n3_380_16270 n3_521_16270 8.952381e-02
R38246 n3_333_18424 n3_380_18424 2.984127e-02
R38247 n3_380_18424 n3_521_18424 8.952381e-02
R38248 n3_333_18520 n3_380_18520 2.984127e-02
R38249 n3_380_18520 n3_521_18520 8.952381e-02
R38250 n3_333_20674 n3_380_20674 2.984127e-02
R38251 n3_380_20674 n3_521_20674 8.952381e-02
R38252 n3_333_20770 n3_380_20770 2.984127e-02
R38253 n3_380_20770 n3_521_20770 8.952381e-02
R38254 n3_333_1727 n3_333_1760 2.095238e-02
R38255 n3_333_1760 n3_333_1943 1.161905e-01
R38256 n3_333_1943 n3_333_1976 2.095238e-02
R38257 n3_333_1976 n3_333_2159 1.161905e-01
R38258 n3_333_2159 n3_333_2192 2.095238e-02
R38259 n3_333_2192 n3_333_2375 1.161905e-01
R38260 n3_333_2375 n3_333_2408 2.095238e-02
R38261 n3_333_2408 n3_333_2543 8.571429e-02
R38262 n3_333_2543 n3_333_2591 3.047619e-02
R38263 n3_333_2591 n3_333_2624 2.095238e-02
R38264 n3_333_2624 n3_333_2674 3.174603e-02
R38265 n3_333_2674 n3_333_2770 6.095238e-02
R38266 n3_333_2770 n3_333_2807 2.349206e-02
R38267 n3_333_2807 n3_333_2840 2.095238e-02
R38268 n3_333_2840 n3_333_3023 1.161905e-01
R38269 n3_333_3023 n3_333_3056 2.095238e-02
R38270 n3_333_3056 n3_333_3239 1.161905e-01
R38271 n3_333_3239 n3_333_3272 2.095238e-02
R38272 n3_333_3272 n3_333_3455 1.161905e-01
R38273 n3_333_3455 n3_333_3488 2.095238e-02
R38274 n3_333_3488 n3_333_3671 1.161905e-01
R38275 n3_333_3671 n3_333_3704 2.095238e-02
R38276 n3_333_4103 n3_333_4136 2.095238e-02
R38277 n3_333_4136 n3_333_4319 1.161905e-01
R38278 n3_333_4319 n3_333_4352 2.095238e-02
R38279 n3_333_4352 n3_333_4486 8.507937e-02
R38280 n3_333_4486 n3_333_4535 3.111111e-02
R38281 n3_333_4535 n3_333_4568 2.095238e-02
R38282 n3_333_4568 n3_333_4751 1.161905e-01
R38283 n3_333_4751 n3_333_4784 2.095238e-02
R38284 n3_333_4784 n3_333_4924 8.888889e-02
R38285 n3_333_4924 n3_333_4967 2.730159e-02
R38286 n3_333_4967 n3_333_5000 2.095238e-02
R38287 n3_333_5000 n3_333_5020 1.269841e-02
R38288 n3_333_5020 n3_333_5183 1.034921e-01
R38289 n3_333_5183 n3_333_5216 2.095238e-02
R38290 n3_333_5216 n3_333_5399 1.161905e-01
R38291 n3_333_5399 n3_333_5432 2.095238e-02
R38292 n3_333_5432 n3_333_5615 1.161905e-01
R38293 n3_333_5615 n3_333_5648 2.095238e-02
R38294 n3_333_5648 n3_333_5831 1.161905e-01
R38295 n3_333_5831 n3_333_5864 2.095238e-02
R38296 n3_333_6263 n3_333_6296 2.095238e-02
R38297 n3_333_6296 n3_333_6479 1.161905e-01
R38298 n3_333_6479 n3_333_6512 2.095238e-02
R38299 n3_333_6512 n3_333_6695 1.161905e-01
R38300 n3_333_6695 n3_333_6728 2.095238e-02
R38301 n3_333_6728 n3_333_6911 1.161905e-01
R38302 n3_333_6911 n3_333_6944 2.095238e-02
R38303 n3_333_6944 n3_333_7127 1.161905e-01
R38304 n3_333_7127 n3_333_7160 2.095238e-02
R38305 n3_333_7160 n3_333_7174 8.888889e-03
R38306 n3_333_7174 n3_333_7270 6.095238e-02
R38307 n3_333_7270 n3_333_7343 4.634921e-02
R38308 n3_333_7343 n3_333_7376 2.095238e-02
R38309 n3_333_7376 n3_333_7559 1.161905e-01
R38310 n3_333_7559 n3_333_7592 2.095238e-02
R38311 n3_333_7592 n3_333_7775 1.161905e-01
R38312 n3_333_7775 n3_333_7808 2.095238e-02
R38313 n3_333_7808 n3_333_7991 1.161905e-01
R38314 n3_333_7991 n3_333_8024 2.095238e-02
R38315 n3_333_8024 n3_333_8207 1.161905e-01
R38316 n3_333_8207 n3_333_8240 2.095238e-02
R38317 n3_333_8456 n3_333_8639 1.161905e-01
R38318 n3_333_8639 n3_333_8672 2.095238e-02
R38319 n3_333_8672 n3_333_8855 1.161905e-01
R38320 n3_333_8855 n3_333_8888 2.095238e-02
R38321 n3_333_8888 n3_333_9071 1.161905e-01
R38322 n3_333_9071 n3_333_9104 2.095238e-02
R38323 n3_333_9104 n3_333_9287 1.161905e-01
R38324 n3_333_9287 n3_333_9320 2.095238e-02
R38325 n3_333_9320 n3_333_9424 6.603175e-02
R38326 n3_333_9424 n3_333_9503 5.015873e-02
R38327 n3_333_9503 n3_333_9520 1.079365e-02
R38328 n3_333_9520 n3_333_9536 1.015873e-02
R38329 n3_333_9536 n3_333_9719 1.161905e-01
R38330 n3_333_9719 n3_333_9752 2.095238e-02
R38331 n3_333_9752 n3_333_9935 1.161905e-01
R38332 n3_333_9935 n3_333_9968 2.095238e-02
R38333 n3_333_9968 n3_333_10151 1.161905e-01
R38334 n3_333_10151 n3_333_10184 2.095238e-02
R38335 n3_333_10184 n3_333_10367 1.161905e-01
R38336 n3_333_10367 n3_333_10400 2.095238e-02
R38337 n3_333_10799 n3_333_10832 2.095238e-02
R38338 n3_333_10832 n3_333_11015 1.161905e-01
R38339 n3_333_11015 n3_333_11048 2.095238e-02
R38340 n3_333_11048 n3_333_11231 1.161905e-01
R38341 n3_333_11231 n3_333_11264 2.095238e-02
R38342 n3_333_11264 n3_333_11447 1.161905e-01
R38343 n3_333_11447 n3_333_11480 2.095238e-02
R38344 n3_333_11480 n3_333_11663 1.161905e-01
R38345 n3_333_11663 n3_333_11674 6.984127e-03
R38346 n3_333_11674 n3_333_11696 1.396825e-02
R38347 n3_333_11696 n3_333_11770 4.698413e-02
R38348 n3_333_11770 n3_333_11879 6.920635e-02
R38349 n3_333_11879 n3_333_11912 2.095238e-02
R38350 n3_333_11912 n3_333_12095 1.161905e-01
R38351 n3_333_12095 n3_333_12128 2.095238e-02
R38352 n3_333_12128 n3_333_12311 1.161905e-01
R38353 n3_333_12311 n3_333_12344 2.095238e-02
R38354 n3_333_12344 n3_333_12527 1.161905e-01
R38355 n3_333_12527 n3_333_12560 2.095238e-02
R38356 n3_333_12560 n3_333_12743 1.161905e-01
R38357 n3_333_12959 n3_333_12992 2.095238e-02
R38358 n3_333_12992 n3_333_13175 1.161905e-01
R38359 n3_333_13175 n3_333_13208 2.095238e-02
R38360 n3_333_13208 n3_333_13391 1.161905e-01
R38361 n3_333_13391 n3_333_13424 2.095238e-02
R38362 n3_333_13424 n3_333_13607 1.161905e-01
R38363 n3_333_13607 n3_333_13640 2.095238e-02
R38364 n3_333_13640 n3_333_13774 8.507937e-02
R38365 n3_333_13774 n3_333_13823 3.111111e-02
R38366 n3_333_13823 n3_333_13856 2.095238e-02
R38367 n3_333_13856 n3_333_13924 4.317460e-02
R38368 n3_333_13924 n3_333_14020 6.095238e-02
R38369 n3_333_14020 n3_333_14039 1.206349e-02
R38370 n3_333_14039 n3_333_14072 2.095238e-02
R38371 n3_333_14072 n3_333_14255 1.161905e-01
R38372 n3_333_14255 n3_333_14288 2.095238e-02
R38373 n3_333_14288 n3_333_14471 1.161905e-01
R38374 n3_333_14471 n3_333_14504 2.095238e-02
R38375 n3_333_14504 n3_333_14687 1.161905e-01
R38376 n3_333_14687 n3_333_14720 2.095238e-02
R38377 n3_333_14720 n3_333_14903 1.161905e-01
R38378 n3_333_14903 n3_333_14936 2.095238e-02
R38379 n3_333_15335 n3_333_15368 2.095238e-02
R38380 n3_333_15368 n3_333_15551 1.161905e-01
R38381 n3_333_15551 n3_333_15584 2.095238e-02
R38382 n3_333_15584 n3_333_15767 1.161905e-01
R38383 n3_333_15767 n3_333_15800 2.095238e-02
R38384 n3_333_15800 n3_333_15983 1.161905e-01
R38385 n3_333_15983 n3_333_16016 2.095238e-02
R38386 n3_333_16016 n3_333_16174 1.003175e-01
R38387 n3_333_16174 n3_333_16199 1.587302e-02
R38388 n3_333_16199 n3_333_16232 2.095238e-02
R38389 n3_333_16232 n3_333_16270 2.412698e-02
R38390 n3_333_16270 n3_333_16415 9.206349e-02
R38391 n3_333_16415 n3_333_16448 2.095238e-02
R38392 n3_333_16448 n3_333_16631 1.161905e-01
R38393 n3_333_16631 n3_333_16664 2.095238e-02
R38394 n3_333_16664 n3_333_16847 1.161905e-01
R38395 n3_333_16847 n3_333_16880 2.095238e-02
R38396 n3_333_16880 n3_333_17063 1.161905e-01
R38397 n3_333_17063 n3_333_17096 2.095238e-02
R38398 n3_333_17495 n3_333_17528 2.095238e-02
R38399 n3_333_17528 n3_333_17711 1.161905e-01
R38400 n3_333_17711 n3_333_17744 2.095238e-02
R38401 n3_333_17744 n3_333_17927 1.161905e-01
R38402 n3_333_17927 n3_333_17960 2.095238e-02
R38403 n3_333_17960 n3_333_18116 9.904762e-02
R38404 n3_333_18116 n3_333_18143 1.714286e-02
R38405 n3_333_18143 n3_333_18176 2.095238e-02
R38406 n3_333_18176 n3_333_18359 1.161905e-01
R38407 n3_333_18359 n3_333_18392 2.095238e-02
R38408 n3_333_18392 n3_333_18424 2.031746e-02
R38409 n3_333_18424 n3_333_18520 6.095238e-02
R38410 n3_333_18520 n3_333_18527 4.444444e-03
R38411 n3_333_18527 n3_333_18575 3.047619e-02
R38412 n3_333_18575 n3_333_18608 2.095238e-02
R38413 n3_333_18608 n3_333_18791 1.161905e-01
R38414 n3_333_18791 n3_333_18824 2.095238e-02
R38415 n3_333_18824 n3_333_19007 1.161905e-01
R38416 n3_333_19007 n3_333_19040 2.095238e-02
R38417 n3_333_19040 n3_333_19196 9.904762e-02
R38418 n3_333_19196 n3_333_19223 1.714286e-02
R38419 n3_333_19223 n3_333_19256 2.095238e-02
R38420 n3_333_19256 n3_333_19412 9.904762e-02
R38421 n3_333_19412 n3_333_19439 1.714286e-02
R38422 n3_333_19439 n3_333_19472 2.095238e-02
R38423 n3_333_19871 n3_333_19904 2.095238e-02
R38424 n3_333_19904 n3_333_20087 1.161905e-01
R38425 n3_333_20087 n3_333_20120 2.095238e-02
R38426 n3_333_20120 n3_333_20303 1.161905e-01
R38427 n3_333_20303 n3_333_20336 2.095238e-02
R38428 n3_333_20336 n3_333_20519 1.161905e-01
R38429 n3_333_20519 n3_333_20552 2.095238e-02
R38430 n3_333_20552 n3_333_20674 7.746032e-02
R38431 n3_333_20674 n3_333_20687 8.253968e-03
R38432 n3_333_20687 n3_333_20735 3.047619e-02
R38433 n3_333_20735 n3_333_20768 2.095238e-02
R38434 n3_333_20768 n3_333_20770 1.269841e-03
R38435 n3_521_215 n3_521_248 2.095238e-02
R38436 n3_521_248 n3_521_383 8.571429e-02
R38437 n3_521_383 n3_521_424 2.603175e-02
R38438 n3_521_424 n3_521_431 4.444444e-03
R38439 n3_521_520 n3_521_647 8.063492e-02
R38440 n3_521_647 n3_521_680 2.095238e-02
R38441 n3_521_680 n3_521_863 1.161905e-01
R38442 n3_521_863 n3_521_896 2.095238e-02
R38443 n3_521_896 n3_521_1079 1.161905e-01
R38444 n3_521_1079 n3_521_1112 2.095238e-02
R38445 n3_521_1112 n3_521_1295 1.161905e-01
R38446 n3_521_1295 n3_521_1328 2.095238e-02
R38447 n3_521_1328 n3_521_1511 1.161905e-01
R38448 n3_521_1511 n3_521_1544 2.095238e-02
R38449 n3_521_1544 n3_521_1727 1.161905e-01
R38450 n3_521_1727 n3_521_1760 2.095238e-02
R38451 n3_521_1760 n3_521_1943 1.161905e-01
R38452 n3_521_1943 n3_521_1976 2.095238e-02
R38453 n3_521_1976 n3_521_2159 1.161905e-01
R38454 n3_521_2159 n3_521_2192 2.095238e-02
R38455 n3_521_2192 n3_521_2375 1.161905e-01
R38456 n3_521_2375 n3_521_2408 2.095238e-02
R38457 n3_521_2408 n3_521_2543 8.571429e-02
R38458 n3_521_2543 n3_521_2591 3.047619e-02
R38459 n3_521_2591 n3_521_2624 2.095238e-02
R38460 n3_521_2624 n3_521_2674 3.174603e-02
R38461 n3_521_2770 n3_521_2807 2.349206e-02
R38462 n3_521_2807 n3_521_2840 2.095238e-02
R38463 n3_521_2840 n3_521_3023 1.161905e-01
R38464 n3_521_3023 n3_521_3056 2.095238e-02
R38465 n3_521_3056 n3_521_3239 1.161905e-01
R38466 n3_521_3239 n3_521_3272 2.095238e-02
R38467 n3_521_3272 n3_521_3455 1.161905e-01
R38468 n3_521_3455 n3_521_3488 2.095238e-02
R38469 n3_521_3488 n3_521_3671 1.161905e-01
R38470 n3_521_3671 n3_521_3704 2.095238e-02
R38471 n3_521_3704 n3_521_3887 1.161905e-01
R38472 n3_521_3887 n3_521_3920 2.095238e-02
R38473 n3_521_3920 n3_521_4103 1.161905e-01
R38474 n3_521_4103 n3_521_4136 2.095238e-02
R38475 n3_521_4136 n3_521_4319 1.161905e-01
R38476 n3_521_4319 n3_521_4352 2.095238e-02
R38477 n3_521_4352 n3_521_4486 8.507937e-02
R38478 n3_521_4486 n3_521_4535 3.111111e-02
R38479 n3_521_4535 n3_521_4568 2.095238e-02
R38480 n3_521_4568 n3_521_4751 1.161905e-01
R38481 n3_521_4751 n3_521_4784 2.095238e-02
R38482 n3_521_4784 n3_521_4924 8.888889e-02
R38483 n3_521_5000 n3_521_5020 1.269841e-02
R38484 n3_521_5020 n3_521_5183 1.034921e-01
R38485 n3_521_5183 n3_521_5216 2.095238e-02
R38486 n3_521_5216 n3_521_5399 1.161905e-01
R38487 n3_521_5399 n3_521_5432 2.095238e-02
R38488 n3_521_5432 n3_521_5615 1.161905e-01
R38489 n3_521_5615 n3_521_5648 2.095238e-02
R38490 n3_521_5648 n3_521_5831 1.161905e-01
R38491 n3_521_5831 n3_521_5864 2.095238e-02
R38492 n3_521_5864 n3_521_6047 1.161905e-01
R38493 n3_521_6047 n3_521_6080 2.095238e-02
R38494 n3_521_6080 n3_521_6263 1.161905e-01
R38495 n3_521_6263 n3_521_6296 2.095238e-02
R38496 n3_521_6296 n3_521_6479 1.161905e-01
R38497 n3_521_6479 n3_521_6512 2.095238e-02
R38498 n3_521_6512 n3_521_6695 1.161905e-01
R38499 n3_521_6695 n3_521_6728 2.095238e-02
R38500 n3_521_6728 n3_521_6911 1.161905e-01
R38501 n3_521_6911 n3_521_6944 2.095238e-02
R38502 n3_521_6944 n3_521_7127 1.161905e-01
R38503 n3_521_7127 n3_521_7160 2.095238e-02
R38504 n3_521_7160 n3_521_7174 8.888889e-03
R38505 n3_521_7270 n3_521_7343 4.634921e-02
R38506 n3_521_7343 n3_521_7376 2.095238e-02
R38507 n3_521_7376 n3_521_7559 1.161905e-01
R38508 n3_521_7559 n3_521_7592 2.095238e-02
R38509 n3_521_7592 n3_521_7775 1.161905e-01
R38510 n3_521_7775 n3_521_7808 2.095238e-02
R38511 n3_521_7808 n3_521_7991 1.161905e-01
R38512 n3_521_7991 n3_521_8024 2.095238e-02
R38513 n3_521_8024 n3_521_8207 1.161905e-01
R38514 n3_521_8207 n3_521_8240 2.095238e-02
R38515 n3_521_8240 n3_521_8423 1.161905e-01
R38516 n3_521_8423 n3_521_8456 2.095238e-02
R38517 n3_521_8456 n3_521_8639 1.161905e-01
R38518 n3_521_8639 n3_521_8672 2.095238e-02
R38519 n3_521_8672 n3_521_8855 1.161905e-01
R38520 n3_521_8855 n3_521_8888 2.095238e-02
R38521 n3_521_8888 n3_521_9071 1.161905e-01
R38522 n3_521_9071 n3_521_9104 2.095238e-02
R38523 n3_521_9104 n3_521_9287 1.161905e-01
R38524 n3_521_9287 n3_521_9320 2.095238e-02
R38525 n3_521_9320 n3_521_9424 6.603175e-02
R38526 n3_521_9503 n3_521_9520 1.079365e-02
R38527 n3_521_9520 n3_521_9536 1.015873e-02
R38528 n3_521_9536 n3_521_9719 1.161905e-01
R38529 n3_521_9719 n3_521_9752 2.095238e-02
R38530 n3_521_9752 n3_521_9935 1.161905e-01
R38531 n3_521_9935 n3_521_9968 2.095238e-02
R38532 n3_521_9968 n3_521_10151 1.161905e-01
R38533 n3_521_10151 n3_521_10184 2.095238e-02
R38534 n3_521_10184 n3_521_10367 1.161905e-01
R38535 n3_521_10367 n3_521_10400 2.095238e-02
R38536 n3_521_10616 n3_521_10799 1.161905e-01
R38537 n3_521_10799 n3_521_10832 2.095238e-02
R38538 n3_521_10832 n3_521_11015 1.161905e-01
R38539 n3_521_11015 n3_521_11048 2.095238e-02
R38540 n3_521_11048 n3_521_11231 1.161905e-01
R38541 n3_521_11231 n3_521_11264 2.095238e-02
R38542 n3_521_11264 n3_521_11447 1.161905e-01
R38543 n3_521_11447 n3_521_11480 2.095238e-02
R38544 n3_521_11480 n3_521_11663 1.161905e-01
R38545 n3_521_11663 n3_521_11674 6.984127e-03
R38546 n3_521_11674 n3_521_11696 1.396825e-02
R38547 n3_521_11770 n3_521_11879 6.920635e-02
R38548 n3_521_11879 n3_521_11912 2.095238e-02
R38549 n3_521_11912 n3_521_12095 1.161905e-01
R38550 n3_521_12095 n3_521_12128 2.095238e-02
R38551 n3_521_12128 n3_521_12311 1.161905e-01
R38552 n3_521_12311 n3_521_12344 2.095238e-02
R38553 n3_521_12344 n3_521_12527 1.161905e-01
R38554 n3_521_12527 n3_521_12560 2.095238e-02
R38555 n3_521_12560 n3_521_12743 1.161905e-01
R38556 n3_521_12743 n3_521_12776 2.095238e-02
R38557 n3_521_12776 n3_521_12959 1.161905e-01
R38558 n3_521_12959 n3_521_12992 2.095238e-02
R38559 n3_521_12992 n3_521_13175 1.161905e-01
R38560 n3_521_13175 n3_521_13208 2.095238e-02
R38561 n3_521_13208 n3_521_13391 1.161905e-01
R38562 n3_521_13391 n3_521_13424 2.095238e-02
R38563 n3_521_13424 n3_521_13607 1.161905e-01
R38564 n3_521_13607 n3_521_13640 2.095238e-02
R38565 n3_521_13640 n3_521_13774 8.507937e-02
R38566 n3_521_13774 n3_521_13823 3.111111e-02
R38567 n3_521_13823 n3_521_13856 2.095238e-02
R38568 n3_521_13856 n3_521_13924 4.317460e-02
R38569 n3_521_14020 n3_521_14039 1.206349e-02
R38570 n3_521_14039 n3_521_14072 2.095238e-02
R38571 n3_521_14072 n3_521_14255 1.161905e-01
R38572 n3_521_14255 n3_521_14288 2.095238e-02
R38573 n3_521_14288 n3_521_14471 1.161905e-01
R38574 n3_521_14471 n3_521_14504 2.095238e-02
R38575 n3_521_14504 n3_521_14687 1.161905e-01
R38576 n3_521_14687 n3_521_14720 2.095238e-02
R38577 n3_521_14720 n3_521_14903 1.161905e-01
R38578 n3_521_14903 n3_521_14936 2.095238e-02
R38579 n3_521_14936 n3_521_15119 1.161905e-01
R38580 n3_521_15119 n3_521_15152 2.095238e-02
R38581 n3_521_15152 n3_521_15335 1.161905e-01
R38582 n3_521_15335 n3_521_15368 2.095238e-02
R38583 n3_521_15368 n3_521_15551 1.161905e-01
R38584 n3_521_15551 n3_521_15584 2.095238e-02
R38585 n3_521_15584 n3_521_15767 1.161905e-01
R38586 n3_521_15767 n3_521_15800 2.095238e-02
R38587 n3_521_15800 n3_521_15983 1.161905e-01
R38588 n3_521_15983 n3_521_16016 2.095238e-02
R38589 n3_521_16016 n3_521_16174 1.003175e-01
R38590 n3_521_16174 n3_521_16199 1.587302e-02
R38591 n3_521_16270 n3_521_16415 9.206349e-02
R38592 n3_521_16415 n3_521_16448 2.095238e-02
R38593 n3_521_16448 n3_521_16631 1.161905e-01
R38594 n3_521_16631 n3_521_16664 2.095238e-02
R38595 n3_521_16664 n3_521_16847 1.161905e-01
R38596 n3_521_16847 n3_521_16880 2.095238e-02
R38597 n3_521_16880 n3_521_17063 1.161905e-01
R38598 n3_521_17063 n3_521_17096 2.095238e-02
R38599 n3_521_17096 n3_521_17279 1.161905e-01
R38600 n3_521_17279 n3_521_17312 2.095238e-02
R38601 n3_521_17312 n3_521_17495 1.161905e-01
R38602 n3_521_17495 n3_521_17528 2.095238e-02
R38603 n3_521_17528 n3_521_17711 1.161905e-01
R38604 n3_521_17711 n3_521_17744 2.095238e-02
R38605 n3_521_17744 n3_521_17927 1.161905e-01
R38606 n3_521_17927 n3_521_17960 2.095238e-02
R38607 n3_521_17960 n3_521_18116 9.904762e-02
R38608 n3_521_18116 n3_521_18143 1.714286e-02
R38609 n3_521_18143 n3_521_18176 2.095238e-02
R38610 n3_521_18176 n3_521_18359 1.161905e-01
R38611 n3_521_18359 n3_521_18392 2.095238e-02
R38612 n3_521_18392 n3_521_18424 2.031746e-02
R38613 n3_521_18520 n3_521_18527 4.444444e-03
R38614 n3_521_18527 n3_521_18575 3.047619e-02
R38615 n3_521_18575 n3_521_18608 2.095238e-02
R38616 n3_521_18608 n3_521_18791 1.161905e-01
R38617 n3_521_18791 n3_521_18824 2.095238e-02
R38618 n3_521_18824 n3_521_19007 1.161905e-01
R38619 n3_521_19007 n3_521_19040 2.095238e-02
R38620 n3_521_19040 n3_521_19196 9.904762e-02
R38621 n3_521_19196 n3_521_19223 1.714286e-02
R38622 n3_521_19223 n3_521_19256 2.095238e-02
R38623 n3_521_19256 n3_521_19412 9.904762e-02
R38624 n3_521_19412 n3_521_19439 1.714286e-02
R38625 n3_521_19439 n3_521_19472 2.095238e-02
R38626 n3_521_19472 n3_521_19655 1.161905e-01
R38627 n3_521_19655 n3_521_19688 2.095238e-02
R38628 n3_521_19688 n3_521_19871 1.161905e-01
R38629 n3_521_19871 n3_521_19904 2.095238e-02
R38630 n3_521_19904 n3_521_20087 1.161905e-01
R38631 n3_521_20087 n3_521_20120 2.095238e-02
R38632 n3_521_20120 n3_521_20303 1.161905e-01
R38633 n3_521_20303 n3_521_20336 2.095238e-02
R38634 n3_521_20336 n3_521_20519 1.161905e-01
R38635 n3_521_20519 n3_521_20552 2.095238e-02
R38636 n3_521_20552 n3_521_20674 7.746032e-02
R38637 n3_521_20674 n3_521_20687 8.253968e-03
R38638 n3_521_20768 n3_521_20770 1.269841e-03
R38639 n3_521_20770 n3_521_20951 1.149206e-01
R38640 n3_521_20951 n3_521_20984 2.095238e-02
R38641 n3_2400_215 n3_2400_248 2.095238e-02
R38642 n3_2400_248 n3_2400_383 8.571429e-02
R38643 n3_2400_383 n3_2400_431 3.047619e-02
R38644 n3_2400_431 n3_2400_464 2.095238e-02
R38645 n3_2400_464 n3_2400_647 1.161905e-01
R38646 n3_2400_647 n3_2400_680 2.095238e-02
R38647 n3_2400_680 n3_2400_863 1.161905e-01
R38648 n3_2400_863 n3_2400_896 2.095238e-02
R38649 n3_2400_896 n3_2400_1079 1.161905e-01
R38650 n3_2400_1079 n3_2400_1112 2.095238e-02
R38651 n3_2400_1112 n3_2400_1295 1.161905e-01
R38652 n3_2400_1295 n3_2400_1328 2.095238e-02
R38653 n3_2400_1328 n3_2400_1511 1.161905e-01
R38654 n3_2400_1511 n3_2400_1544 2.095238e-02
R38655 n3_2400_1544 n3_2400_1727 1.161905e-01
R38656 n3_2400_1727 n3_2400_1760 2.095238e-02
R38657 n3_2400_1760 n3_2400_1943 1.161905e-01
R38658 n3_2400_1943 n3_2400_1976 2.095238e-02
R38659 n3_2400_1976 n3_2400_2159 1.161905e-01
R38660 n3_2400_2159 n3_2400_2192 2.095238e-02
R38661 n3_2400_2192 n3_2400_2375 1.161905e-01
R38662 n3_2400_2375 n3_2400_2408 2.095238e-02
R38663 n3_2400_2408 n3_2400_2543 8.571429e-02
R38664 n3_2400_2543 n3_2400_2591 3.047619e-02
R38665 n3_2400_2591 n3_2400_2624 2.095238e-02
R38666 n3_2400_18527 n3_2400_18575 3.047619e-02
R38667 n3_2400_18575 n3_2400_18608 2.095238e-02
R38668 n3_2400_18608 n3_2400_18791 1.161905e-01
R38669 n3_2400_18791 n3_2400_18824 2.095238e-02
R38670 n3_2400_18824 n3_2400_19007 1.161905e-01
R38671 n3_2400_19007 n3_2400_19040 2.095238e-02
R38672 n3_2400_19040 n3_2400_19223 1.161905e-01
R38673 n3_2400_19223 n3_2400_19256 2.095238e-02
R38674 n3_2400_19256 n3_2400_19439 1.161905e-01
R38675 n3_2400_19439 n3_2400_19472 2.095238e-02
R38676 n3_2400_19472 n3_2400_19655 1.161905e-01
R38677 n3_2400_19655 n3_2400_19688 2.095238e-02
R38678 n3_2400_19688 n3_2400_19871 1.161905e-01
R38679 n3_2400_19871 n3_2400_19904 2.095238e-02
R38680 n3_2400_19904 n3_2400_20087 1.161905e-01
R38681 n3_2400_20087 n3_2400_20120 2.095238e-02
R38682 n3_2400_20120 n3_2400_20303 1.161905e-01
R38683 n3_2400_20303 n3_2400_20336 2.095238e-02
R38684 n3_2400_20336 n3_2400_20519 1.161905e-01
R38685 n3_2400_20519 n3_2400_20552 2.095238e-02
R38686 n3_2400_20552 n3_2400_20687 8.571429e-02
R38687 n3_2400_20687 n3_2400_20735 3.047619e-02
R38688 n3_2400_20735 n3_2400_20768 2.095238e-02
R38689 n3_2400_20768 n3_2400_20951 1.161905e-01
R38690 n3_2400_20951 n3_2400_20984 2.095238e-02
R38691 n3_2583_424 n3_2630_424 2.984127e-02
R38692 n3_2630_424 n3_2771_424 8.952381e-02
R38693 n3_2583_520 n3_2630_520 2.984127e-02
R38694 n3_2630_520 n3_2771_520 8.952381e-02
R38695 n3_2583_2674 n3_2630_2674 2.984127e-02
R38696 n3_2630_2674 n3_2771_2674 8.952381e-02
R38697 n3_2583_2770 n3_2630_2770 2.984127e-02
R38698 n3_2630_2770 n3_2771_2770 8.952381e-02
R38699 n3_2583_4924 n3_2630_4924 2.984127e-02
R38700 n3_2630_4924 n3_2771_4924 8.952381e-02
R38701 n3_2583_5020 n3_2630_5020 2.984127e-02
R38702 n3_2630_5020 n3_2771_5020 8.952381e-02
R38703 n3_2583_7174 n3_2630_7174 2.984127e-02
R38704 n3_2630_7174 n3_2771_7174 8.952381e-02
R38705 n3_2583_7270 n3_2630_7270 2.984127e-02
R38706 n3_2630_7270 n3_2771_7270 8.952381e-02
R38707 n3_2583_9424 n3_2630_9424 2.984127e-02
R38708 n3_2630_9424 n3_2771_9424 8.952381e-02
R38709 n3_2583_9520 n3_2630_9520 2.984127e-02
R38710 n3_2630_9520 n3_2771_9520 8.952381e-02
R38711 n3_2583_11674 n3_2630_11674 2.984127e-02
R38712 n3_2630_11674 n3_2771_11674 8.952381e-02
R38713 n3_2583_11770 n3_2630_11770 2.984127e-02
R38714 n3_2630_11770 n3_2771_11770 8.952381e-02
R38715 n3_2583_13924 n3_2630_13924 2.984127e-02
R38716 n3_2630_13924 n3_2771_13924 8.952381e-02
R38717 n3_2583_14020 n3_2630_14020 2.984127e-02
R38718 n3_2630_14020 n3_2771_14020 8.952381e-02
R38719 n3_2583_16174 n3_2630_16174 2.984127e-02
R38720 n3_2630_16174 n3_2771_16174 8.952381e-02
R38721 n3_2583_16270 n3_2630_16270 2.984127e-02
R38722 n3_2630_16270 n3_2771_16270 8.952381e-02
R38723 n3_2583_18424 n3_2630_18424 2.984127e-02
R38724 n3_2630_18424 n3_2771_18424 8.952381e-02
R38725 n3_2583_18520 n3_2630_18520 2.984127e-02
R38726 n3_2630_18520 n3_2771_18520 8.952381e-02
R38727 n3_2583_20674 n3_2630_20674 2.984127e-02
R38728 n3_2630_20674 n3_2771_20674 8.952381e-02
R38729 n3_2583_20770 n3_2630_20770 2.984127e-02
R38730 n3_2630_20770 n3_2771_20770 8.952381e-02
R38731 n3_2583_215 n3_2583_248 2.095238e-02
R38732 n3_2583_248 n3_2583_383 8.571429e-02
R38733 n3_2583_383 n3_2583_424 2.603175e-02
R38734 n3_2583_424 n3_2583_431 4.444444e-03
R38735 n3_2583_431 n3_2583_464 2.095238e-02
R38736 n3_2583_464 n3_2583_520 3.555556e-02
R38737 n3_2583_520 n3_2583_647 8.063492e-02
R38738 n3_2583_647 n3_2583_680 2.095238e-02
R38739 n3_2583_680 n3_2583_863 1.161905e-01
R38740 n3_2583_863 n3_2583_896 2.095238e-02
R38741 n3_2583_896 n3_2583_1079 1.161905e-01
R38742 n3_2583_1079 n3_2583_1112 2.095238e-02
R38743 n3_2583_1112 n3_2583_1295 1.161905e-01
R38744 n3_2583_1295 n3_2583_1328 2.095238e-02
R38745 n3_2583_1727 n3_2583_1760 2.095238e-02
R38746 n3_2583_1760 n3_2583_1943 1.161905e-01
R38747 n3_2583_1943 n3_2583_1976 2.095238e-02
R38748 n3_2583_1976 n3_2583_2159 1.161905e-01
R38749 n3_2583_2159 n3_2583_2192 2.095238e-02
R38750 n3_2583_2192 n3_2583_2375 1.161905e-01
R38751 n3_2583_2375 n3_2583_2408 2.095238e-02
R38752 n3_2583_2408 n3_2583_2543 8.571429e-02
R38753 n3_2583_2543 n3_2583_2591 3.047619e-02
R38754 n3_2583_2591 n3_2583_2624 2.095238e-02
R38755 n3_2583_2624 n3_2583_2674 3.174603e-02
R38756 n3_2583_2674 n3_2583_2770 6.095238e-02
R38757 n3_2583_2770 n3_2583_2807 2.349206e-02
R38758 n3_2583_2807 n3_2583_2840 2.095238e-02
R38759 n3_2583_2840 n3_2583_3023 1.161905e-01
R38760 n3_2583_3023 n3_2583_3056 2.095238e-02
R38761 n3_2583_3056 n3_2583_3239 1.161905e-01
R38762 n3_2583_3239 n3_2583_3272 2.095238e-02
R38763 n3_2583_3272 n3_2583_3428 9.904762e-02
R38764 n3_2583_3428 n3_2583_3455 1.714286e-02
R38765 n3_2583_3455 n3_2583_3488 2.095238e-02
R38766 n3_2583_3488 n3_2583_3671 1.161905e-01
R38767 n3_2583_3671 n3_2583_3704 2.095238e-02
R38768 n3_2583_4076 n3_2583_4103 1.714286e-02
R38769 n3_2583_4103 n3_2583_4136 2.095238e-02
R38770 n3_2583_4136 n3_2583_4270 8.507937e-02
R38771 n3_2583_4270 n3_2583_4319 3.111111e-02
R38772 n3_2583_4319 n3_2583_4352 2.095238e-02
R38773 n3_2583_4352 n3_2583_4508 9.904762e-02
R38774 n3_2583_4508 n3_2583_4535 1.714286e-02
R38775 n3_2583_4535 n3_2583_4568 2.095238e-02
R38776 n3_2583_4568 n3_2583_4751 1.161905e-01
R38777 n3_2583_4751 n3_2583_4784 2.095238e-02
R38778 n3_2583_4784 n3_2583_4924 8.888889e-02
R38779 n3_2583_4924 n3_2583_4967 2.730159e-02
R38780 n3_2583_4967 n3_2583_5000 2.095238e-02
R38781 n3_2583_5000 n3_2583_5020 1.269841e-02
R38782 n3_2583_5020 n3_2583_5183 1.034921e-01
R38783 n3_2583_5183 n3_2583_5216 2.095238e-02
R38784 n3_2583_5216 n3_2583_5399 1.161905e-01
R38785 n3_2583_5399 n3_2583_5432 2.095238e-02
R38786 n3_2583_5432 n3_2583_5446 8.888889e-03
R38787 n3_2583_5446 n3_2583_5588 9.015873e-02
R38788 n3_2583_5588 n3_2583_5615 1.714286e-02
R38789 n3_2583_5615 n3_2583_5648 2.095238e-02
R38790 n3_2583_5648 n3_2583_5831 1.161905e-01
R38791 n3_2583_5831 n3_2583_5864 2.095238e-02
R38792 n3_2583_6263 n3_2583_6296 2.095238e-02
R38793 n3_2583_6296 n3_2583_6479 1.161905e-01
R38794 n3_2583_6479 n3_2583_6512 2.095238e-02
R38795 n3_2583_6512 n3_2583_6549 2.349206e-02
R38796 n3_2583_6549 n3_2583_6646 6.158730e-02
R38797 n3_2583_6646 n3_2583_6695 3.111111e-02
R38798 n3_2583_6695 n3_2583_6728 2.095238e-02
R38799 n3_2583_6728 n3_2583_6911 1.161905e-01
R38800 n3_2583_6911 n3_2583_6944 2.095238e-02
R38801 n3_2583_6944 n3_2583_7127 1.161905e-01
R38802 n3_2583_7127 n3_2583_7160 2.095238e-02
R38803 n3_2583_7160 n3_2583_7174 8.888889e-03
R38804 n3_2583_7174 n3_2583_7270 6.095238e-02
R38805 n3_2583_7270 n3_2583_7343 4.634921e-02
R38806 n3_2583_7343 n3_2583_7376 2.095238e-02
R38807 n3_2583_7376 n3_2583_7559 1.161905e-01
R38808 n3_2583_7559 n3_2583_7592 2.095238e-02
R38809 n3_2583_7592 n3_2583_7775 1.161905e-01
R38810 n3_2583_7775 n3_2583_7808 2.095238e-02
R38811 n3_2583_7808 n3_2583_7822 8.888889e-03
R38812 n3_2583_7822 n3_2583_7964 9.015873e-02
R38813 n3_2583_7964 n3_2583_7991 1.714286e-02
R38814 n3_2583_7991 n3_2583_8024 2.095238e-02
R38815 n3_2583_8024 n3_2583_8207 1.161905e-01
R38816 n3_2583_8207 n3_2583_8240 2.095238e-02
R38817 n3_2583_8456 n3_2583_8639 1.161905e-01
R38818 n3_2583_8639 n3_2583_8672 2.095238e-02
R38819 n3_2583_8672 n3_2583_8855 1.161905e-01
R38820 n3_2583_8855 n3_2583_8888 2.095238e-02
R38821 n3_2583_8888 n3_2583_8902 8.888889e-03
R38822 n3_2583_8902 n3_2583_9022 7.619048e-02
R38823 n3_2583_9022 n3_2583_9044 1.396825e-02
R38824 n3_2583_9044 n3_2583_9071 1.714286e-02
R38825 n3_2583_9071 n3_2583_9104 2.095238e-02
R38826 n3_2583_9104 n3_2583_9287 1.161905e-01
R38827 n3_2583_9287 n3_2583_9320 2.095238e-02
R38828 n3_2583_9320 n3_2583_9424 6.603175e-02
R38829 n3_2583_9424 n3_2583_9503 5.015873e-02
R38830 n3_2583_9503 n3_2583_9520 1.079365e-02
R38831 n3_2583_9520 n3_2583_9536 1.015873e-02
R38832 n3_2583_9536 n3_2583_9719 1.161905e-01
R38833 n3_2583_9719 n3_2583_9752 2.095238e-02
R38834 n3_2583_9752 n3_2583_9935 1.161905e-01
R38835 n3_2583_9935 n3_2583_9968 2.095238e-02
R38836 n3_2583_9968 n3_2583_9982 8.888889e-03
R38837 n3_2583_9982 n3_2583_10124 9.015873e-02
R38838 n3_2583_10124 n3_2583_10151 1.714286e-02
R38839 n3_2583_10151 n3_2583_10184 2.095238e-02
R38840 n3_2583_10184 n3_2583_10367 1.161905e-01
R38841 n3_2583_10367 n3_2583_10400 2.095238e-02
R38842 n3_2583_10799 n3_2583_10832 2.095238e-02
R38843 n3_2583_10832 n3_2583_11015 1.161905e-01
R38844 n3_2583_11015 n3_2583_11048 2.095238e-02
R38845 n3_2583_11048 n3_2583_11182 8.507937e-02
R38846 n3_2583_11182 n3_2583_11204 1.396825e-02
R38847 n3_2583_11204 n3_2583_11231 1.714286e-02
R38848 n3_2583_11231 n3_2583_11264 2.095238e-02
R38849 n3_2583_11264 n3_2583_11447 1.161905e-01
R38850 n3_2583_11447 n3_2583_11480 2.095238e-02
R38851 n3_2583_11480 n3_2583_11663 1.161905e-01
R38852 n3_2583_11663 n3_2583_11674 6.984127e-03
R38853 n3_2583_11674 n3_2583_11696 1.396825e-02
R38854 n3_2583_11696 n3_2583_11770 4.698413e-02
R38855 n3_2583_11770 n3_2583_11879 6.920635e-02
R38856 n3_2583_11879 n3_2583_11912 2.095238e-02
R38857 n3_2583_11912 n3_2583_12095 1.161905e-01
R38858 n3_2583_12095 n3_2583_12128 2.095238e-02
R38859 n3_2583_12128 n3_2583_12262 8.507937e-02
R38860 n3_2583_12262 n3_2583_12284 1.396825e-02
R38861 n3_2583_12284 n3_2583_12311 1.714286e-02
R38862 n3_2583_12311 n3_2583_12344 2.095238e-02
R38863 n3_2583_12344 n3_2583_12527 1.161905e-01
R38864 n3_2583_12527 n3_2583_12560 2.095238e-02
R38865 n3_2583_12560 n3_2583_12743 1.161905e-01
R38866 n3_2583_12959 n3_2583_12992 2.095238e-02
R38867 n3_2583_12992 n3_2583_13175 1.161905e-01
R38868 n3_2583_13175 n3_2583_13208 2.095238e-02
R38869 n3_2583_13208 n3_2583_13391 1.161905e-01
R38870 n3_2583_13391 n3_2583_13424 2.095238e-02
R38871 n3_2583_13424 n3_2583_13558 8.507937e-02
R38872 n3_2583_13558 n3_2583_13580 1.396825e-02
R38873 n3_2583_13580 n3_2583_13607 1.714286e-02
R38874 n3_2583_13607 n3_2583_13640 2.095238e-02
R38875 n3_2583_13640 n3_2583_13796 9.904762e-02
R38876 n3_2583_13796 n3_2583_13823 1.714286e-02
R38877 n3_2583_13823 n3_2583_13856 2.095238e-02
R38878 n3_2583_13856 n3_2583_13924 4.317460e-02
R38879 n3_2583_13924 n3_2583_13990 4.190476e-02
R38880 n3_2583_13990 n3_2583_14020 1.904762e-02
R38881 n3_2583_14020 n3_2583_14039 1.206349e-02
R38882 n3_2583_14039 n3_2583_14072 2.095238e-02
R38883 n3_2583_14072 n3_2583_14206 8.507937e-02
R38884 n3_2583_14206 n3_2583_14255 3.111111e-02
R38885 n3_2583_14255 n3_2583_14288 2.095238e-02
R38886 n3_2583_14288 n3_2583_14471 1.161905e-01
R38887 n3_2583_14471 n3_2583_14504 2.095238e-02
R38888 n3_2583_14504 n3_2583_14660 9.904762e-02
R38889 n3_2583_14660 n3_2583_14687 1.714286e-02
R38890 n3_2583_14687 n3_2583_14720 2.095238e-02
R38891 n3_2583_14720 n3_2583_14903 1.161905e-01
R38892 n3_2583_14903 n3_2583_14936 2.095238e-02
R38893 n3_2583_15335 n3_2583_15368 2.095238e-02
R38894 n3_2583_15368 n3_2583_15524 9.904762e-02
R38895 n3_2583_15524 n3_2583_15551 1.714286e-02
R38896 n3_2583_15551 n3_2583_15584 2.095238e-02
R38897 n3_2583_15584 n3_2583_15740 9.904762e-02
R38898 n3_2583_15740 n3_2583_15767 1.714286e-02
R38899 n3_2583_15767 n3_2583_15800 2.095238e-02
R38900 n3_2583_15800 n3_2583_15983 1.161905e-01
R38901 n3_2583_15983 n3_2583_16016 2.095238e-02
R38902 n3_2583_16016 n3_2583_16174 1.003175e-01
R38903 n3_2583_16174 n3_2583_16199 1.587302e-02
R38904 n3_2583_16199 n3_2583_16232 2.095238e-02
R38905 n3_2583_16232 n3_2583_16270 2.412698e-02
R38906 n3_2583_16270 n3_2583_16415 9.206349e-02
R38907 n3_2583_16415 n3_2583_16448 2.095238e-02
R38908 n3_2583_16448 n3_2583_16582 8.507937e-02
R38909 n3_2583_16582 n3_2583_16631 3.111111e-02
R38910 n3_2583_16631 n3_2583_16664 2.095238e-02
R38911 n3_2583_16664 n3_2583_16798 8.507937e-02
R38912 n3_2583_16798 n3_2583_16820 1.396825e-02
R38913 n3_2583_16820 n3_2583_16847 1.714286e-02
R38914 n3_2583_16847 n3_2583_16880 2.095238e-02
R38915 n3_2583_16880 n3_2583_17036 9.904762e-02
R38916 n3_2583_17036 n3_2583_17063 1.714286e-02
R38917 n3_2583_17063 n3_2583_17096 2.095238e-02
R38918 n3_2583_17495 n3_2583_17528 2.095238e-02
R38919 n3_2583_17528 n3_2583_17662 8.507937e-02
R38920 n3_2583_17662 n3_2583_17684 1.396825e-02
R38921 n3_2583_17684 n3_2583_17711 1.714286e-02
R38922 n3_2583_17711 n3_2583_17744 2.095238e-02
R38923 n3_2583_17744 n3_2583_17927 1.161905e-01
R38924 n3_2583_17927 n3_2583_17960 2.095238e-02
R38925 n3_2583_17960 n3_2583_18143 1.161905e-01
R38926 n3_2583_18143 n3_2583_18176 2.095238e-02
R38927 n3_2583_18176 n3_2583_18359 1.161905e-01
R38928 n3_2583_18359 n3_2583_18392 2.095238e-02
R38929 n3_2583_18392 n3_2583_18424 2.031746e-02
R38930 n3_2583_18424 n3_2583_18520 6.095238e-02
R38931 n3_2583_18520 n3_2583_18527 4.444444e-03
R38932 n3_2583_18527 n3_2583_18575 3.047619e-02
R38933 n3_2583_18575 n3_2583_18608 2.095238e-02
R38934 n3_2583_18608 n3_2583_18791 1.161905e-01
R38935 n3_2583_18791 n3_2583_18824 2.095238e-02
R38936 n3_2583_18824 n3_2583_19007 1.161905e-01
R38937 n3_2583_19007 n3_2583_19040 2.095238e-02
R38938 n3_2583_19040 n3_2583_19223 1.161905e-01
R38939 n3_2583_19223 n3_2583_19256 2.095238e-02
R38940 n3_2583_19256 n3_2583_19439 1.161905e-01
R38941 n3_2583_19439 n3_2583_19472 2.095238e-02
R38942 n3_2583_19871 n3_2583_19904 2.095238e-02
R38943 n3_2583_19904 n3_2583_20087 1.161905e-01
R38944 n3_2583_20087 n3_2583_20120 2.095238e-02
R38945 n3_2583_20120 n3_2583_20303 1.161905e-01
R38946 n3_2583_20303 n3_2583_20336 2.095238e-02
R38947 n3_2583_20336 n3_2583_20519 1.161905e-01
R38948 n3_2583_20519 n3_2583_20552 2.095238e-02
R38949 n3_2583_20552 n3_2583_20674 7.746032e-02
R38950 n3_2583_20674 n3_2583_20687 8.253968e-03
R38951 n3_2583_20687 n3_2583_20735 3.047619e-02
R38952 n3_2583_20735 n3_2583_20768 2.095238e-02
R38953 n3_2583_20768 n3_2583_20770 1.269841e-03
R38954 n3_2583_20770 n3_2583_20951 1.149206e-01
R38955 n3_2583_20951 n3_2583_20984 2.095238e-02
R38956 n3_2771_215 n3_2771_248 2.095238e-02
R38957 n3_2771_248 n3_2771_383 8.571429e-02
R38958 n3_2771_383 n3_2771_424 2.603175e-02
R38959 n3_2771_424 n3_2771_431 4.444444e-03
R38960 n3_2771_520 n3_2771_647 8.063492e-02
R38961 n3_2771_647 n3_2771_680 2.095238e-02
R38962 n3_2771_680 n3_2771_863 1.161905e-01
R38963 n3_2771_863 n3_2771_896 2.095238e-02
R38964 n3_2771_896 n3_2771_1079 1.161905e-01
R38965 n3_2771_1079 n3_2771_1112 2.095238e-02
R38966 n3_2771_1112 n3_2771_1295 1.161905e-01
R38967 n3_2771_1295 n3_2771_1328 2.095238e-02
R38968 n3_2771_1328 n3_2771_1511 1.161905e-01
R38969 n3_2771_1511 n3_2771_1544 2.095238e-02
R38970 n3_2771_1544 n3_2771_1727 1.161905e-01
R38971 n3_2771_1727 n3_2771_1760 2.095238e-02
R38972 n3_2771_1760 n3_2771_1943 1.161905e-01
R38973 n3_2771_1943 n3_2771_1976 2.095238e-02
R38974 n3_2771_1976 n3_2771_2159 1.161905e-01
R38975 n3_2771_2159 n3_2771_2192 2.095238e-02
R38976 n3_2771_2192 n3_2771_2375 1.161905e-01
R38977 n3_2771_2375 n3_2771_2408 2.095238e-02
R38978 n3_2771_2408 n3_2771_2543 8.571429e-02
R38979 n3_2771_2543 n3_2771_2591 3.047619e-02
R38980 n3_2771_2591 n3_2771_2624 2.095238e-02
R38981 n3_2771_2624 n3_2771_2674 3.174603e-02
R38982 n3_2771_2770 n3_2771_2807 2.349206e-02
R38983 n3_2771_2807 n3_2771_2840 2.095238e-02
R38984 n3_2771_2840 n3_2771_3023 1.161905e-01
R38985 n3_2771_3023 n3_2771_3056 2.095238e-02
R38986 n3_2771_3056 n3_2771_3239 1.161905e-01
R38987 n3_2771_3239 n3_2771_3272 2.095238e-02
R38988 n3_2771_3272 n3_2771_3428 9.904762e-02
R38989 n3_2771_3428 n3_2771_3455 1.714286e-02
R38990 n3_2771_3455 n3_2771_3488 2.095238e-02
R38991 n3_2771_3488 n3_2771_3671 1.161905e-01
R38992 n3_2771_3671 n3_2771_3704 2.095238e-02
R38993 n3_2771_3704 n3_2771_3860 9.904762e-02
R38994 n3_2771_3860 n3_2771_3887 1.714286e-02
R38995 n3_2771_3887 n3_2771_3920 2.095238e-02
R38996 n3_2771_3920 n3_2771_4076 9.904762e-02
R38997 n3_2771_4076 n3_2771_4103 1.714286e-02
R38998 n3_2771_4103 n3_2771_4136 2.095238e-02
R38999 n3_2771_4136 n3_2771_4270 8.507937e-02
R39000 n3_2771_4270 n3_2771_4319 3.111111e-02
R39001 n3_2771_4319 n3_2771_4352 2.095238e-02
R39002 n3_2771_4352 n3_2771_4508 9.904762e-02
R39003 n3_2771_4508 n3_2771_4535 1.714286e-02
R39004 n3_2771_4535 n3_2771_4568 2.095238e-02
R39005 n3_2771_4568 n3_2771_4751 1.161905e-01
R39006 n3_2771_4751 n3_2771_4784 2.095238e-02
R39007 n3_2771_4784 n3_2771_4924 8.888889e-02
R39008 n3_2771_5000 n3_2771_5020 1.269841e-02
R39009 n3_2771_5020 n3_2771_5183 1.034921e-01
R39010 n3_2771_5183 n3_2771_5216 2.095238e-02
R39011 n3_2771_5216 n3_2771_5399 1.161905e-01
R39012 n3_2771_5399 n3_2771_5432 2.095238e-02
R39013 n3_2771_5432 n3_2771_5446 8.888889e-03
R39014 n3_2771_5446 n3_2771_5588 9.015873e-02
R39015 n3_2771_5588 n3_2771_5615 1.714286e-02
R39016 n3_2771_5615 n3_2771_5648 2.095238e-02
R39017 n3_2771_5648 n3_2771_5831 1.161905e-01
R39018 n3_2771_5831 n3_2771_5864 2.095238e-02
R39019 n3_2771_5864 n3_2771_6047 1.161905e-01
R39020 n3_2771_6047 n3_2771_6080 2.095238e-02
R39021 n3_2771_6080 n3_2771_6263 1.161905e-01
R39022 n3_2771_6263 n3_2771_6296 2.095238e-02
R39023 n3_2771_6296 n3_2771_6479 1.161905e-01
R39024 n3_2771_6479 n3_2771_6512 2.095238e-02
R39025 n3_2771_6512 n3_2771_6549 2.349206e-02
R39026 n3_2771_6549 n3_2771_6646 6.158730e-02
R39027 n3_2771_6646 n3_2771_6695 3.111111e-02
R39028 n3_2771_6695 n3_2771_6728 2.095238e-02
R39029 n3_2771_6728 n3_2771_6911 1.161905e-01
R39030 n3_2771_6911 n3_2771_6944 2.095238e-02
R39031 n3_2771_6944 n3_2771_7127 1.161905e-01
R39032 n3_2771_7127 n3_2771_7160 2.095238e-02
R39033 n3_2771_7160 n3_2771_7174 8.888889e-03
R39034 n3_2771_7270 n3_2771_7343 4.634921e-02
R39035 n3_2771_7343 n3_2771_7376 2.095238e-02
R39036 n3_2771_7376 n3_2771_7559 1.161905e-01
R39037 n3_2771_7559 n3_2771_7592 2.095238e-02
R39038 n3_2771_7592 n3_2771_7775 1.161905e-01
R39039 n3_2771_7775 n3_2771_7808 2.095238e-02
R39040 n3_2771_7808 n3_2771_7822 8.888889e-03
R39041 n3_2771_7822 n3_2771_7964 9.015873e-02
R39042 n3_2771_7964 n3_2771_7991 1.714286e-02
R39043 n3_2771_7991 n3_2771_8024 2.095238e-02
R39044 n3_2771_8024 n3_2771_8207 1.161905e-01
R39045 n3_2771_8207 n3_2771_8240 2.095238e-02
R39046 n3_2771_8240 n3_2771_8423 1.161905e-01
R39047 n3_2771_8423 n3_2771_8456 2.095238e-02
R39048 n3_2771_8456 n3_2771_8639 1.161905e-01
R39049 n3_2771_8639 n3_2771_8672 2.095238e-02
R39050 n3_2771_8672 n3_2771_8855 1.161905e-01
R39051 n3_2771_8855 n3_2771_8888 2.095238e-02
R39052 n3_2771_8888 n3_2771_8902 8.888889e-03
R39053 n3_2771_8902 n3_2771_9022 7.619048e-02
R39054 n3_2771_9022 n3_2771_9044 1.396825e-02
R39055 n3_2771_9044 n3_2771_9071 1.714286e-02
R39056 n3_2771_9071 n3_2771_9104 2.095238e-02
R39057 n3_2771_9104 n3_2771_9287 1.161905e-01
R39058 n3_2771_9287 n3_2771_9320 2.095238e-02
R39059 n3_2771_9320 n3_2771_9424 6.603175e-02
R39060 n3_2771_9503 n3_2771_9520 1.079365e-02
R39061 n3_2771_9520 n3_2771_9536 1.015873e-02
R39062 n3_2771_9536 n3_2771_9719 1.161905e-01
R39063 n3_2771_9719 n3_2771_9752 2.095238e-02
R39064 n3_2771_9752 n3_2771_9935 1.161905e-01
R39065 n3_2771_9935 n3_2771_9968 2.095238e-02
R39066 n3_2771_9968 n3_2771_9982 8.888889e-03
R39067 n3_2771_9982 n3_2771_10124 9.015873e-02
R39068 n3_2771_10124 n3_2771_10151 1.714286e-02
R39069 n3_2771_10151 n3_2771_10184 2.095238e-02
R39070 n3_2771_10184 n3_2771_10367 1.161905e-01
R39071 n3_2771_10367 n3_2771_10400 2.095238e-02
R39072 n3_2771_10616 n3_2771_10799 1.161905e-01
R39073 n3_2771_10799 n3_2771_10832 2.095238e-02
R39074 n3_2771_10832 n3_2771_11015 1.161905e-01
R39075 n3_2771_11015 n3_2771_11048 2.095238e-02
R39076 n3_2771_11048 n3_2771_11182 8.507937e-02
R39077 n3_2771_11182 n3_2771_11204 1.396825e-02
R39078 n3_2771_11204 n3_2771_11231 1.714286e-02
R39079 n3_2771_11231 n3_2771_11264 2.095238e-02
R39080 n3_2771_11264 n3_2771_11447 1.161905e-01
R39081 n3_2771_11447 n3_2771_11480 2.095238e-02
R39082 n3_2771_11480 n3_2771_11663 1.161905e-01
R39083 n3_2771_11663 n3_2771_11674 6.984127e-03
R39084 n3_2771_11674 n3_2771_11696 1.396825e-02
R39085 n3_2771_11770 n3_2771_11879 6.920635e-02
R39086 n3_2771_11879 n3_2771_11912 2.095238e-02
R39087 n3_2771_11912 n3_2771_12095 1.161905e-01
R39088 n3_2771_12095 n3_2771_12128 2.095238e-02
R39089 n3_2771_12128 n3_2771_12262 8.507937e-02
R39090 n3_2771_12262 n3_2771_12284 1.396825e-02
R39091 n3_2771_12284 n3_2771_12311 1.714286e-02
R39092 n3_2771_12311 n3_2771_12344 2.095238e-02
R39093 n3_2771_12344 n3_2771_12527 1.161905e-01
R39094 n3_2771_12527 n3_2771_12560 2.095238e-02
R39095 n3_2771_12560 n3_2771_12743 1.161905e-01
R39096 n3_2771_12743 n3_2771_12776 2.095238e-02
R39097 n3_2771_12776 n3_2771_12959 1.161905e-01
R39098 n3_2771_12959 n3_2771_12992 2.095238e-02
R39099 n3_2771_12992 n3_2771_13175 1.161905e-01
R39100 n3_2771_13175 n3_2771_13208 2.095238e-02
R39101 n3_2771_13208 n3_2771_13391 1.161905e-01
R39102 n3_2771_13391 n3_2771_13424 2.095238e-02
R39103 n3_2771_13424 n3_2771_13558 8.507937e-02
R39104 n3_2771_13558 n3_2771_13580 1.396825e-02
R39105 n3_2771_13580 n3_2771_13607 1.714286e-02
R39106 n3_2771_13607 n3_2771_13640 2.095238e-02
R39107 n3_2771_13640 n3_2771_13796 9.904762e-02
R39108 n3_2771_13796 n3_2771_13823 1.714286e-02
R39109 n3_2771_13823 n3_2771_13856 2.095238e-02
R39110 n3_2771_13856 n3_2771_13924 4.317460e-02
R39111 n3_2771_13990 n3_2771_14020 1.904762e-02
R39112 n3_2771_14020 n3_2771_14039 1.206349e-02
R39113 n3_2771_14039 n3_2771_14072 2.095238e-02
R39114 n3_2771_14072 n3_2771_14206 8.507937e-02
R39115 n3_2771_14206 n3_2771_14255 3.111111e-02
R39116 n3_2771_14255 n3_2771_14288 2.095238e-02
R39117 n3_2771_14288 n3_2771_14471 1.161905e-01
R39118 n3_2771_14471 n3_2771_14504 2.095238e-02
R39119 n3_2771_14504 n3_2771_14660 9.904762e-02
R39120 n3_2771_14660 n3_2771_14687 1.714286e-02
R39121 n3_2771_14687 n3_2771_14720 2.095238e-02
R39122 n3_2771_14720 n3_2771_14903 1.161905e-01
R39123 n3_2771_14903 n3_2771_14936 2.095238e-02
R39124 n3_2771_14936 n3_2771_15119 1.161905e-01
R39125 n3_2771_15119 n3_2771_15152 2.095238e-02
R39126 n3_2771_15152 n3_2771_15335 1.161905e-01
R39127 n3_2771_15335 n3_2771_15368 2.095238e-02
R39128 n3_2771_15368 n3_2771_15524 9.904762e-02
R39129 n3_2771_15524 n3_2771_15551 1.714286e-02
R39130 n3_2771_15551 n3_2771_15584 2.095238e-02
R39131 n3_2771_15584 n3_2771_15740 9.904762e-02
R39132 n3_2771_15740 n3_2771_15767 1.714286e-02
R39133 n3_2771_15767 n3_2771_15800 2.095238e-02
R39134 n3_2771_15800 n3_2771_15983 1.161905e-01
R39135 n3_2771_15983 n3_2771_16016 2.095238e-02
R39136 n3_2771_16016 n3_2771_16174 1.003175e-01
R39137 n3_2771_16174 n3_2771_16199 1.587302e-02
R39138 n3_2771_16270 n3_2771_16415 9.206349e-02
R39139 n3_2771_16415 n3_2771_16448 2.095238e-02
R39140 n3_2771_16448 n3_2771_16582 8.507937e-02
R39141 n3_2771_16582 n3_2771_16631 3.111111e-02
R39142 n3_2771_16631 n3_2771_16664 2.095238e-02
R39143 n3_2771_16664 n3_2771_16798 8.507937e-02
R39144 n3_2771_16798 n3_2771_16820 1.396825e-02
R39145 n3_2771_16820 n3_2771_16847 1.714286e-02
R39146 n3_2771_16847 n3_2771_16880 2.095238e-02
R39147 n3_2771_16880 n3_2771_17036 9.904762e-02
R39148 n3_2771_17036 n3_2771_17063 1.714286e-02
R39149 n3_2771_17063 n3_2771_17096 2.095238e-02
R39150 n3_2771_17096 n3_2771_17279 1.161905e-01
R39151 n3_2771_17279 n3_2771_17312 2.095238e-02
R39152 n3_2771_17312 n3_2771_17495 1.161905e-01
R39153 n3_2771_17495 n3_2771_17528 2.095238e-02
R39154 n3_2771_17528 n3_2771_17662 8.507937e-02
R39155 n3_2771_17662 n3_2771_17684 1.396825e-02
R39156 n3_2771_17684 n3_2771_17711 1.714286e-02
R39157 n3_2771_17711 n3_2771_17744 2.095238e-02
R39158 n3_2771_17744 n3_2771_17927 1.161905e-01
R39159 n3_2771_17927 n3_2771_17960 2.095238e-02
R39160 n3_2771_17960 n3_2771_18143 1.161905e-01
R39161 n3_2771_18143 n3_2771_18176 2.095238e-02
R39162 n3_2771_18176 n3_2771_18359 1.161905e-01
R39163 n3_2771_18359 n3_2771_18392 2.095238e-02
R39164 n3_2771_18392 n3_2771_18424 2.031746e-02
R39165 n3_2771_18520 n3_2771_18527 4.444444e-03
R39166 n3_2771_18527 n3_2771_18575 3.047619e-02
R39167 n3_2771_18575 n3_2771_18608 2.095238e-02
R39168 n3_2771_18608 n3_2771_18791 1.161905e-01
R39169 n3_2771_18791 n3_2771_18824 2.095238e-02
R39170 n3_2771_18824 n3_2771_19007 1.161905e-01
R39171 n3_2771_19007 n3_2771_19040 2.095238e-02
R39172 n3_2771_19040 n3_2771_19223 1.161905e-01
R39173 n3_2771_19223 n3_2771_19256 2.095238e-02
R39174 n3_2771_19256 n3_2771_19439 1.161905e-01
R39175 n3_2771_19439 n3_2771_19472 2.095238e-02
R39176 n3_2771_19472 n3_2771_19655 1.161905e-01
R39177 n3_2771_19655 n3_2771_19688 2.095238e-02
R39178 n3_2771_19688 n3_2771_19871 1.161905e-01
R39179 n3_2771_19871 n3_2771_19904 2.095238e-02
R39180 n3_2771_19904 n3_2771_20087 1.161905e-01
R39181 n3_2771_20087 n3_2771_20120 2.095238e-02
R39182 n3_2771_20120 n3_2771_20303 1.161905e-01
R39183 n3_2771_20303 n3_2771_20336 2.095238e-02
R39184 n3_2771_20336 n3_2771_20519 1.161905e-01
R39185 n3_2771_20519 n3_2771_20552 2.095238e-02
R39186 n3_2771_20552 n3_2771_20674 7.746032e-02
R39187 n3_2771_20674 n3_2771_20687 8.253968e-03
R39188 n3_2771_20768 n3_2771_20770 1.269841e-03
R39189 n3_2771_20770 n3_2771_20951 1.149206e-01
R39190 n3_2771_20951 n3_2771_20984 2.095238e-02
R39191 n3_2864_215 n3_2864_248 2.095238e-02
R39192 n3_2864_248 n3_2864_383 8.571429e-02
R39193 n3_2864_383 n3_2864_431 3.047619e-02
R39194 n3_2864_431 n3_2864_464 2.095238e-02
R39195 n3_2864_464 n3_2864_647 1.161905e-01
R39196 n3_2864_647 n3_2864_680 2.095238e-02
R39197 n3_2864_680 n3_2864_863 1.161905e-01
R39198 n3_2864_863 n3_2864_896 2.095238e-02
R39199 n3_2864_896 n3_2864_1079 1.161905e-01
R39200 n3_2864_1079 n3_2864_1112 2.095238e-02
R39201 n3_2864_1112 n3_2864_1295 1.161905e-01
R39202 n3_2864_1295 n3_2864_1328 2.095238e-02
R39203 n3_2864_1328 n3_2864_1511 1.161905e-01
R39204 n3_2864_1511 n3_2864_1544 2.095238e-02
R39205 n3_2864_1544 n3_2864_1727 1.161905e-01
R39206 n3_2864_1727 n3_2864_1760 2.095238e-02
R39207 n3_2864_1760 n3_2864_1943 1.161905e-01
R39208 n3_2864_1943 n3_2864_1976 2.095238e-02
R39209 n3_2864_1976 n3_2864_2159 1.161905e-01
R39210 n3_2864_2159 n3_2864_2192 2.095238e-02
R39211 n3_2864_2192 n3_2864_2375 1.161905e-01
R39212 n3_2864_2375 n3_2864_2408 2.095238e-02
R39213 n3_2864_2408 n3_2864_2543 8.571429e-02
R39214 n3_2864_2543 n3_2864_2591 3.047619e-02
R39215 n3_2864_2591 n3_2864_2624 2.095238e-02
R39216 n3_2864_18527 n3_2864_18575 3.047619e-02
R39217 n3_2864_18575 n3_2864_18608 2.095238e-02
R39218 n3_2864_18608 n3_2864_18791 1.161905e-01
R39219 n3_2864_18791 n3_2864_18824 2.095238e-02
R39220 n3_2864_18824 n3_2864_19007 1.161905e-01
R39221 n3_2864_19007 n3_2864_19040 2.095238e-02
R39222 n3_2864_19040 n3_2864_19223 1.161905e-01
R39223 n3_2864_19223 n3_2864_19256 2.095238e-02
R39224 n3_2864_19256 n3_2864_19439 1.161905e-01
R39225 n3_2864_19439 n3_2864_19472 2.095238e-02
R39226 n3_2864_19472 n3_2864_19655 1.161905e-01
R39227 n3_2864_19655 n3_2864_19688 2.095238e-02
R39228 n3_2864_19688 n3_2864_19871 1.161905e-01
R39229 n3_2864_19871 n3_2864_19904 2.095238e-02
R39230 n3_2864_19904 n3_2864_20087 1.161905e-01
R39231 n3_2864_20087 n3_2864_20120 2.095238e-02
R39232 n3_2864_20120 n3_2864_20303 1.161905e-01
R39233 n3_2864_20303 n3_2864_20336 2.095238e-02
R39234 n3_2864_20336 n3_2864_20519 1.161905e-01
R39235 n3_2864_20519 n3_2864_20552 2.095238e-02
R39236 n3_2864_20552 n3_2864_20687 8.571429e-02
R39237 n3_2864_20687 n3_2864_20735 3.047619e-02
R39238 n3_2864_20735 n3_2864_20768 2.095238e-02
R39239 n3_2864_20768 n3_2864_20951 1.161905e-01
R39240 n3_2864_20951 n3_2864_20984 2.095238e-02
R39241 n3_4650_215 n3_4650_248 2.095238e-02
R39242 n3_4650_248 n3_4650_431 1.161905e-01
R39243 n3_4650_431 n3_4650_464 2.095238e-02
R39244 n3_4650_464 n3_4650_513 3.111111e-02
R39245 n3_4650_513 n3_4650_647 8.507937e-02
R39246 n3_4650_647 n3_4650_680 2.095238e-02
R39247 n3_4650_680 n3_4650_863 1.161905e-01
R39248 n3_4650_863 n3_4650_896 2.095238e-02
R39249 n3_4650_896 n3_4650_945 3.111111e-02
R39250 n3_4650_945 n3_4650_1079 8.507937e-02
R39251 n3_4650_1079 n3_4650_1112 2.095238e-02
R39252 n3_4650_1112 n3_4650_1295 1.161905e-01
R39253 n3_4650_1295 n3_4650_1328 2.095238e-02
R39254 n3_4650_1328 n3_4650_1511 1.161905e-01
R39255 n3_4650_1511 n3_4650_1544 2.095238e-02
R39256 n3_4650_1544 n3_4650_1727 1.161905e-01
R39257 n3_4650_1727 n3_4650_1760 2.095238e-02
R39258 n3_4650_1760 n3_4650_1943 1.161905e-01
R39259 n3_4650_1943 n3_4650_1976 2.095238e-02
R39260 n3_4650_1976 n3_4650_2132 9.904762e-02
R39261 n3_4650_2132 n3_4650_2159 1.714286e-02
R39262 n3_4650_2159 n3_4650_2192 2.095238e-02
R39263 n3_4650_2192 n3_4650_2375 1.161905e-01
R39264 n3_4650_2375 n3_4650_2408 2.095238e-02
R39265 n3_4650_2408 n3_4650_2543 8.571429e-02
R39266 n3_4650_2543 n3_4650_2591 3.047619e-02
R39267 n3_4650_2591 n3_4650_2624 2.095238e-02
R39268 n3_4650_18527 n3_4650_18575 3.047619e-02
R39269 n3_4650_18575 n3_4650_18608 2.095238e-02
R39270 n3_4650_18608 n3_4650_18791 1.161905e-01
R39271 n3_4650_18791 n3_4650_18824 2.095238e-02
R39272 n3_4650_18824 n3_4650_19007 1.161905e-01
R39273 n3_4650_19007 n3_4650_19040 2.095238e-02
R39274 n3_4650_19040 n3_4650_19223 1.161905e-01
R39275 n3_4650_19223 n3_4650_19256 2.095238e-02
R39276 n3_4650_19256 n3_4650_19439 1.161905e-01
R39277 n3_4650_19439 n3_4650_19472 2.095238e-02
R39278 n3_4650_19472 n3_4650_19655 1.161905e-01
R39279 n3_4650_19655 n3_4650_19688 2.095238e-02
R39280 n3_4650_19688 n3_4650_19871 1.161905e-01
R39281 n3_4650_19871 n3_4650_19904 2.095238e-02
R39282 n3_4650_19904 n3_4650_20087 1.161905e-01
R39283 n3_4650_20087 n3_4650_20120 2.095238e-02
R39284 n3_4650_20120 n3_4650_20303 1.161905e-01
R39285 n3_4650_20303 n3_4650_20336 2.095238e-02
R39286 n3_4650_20336 n3_4650_20519 1.161905e-01
R39287 n3_4650_20519 n3_4650_20552 2.095238e-02
R39288 n3_4650_20552 n3_4650_20687 8.571429e-02
R39289 n3_4650_20687 n3_4650_20735 3.047619e-02
R39290 n3_4650_20735 n3_4650_20768 2.095238e-02
R39291 n3_4650_20768 n3_4650_20951 1.161905e-01
R39292 n3_4650_20951 n3_4650_20984 2.095238e-02
R39293 n3_4833_424 n3_4880_424 2.984127e-02
R39294 n3_4880_424 n3_5021_424 8.952381e-02
R39295 n3_4833_520 n3_4880_520 2.984127e-02
R39296 n3_4880_520 n3_5021_520 8.952381e-02
R39297 n3_4833_2674 n3_4880_2674 2.984127e-02
R39298 n3_4880_2674 n3_5021_2674 8.952381e-02
R39299 n3_4833_2770 n3_4880_2770 2.984127e-02
R39300 n3_4880_2770 n3_5021_2770 8.952381e-02
R39301 n3_4833_4924 n3_4880_4924 2.984127e-02
R39302 n3_4880_4924 n3_5021_4924 8.952381e-02
R39303 n3_4833_5020 n3_4880_5020 2.984127e-02
R39304 n3_4880_5020 n3_5021_5020 8.952381e-02
R39305 n3_4833_7174 n3_4880_7174 2.984127e-02
R39306 n3_4880_7174 n3_5021_7174 8.952381e-02
R39307 n3_4833_7270 n3_4880_7270 2.984127e-02
R39308 n3_4880_7270 n3_5021_7270 8.952381e-02
R39309 n3_4833_9424 n3_4880_9424 2.984127e-02
R39310 n3_4880_9424 n3_5021_9424 8.952381e-02
R39311 n3_4833_9520 n3_4880_9520 2.984127e-02
R39312 n3_4880_9520 n3_5021_9520 8.952381e-02
R39313 n3_4833_11674 n3_4880_11674 2.984127e-02
R39314 n3_4880_11674 n3_5021_11674 8.952381e-02
R39315 n3_4833_11770 n3_4880_11770 2.984127e-02
R39316 n3_4880_11770 n3_5021_11770 8.952381e-02
R39317 n3_4833_13924 n3_4880_13924 2.984127e-02
R39318 n3_4880_13924 n3_5021_13924 8.952381e-02
R39319 n3_4833_14020 n3_4880_14020 2.984127e-02
R39320 n3_4880_14020 n3_5021_14020 8.952381e-02
R39321 n3_4833_16174 n3_4880_16174 2.984127e-02
R39322 n3_4880_16174 n3_5021_16174 8.952381e-02
R39323 n3_4833_16270 n3_4880_16270 2.984127e-02
R39324 n3_4880_16270 n3_5021_16270 8.952381e-02
R39325 n3_4833_18424 n3_4880_18424 2.984127e-02
R39326 n3_4880_18424 n3_5021_18424 8.952381e-02
R39327 n3_4833_18520 n3_4880_18520 2.984127e-02
R39328 n3_4880_18520 n3_5021_18520 8.952381e-02
R39329 n3_4833_20674 n3_4880_20674 2.984127e-02
R39330 n3_4880_20674 n3_5021_20674 8.952381e-02
R39331 n3_4833_20770 n3_4880_20770 2.984127e-02
R39332 n3_4880_20770 n3_5021_20770 8.952381e-02
R39333 n3_4833_215 n3_4833_248 2.095238e-02
R39334 n3_4833_248 n3_4833_424 1.117460e-01
R39335 n3_4833_424 n3_4833_431 4.444444e-03
R39336 n3_4833_431 n3_4833_464 2.095238e-02
R39337 n3_4833_464 n3_4833_513 3.111111e-02
R39338 n3_4833_513 n3_4833_520 4.444444e-03
R39339 n3_4833_520 n3_4833_647 8.063492e-02
R39340 n3_4833_647 n3_4833_680 2.095238e-02
R39341 n3_4833_680 n3_4833_863 1.161905e-01
R39342 n3_4833_863 n3_4833_896 2.095238e-02
R39343 n3_4833_896 n3_4833_945 3.111111e-02
R39344 n3_4833_945 n3_4833_1079 8.507937e-02
R39345 n3_4833_1079 n3_4833_1112 2.095238e-02
R39346 n3_4833_1112 n3_4833_1295 1.161905e-01
R39347 n3_4833_1295 n3_4833_1328 2.095238e-02
R39348 n3_4833_1727 n3_4833_1760 2.095238e-02
R39349 n3_4833_1760 n3_4833_1916 9.904762e-02
R39350 n3_4833_1916 n3_4833_1943 1.714286e-02
R39351 n3_4833_1943 n3_4833_1976 2.095238e-02
R39352 n3_4833_1976 n3_4833_2132 9.904762e-02
R39353 n3_4833_2132 n3_4833_2159 1.714286e-02
R39354 n3_4833_2159 n3_4833_2192 2.095238e-02
R39355 n3_4833_2192 n3_4833_2375 1.161905e-01
R39356 n3_4833_2375 n3_4833_2408 2.095238e-02
R39357 n3_4833_2408 n3_4833_2543 8.571429e-02
R39358 n3_4833_2543 n3_4833_2564 1.333333e-02
R39359 n3_4833_2564 n3_4833_2591 1.714286e-02
R39360 n3_4833_2591 n3_4833_2624 2.095238e-02
R39361 n3_4833_2624 n3_4833_2674 3.174603e-02
R39362 n3_4833_2674 n3_4833_2770 6.095238e-02
R39363 n3_4833_2770 n3_4833_2807 2.349206e-02
R39364 n3_4833_2807 n3_4833_2840 2.095238e-02
R39365 n3_4833_2840 n3_4833_2996 9.904762e-02
R39366 n3_4833_2996 n3_4833_3023 1.714286e-02
R39367 n3_4833_3023 n3_4833_3056 2.095238e-02
R39368 n3_4833_3056 n3_4833_3212 9.904762e-02
R39369 n3_4833_3212 n3_4833_3239 1.714286e-02
R39370 n3_4833_3239 n3_4833_3272 2.095238e-02
R39371 n3_4833_3272 n3_4833_3455 1.161905e-01
R39372 n3_4833_3455 n3_4833_3488 2.095238e-02
R39373 n3_4833_3488 n3_4833_3644 9.904762e-02
R39374 n3_4833_3644 n3_4833_3671 1.714286e-02
R39375 n3_4833_3671 n3_4833_3704 2.095238e-02
R39376 n3_4833_4103 n3_4833_4136 2.095238e-02
R39377 n3_4833_4136 n3_4833_4292 9.904762e-02
R39378 n3_4833_4292 n3_4833_4319 1.714286e-02
R39379 n3_4833_4319 n3_4833_4352 2.095238e-02
R39380 n3_4833_4352 n3_4833_4486 8.507937e-02
R39381 n3_4833_4486 n3_4833_4508 1.396825e-02
R39382 n3_4833_4508 n3_4833_4535 1.714286e-02
R39383 n3_4833_4535 n3_4833_4568 2.095238e-02
R39384 n3_4833_4568 n3_4833_4751 1.161905e-01
R39385 n3_4833_4751 n3_4833_4784 2.095238e-02
R39386 n3_4833_4784 n3_4833_4924 8.888889e-02
R39387 n3_4833_4924 n3_4833_4967 2.730159e-02
R39388 n3_4833_4967 n3_4833_5000 2.095238e-02
R39389 n3_4833_5000 n3_4833_5020 1.269841e-02
R39390 n3_4833_5020 n3_4833_5183 1.034921e-01
R39391 n3_4833_5183 n3_4833_5216 2.095238e-02
R39392 n3_4833_5216 n3_4833_5399 1.161905e-01
R39393 n3_4833_5399 n3_4833_5432 2.095238e-02
R39394 n3_4833_5432 n3_4833_5446 8.888889e-03
R39395 n3_4833_5446 n3_4833_5588 9.015873e-02
R39396 n3_4833_5588 n3_4833_5615 1.714286e-02
R39397 n3_4833_5615 n3_4833_5648 2.095238e-02
R39398 n3_4833_5648 n3_4833_5831 1.161905e-01
R39399 n3_4833_5831 n3_4833_5864 2.095238e-02
R39400 n3_4833_6263 n3_4833_6296 2.095238e-02
R39401 n3_4833_6296 n3_4833_6479 1.161905e-01
R39402 n3_4833_6479 n3_4833_6512 2.095238e-02
R39403 n3_4833_6512 n3_4833_6549 2.349206e-02
R39404 n3_4833_6549 n3_4833_6646 6.158730e-02
R39405 n3_4833_6646 n3_4833_6695 3.111111e-02
R39406 n3_4833_6695 n3_4833_6728 2.095238e-02
R39407 n3_4833_6728 n3_4833_6911 1.161905e-01
R39408 n3_4833_6911 n3_4833_6944 2.095238e-02
R39409 n3_4833_6944 n3_4833_7127 1.161905e-01
R39410 n3_4833_7127 n3_4833_7160 2.095238e-02
R39411 n3_4833_7160 n3_4833_7174 8.888889e-03
R39412 n3_4833_7174 n3_4833_7270 6.095238e-02
R39413 n3_4833_7270 n3_4833_7343 4.634921e-02
R39414 n3_4833_7343 n3_4833_7376 2.095238e-02
R39415 n3_4833_7376 n3_4833_7559 1.161905e-01
R39416 n3_4833_7559 n3_4833_7592 2.095238e-02
R39417 n3_4833_7592 n3_4833_7775 1.161905e-01
R39418 n3_4833_7775 n3_4833_7808 2.095238e-02
R39419 n3_4833_7808 n3_4833_7822 8.888889e-03
R39420 n3_4833_7822 n3_4833_7964 9.015873e-02
R39421 n3_4833_7964 n3_4833_7991 1.714286e-02
R39422 n3_4833_7991 n3_4833_8024 2.095238e-02
R39423 n3_4833_8024 n3_4833_8207 1.161905e-01
R39424 n3_4833_8207 n3_4833_8240 2.095238e-02
R39425 n3_4833_8456 n3_4833_8639 1.161905e-01
R39426 n3_4833_8639 n3_4833_8672 2.095238e-02
R39427 n3_4833_8672 n3_4833_8855 1.161905e-01
R39428 n3_4833_8855 n3_4833_8888 2.095238e-02
R39429 n3_4833_8888 n3_4833_8902 8.888889e-03
R39430 n3_4833_8902 n3_4833_9022 7.619048e-02
R39431 n3_4833_9022 n3_4833_9044 1.396825e-02
R39432 n3_4833_9044 n3_4833_9071 1.714286e-02
R39433 n3_4833_9071 n3_4833_9104 2.095238e-02
R39434 n3_4833_9104 n3_4833_9287 1.161905e-01
R39435 n3_4833_9287 n3_4833_9320 2.095238e-02
R39436 n3_4833_9320 n3_4833_9424 6.603175e-02
R39437 n3_4833_9424 n3_4833_9503 5.015873e-02
R39438 n3_4833_9503 n3_4833_9520 1.079365e-02
R39439 n3_4833_9520 n3_4833_9536 1.015873e-02
R39440 n3_4833_9536 n3_4833_9719 1.161905e-01
R39441 n3_4833_9719 n3_4833_9752 2.095238e-02
R39442 n3_4833_9752 n3_4833_9935 1.161905e-01
R39443 n3_4833_9935 n3_4833_9968 2.095238e-02
R39444 n3_4833_9968 n3_4833_9982 8.888889e-03
R39445 n3_4833_9982 n3_4833_10124 9.015873e-02
R39446 n3_4833_10124 n3_4833_10151 1.714286e-02
R39447 n3_4833_10151 n3_4833_10184 2.095238e-02
R39448 n3_4833_10184 n3_4833_10367 1.161905e-01
R39449 n3_4833_10367 n3_4833_10400 2.095238e-02
R39450 n3_4833_10799 n3_4833_10832 2.095238e-02
R39451 n3_4833_10832 n3_4833_11015 1.161905e-01
R39452 n3_4833_11015 n3_4833_11048 2.095238e-02
R39453 n3_4833_11048 n3_4833_11182 8.507937e-02
R39454 n3_4833_11182 n3_4833_11204 1.396825e-02
R39455 n3_4833_11204 n3_4833_11231 1.714286e-02
R39456 n3_4833_11231 n3_4833_11264 2.095238e-02
R39457 n3_4833_11264 n3_4833_11447 1.161905e-01
R39458 n3_4833_11447 n3_4833_11480 2.095238e-02
R39459 n3_4833_11480 n3_4833_11663 1.161905e-01
R39460 n3_4833_11663 n3_4833_11674 6.984127e-03
R39461 n3_4833_11674 n3_4833_11696 1.396825e-02
R39462 n3_4833_11696 n3_4833_11770 4.698413e-02
R39463 n3_4833_11770 n3_4833_11879 6.920635e-02
R39464 n3_4833_11879 n3_4833_11912 2.095238e-02
R39465 n3_4833_11912 n3_4833_12095 1.161905e-01
R39466 n3_4833_12095 n3_4833_12128 2.095238e-02
R39467 n3_4833_12128 n3_4833_12284 9.904762e-02
R39468 n3_4833_12284 n3_4833_12311 1.714286e-02
R39469 n3_4833_12311 n3_4833_12344 2.095238e-02
R39470 n3_4833_12344 n3_4833_12527 1.161905e-01
R39471 n3_4833_12527 n3_4833_12560 2.095238e-02
R39472 n3_4833_12560 n3_4833_12743 1.161905e-01
R39473 n3_4833_12959 n3_4833_12992 2.095238e-02
R39474 n3_4833_12992 n3_4833_13175 1.161905e-01
R39475 n3_4833_13175 n3_4833_13208 2.095238e-02
R39476 n3_4833_13208 n3_4833_13391 1.161905e-01
R39477 n3_4833_13391 n3_4833_13424 2.095238e-02
R39478 n3_4833_13424 n3_4833_13580 9.904762e-02
R39479 n3_4833_13580 n3_4833_13607 1.714286e-02
R39480 n3_4833_13607 n3_4833_13640 2.095238e-02
R39481 n3_4833_13640 n3_4833_13823 1.161905e-01
R39482 n3_4833_13823 n3_4833_13856 2.095238e-02
R39483 n3_4833_13856 n3_4833_13924 4.317460e-02
R39484 n3_4833_13924 n3_4833_13990 4.190476e-02
R39485 n3_4833_13990 n3_4833_14020 1.904762e-02
R39486 n3_4833_14020 n3_4833_14039 1.206349e-02
R39487 n3_4833_14039 n3_4833_14072 2.095238e-02
R39488 n3_4833_14072 n3_4833_14206 8.507937e-02
R39489 n3_4833_14206 n3_4833_14255 3.111111e-02
R39490 n3_4833_14255 n3_4833_14288 2.095238e-02
R39491 n3_4833_14288 n3_4833_14471 1.161905e-01
R39492 n3_4833_14471 n3_4833_14504 2.095238e-02
R39493 n3_4833_14504 n3_4833_14687 1.161905e-01
R39494 n3_4833_14687 n3_4833_14720 2.095238e-02
R39495 n3_4833_14720 n3_4833_14903 1.161905e-01
R39496 n3_4833_14903 n3_4833_14936 2.095238e-02
R39497 n3_4833_15335 n3_4833_15368 2.095238e-02
R39498 n3_4833_15368 n3_4833_15524 9.904762e-02
R39499 n3_4833_15524 n3_4833_15551 1.714286e-02
R39500 n3_4833_15551 n3_4833_15584 2.095238e-02
R39501 n3_4833_15584 n3_4833_15740 9.904762e-02
R39502 n3_4833_15740 n3_4833_15767 1.714286e-02
R39503 n3_4833_15767 n3_4833_15800 2.095238e-02
R39504 n3_4833_15800 n3_4833_15983 1.161905e-01
R39505 n3_4833_15983 n3_4833_16016 2.095238e-02
R39506 n3_4833_16016 n3_4833_16172 9.904762e-02
R39507 n3_4833_16172 n3_4833_16174 1.269841e-03
R39508 n3_4833_16174 n3_4833_16199 1.587302e-02
R39509 n3_4833_16199 n3_4833_16232 2.095238e-02
R39510 n3_4833_16232 n3_4833_16270 2.412698e-02
R39511 n3_4833_16270 n3_4833_16415 9.206349e-02
R39512 n3_4833_16415 n3_4833_16448 2.095238e-02
R39513 n3_4833_16448 n3_4833_16631 1.161905e-01
R39514 n3_4833_16631 n3_4833_16664 2.095238e-02
R39515 n3_4833_16664 n3_4833_16847 1.161905e-01
R39516 n3_4833_16847 n3_4833_16880 2.095238e-02
R39517 n3_4833_16880 n3_4833_17036 9.904762e-02
R39518 n3_4833_17036 n3_4833_17063 1.714286e-02
R39519 n3_4833_17063 n3_4833_17096 2.095238e-02
R39520 n3_4833_17468 n3_4833_17495 1.714286e-02
R39521 n3_4833_17495 n3_4833_17528 2.095238e-02
R39522 n3_4833_17528 n3_4833_17684 9.904762e-02
R39523 n3_4833_17684 n3_4833_17711 1.714286e-02
R39524 n3_4833_17711 n3_4833_17744 2.095238e-02
R39525 n3_4833_17744 n3_4833_17927 1.161905e-01
R39526 n3_4833_17927 n3_4833_17960 2.095238e-02
R39527 n3_4833_17960 n3_4833_18143 1.161905e-01
R39528 n3_4833_18143 n3_4833_18176 2.095238e-02
R39529 n3_4833_18176 n3_4833_18359 1.161905e-01
R39530 n3_4833_18359 n3_4833_18392 2.095238e-02
R39531 n3_4833_18392 n3_4833_18424 2.031746e-02
R39532 n3_4833_18424 n3_4833_18520 6.095238e-02
R39533 n3_4833_18520 n3_4833_18527 4.444444e-03
R39534 n3_4833_18527 n3_4833_18548 1.333333e-02
R39535 n3_4833_18548 n3_4833_18575 1.714286e-02
R39536 n3_4833_18575 n3_4833_18608 2.095238e-02
R39537 n3_4833_18608 n3_4833_18764 9.904762e-02
R39538 n3_4833_18764 n3_4833_18791 1.714286e-02
R39539 n3_4833_18791 n3_4833_18824 2.095238e-02
R39540 n3_4833_18824 n3_4833_18980 9.904762e-02
R39541 n3_4833_18980 n3_4833_19007 1.714286e-02
R39542 n3_4833_19007 n3_4833_19040 2.095238e-02
R39543 n3_4833_19040 n3_4833_19196 9.904762e-02
R39544 n3_4833_19196 n3_4833_19223 1.714286e-02
R39545 n3_4833_19223 n3_4833_19256 2.095238e-02
R39546 n3_4833_19256 n3_4833_19439 1.161905e-01
R39547 n3_4833_19439 n3_4833_19472 2.095238e-02
R39548 n3_4833_19871 n3_4833_19904 2.095238e-02
R39549 n3_4833_19904 n3_4833_20087 1.161905e-01
R39550 n3_4833_20087 n3_4833_20120 2.095238e-02
R39551 n3_4833_20120 n3_4833_20303 1.161905e-01
R39552 n3_4833_20303 n3_4833_20336 2.095238e-02
R39553 n3_4833_20336 n3_4833_20519 1.161905e-01
R39554 n3_4833_20519 n3_4833_20552 2.095238e-02
R39555 n3_4833_20552 n3_4833_20674 7.746032e-02
R39556 n3_4833_20674 n3_4833_20687 8.253968e-03
R39557 n3_4833_20687 n3_4833_20735 3.047619e-02
R39558 n3_4833_20735 n3_4833_20768 2.095238e-02
R39559 n3_4833_20768 n3_4833_20770 1.269841e-03
R39560 n3_4833_20770 n3_4833_20951 1.149206e-01
R39561 n3_4833_20951 n3_4833_20984 2.095238e-02
R39562 n3_5021_215 n3_5021_248 2.095238e-02
R39563 n3_5021_248 n3_5021_424 1.117460e-01
R39564 n3_5021_424 n3_5021_431 4.444444e-03
R39565 n3_5021_513 n3_5021_520 4.444444e-03
R39566 n3_5021_520 n3_5021_647 8.063492e-02
R39567 n3_5021_647 n3_5021_680 2.095238e-02
R39568 n3_5021_680 n3_5021_863 1.161905e-01
R39569 n3_5021_863 n3_5021_896 2.095238e-02
R39570 n3_5021_896 n3_5021_945 3.111111e-02
R39571 n3_5021_945 n3_5021_1079 8.507937e-02
R39572 n3_5021_1079 n3_5021_1112 2.095238e-02
R39573 n3_5021_1112 n3_5021_1295 1.161905e-01
R39574 n3_5021_1295 n3_5021_1328 2.095238e-02
R39575 n3_5021_1328 n3_5021_1511 1.161905e-01
R39576 n3_5021_1511 n3_5021_1544 2.095238e-02
R39577 n3_5021_1544 n3_5021_1727 1.161905e-01
R39578 n3_5021_1727 n3_5021_1760 2.095238e-02
R39579 n3_5021_1760 n3_5021_1916 9.904762e-02
R39580 n3_5021_1916 n3_5021_1943 1.714286e-02
R39581 n3_5021_1943 n3_5021_1976 2.095238e-02
R39582 n3_5021_1976 n3_5021_2132 9.904762e-02
R39583 n3_5021_2132 n3_5021_2159 1.714286e-02
R39584 n3_5021_2159 n3_5021_2192 2.095238e-02
R39585 n3_5021_2192 n3_5021_2375 1.161905e-01
R39586 n3_5021_2375 n3_5021_2408 2.095238e-02
R39587 n3_5021_2408 n3_5021_2543 8.571429e-02
R39588 n3_5021_2543 n3_5021_2564 1.333333e-02
R39589 n3_5021_2564 n3_5021_2591 1.714286e-02
R39590 n3_5021_2591 n3_5021_2624 2.095238e-02
R39591 n3_5021_2624 n3_5021_2674 3.174603e-02
R39592 n3_5021_2770 n3_5021_2807 2.349206e-02
R39593 n3_5021_2807 n3_5021_2840 2.095238e-02
R39594 n3_5021_2840 n3_5021_2996 9.904762e-02
R39595 n3_5021_2996 n3_5021_3023 1.714286e-02
R39596 n3_5021_3023 n3_5021_3056 2.095238e-02
R39597 n3_5021_3056 n3_5021_3212 9.904762e-02
R39598 n3_5021_3212 n3_5021_3239 1.714286e-02
R39599 n3_5021_3239 n3_5021_3272 2.095238e-02
R39600 n3_5021_3272 n3_5021_3455 1.161905e-01
R39601 n3_5021_3455 n3_5021_3488 2.095238e-02
R39602 n3_5021_3488 n3_5021_3644 9.904762e-02
R39603 n3_5021_3644 n3_5021_3671 1.714286e-02
R39604 n3_5021_3671 n3_5021_3704 2.095238e-02
R39605 n3_5021_3704 n3_5021_3887 1.161905e-01
R39606 n3_5021_3887 n3_5021_3920 2.095238e-02
R39607 n3_5021_3920 n3_5021_4103 1.161905e-01
R39608 n3_5021_4103 n3_5021_4136 2.095238e-02
R39609 n3_5021_4136 n3_5021_4292 9.904762e-02
R39610 n3_5021_4292 n3_5021_4319 1.714286e-02
R39611 n3_5021_4319 n3_5021_4352 2.095238e-02
R39612 n3_5021_4352 n3_5021_4486 8.507937e-02
R39613 n3_5021_4486 n3_5021_4508 1.396825e-02
R39614 n3_5021_4508 n3_5021_4535 1.714286e-02
R39615 n3_5021_4535 n3_5021_4568 2.095238e-02
R39616 n3_5021_4568 n3_5021_4751 1.161905e-01
R39617 n3_5021_4751 n3_5021_4784 2.095238e-02
R39618 n3_5021_4784 n3_5021_4924 8.888889e-02
R39619 n3_5021_5000 n3_5021_5020 1.269841e-02
R39620 n3_5021_5020 n3_5021_5183 1.034921e-01
R39621 n3_5021_5183 n3_5021_5216 2.095238e-02
R39622 n3_5021_5216 n3_5021_5399 1.161905e-01
R39623 n3_5021_5399 n3_5021_5432 2.095238e-02
R39624 n3_5021_5432 n3_5021_5446 8.888889e-03
R39625 n3_5021_5446 n3_5021_5588 9.015873e-02
R39626 n3_5021_5588 n3_5021_5615 1.714286e-02
R39627 n3_5021_5615 n3_5021_5648 2.095238e-02
R39628 n3_5021_5648 n3_5021_5831 1.161905e-01
R39629 n3_5021_5831 n3_5021_5864 2.095238e-02
R39630 n3_5021_5864 n3_5021_6047 1.161905e-01
R39631 n3_5021_6047 n3_5021_6080 2.095238e-02
R39632 n3_5021_6080 n3_5021_6263 1.161905e-01
R39633 n3_5021_6263 n3_5021_6296 2.095238e-02
R39634 n3_5021_6296 n3_5021_6479 1.161905e-01
R39635 n3_5021_6479 n3_5021_6512 2.095238e-02
R39636 n3_5021_6512 n3_5021_6549 2.349206e-02
R39637 n3_5021_6549 n3_5021_6646 6.158730e-02
R39638 n3_5021_6646 n3_5021_6695 3.111111e-02
R39639 n3_5021_6695 n3_5021_6728 2.095238e-02
R39640 n3_5021_6728 n3_5021_6911 1.161905e-01
R39641 n3_5021_6911 n3_5021_6944 2.095238e-02
R39642 n3_5021_6944 n3_5021_7127 1.161905e-01
R39643 n3_5021_7127 n3_5021_7160 2.095238e-02
R39644 n3_5021_7160 n3_5021_7174 8.888889e-03
R39645 n3_5021_7270 n3_5021_7343 4.634921e-02
R39646 n3_5021_7343 n3_5021_7376 2.095238e-02
R39647 n3_5021_7376 n3_5021_7559 1.161905e-01
R39648 n3_5021_7559 n3_5021_7592 2.095238e-02
R39649 n3_5021_7592 n3_5021_7775 1.161905e-01
R39650 n3_5021_7775 n3_5021_7808 2.095238e-02
R39651 n3_5021_7808 n3_5021_7822 8.888889e-03
R39652 n3_5021_7822 n3_5021_7964 9.015873e-02
R39653 n3_5021_7964 n3_5021_7991 1.714286e-02
R39654 n3_5021_7991 n3_5021_8024 2.095238e-02
R39655 n3_5021_8024 n3_5021_8207 1.161905e-01
R39656 n3_5021_8207 n3_5021_8240 2.095238e-02
R39657 n3_5021_8240 n3_5021_8423 1.161905e-01
R39658 n3_5021_8423 n3_5021_8456 2.095238e-02
R39659 n3_5021_8456 n3_5021_8639 1.161905e-01
R39660 n3_5021_8639 n3_5021_8672 2.095238e-02
R39661 n3_5021_8672 n3_5021_8855 1.161905e-01
R39662 n3_5021_8855 n3_5021_8888 2.095238e-02
R39663 n3_5021_8888 n3_5021_8902 8.888889e-03
R39664 n3_5021_8902 n3_5021_9022 7.619048e-02
R39665 n3_5021_9022 n3_5021_9044 1.396825e-02
R39666 n3_5021_9044 n3_5021_9071 1.714286e-02
R39667 n3_5021_9071 n3_5021_9104 2.095238e-02
R39668 n3_5021_9104 n3_5021_9287 1.161905e-01
R39669 n3_5021_9287 n3_5021_9320 2.095238e-02
R39670 n3_5021_9320 n3_5021_9424 6.603175e-02
R39671 n3_5021_9503 n3_5021_9520 1.079365e-02
R39672 n3_5021_9520 n3_5021_9536 1.015873e-02
R39673 n3_5021_9536 n3_5021_9719 1.161905e-01
R39674 n3_5021_9719 n3_5021_9752 2.095238e-02
R39675 n3_5021_9752 n3_5021_9935 1.161905e-01
R39676 n3_5021_9935 n3_5021_9968 2.095238e-02
R39677 n3_5021_9968 n3_5021_9982 8.888889e-03
R39678 n3_5021_9982 n3_5021_10124 9.015873e-02
R39679 n3_5021_10124 n3_5021_10151 1.714286e-02
R39680 n3_5021_10151 n3_5021_10184 2.095238e-02
R39681 n3_5021_10184 n3_5021_10367 1.161905e-01
R39682 n3_5021_10367 n3_5021_10400 2.095238e-02
R39683 n3_5021_10616 n3_5021_10799 1.161905e-01
R39684 n3_5021_10799 n3_5021_10832 2.095238e-02
R39685 n3_5021_10832 n3_5021_11015 1.161905e-01
R39686 n3_5021_11015 n3_5021_11048 2.095238e-02
R39687 n3_5021_11048 n3_5021_11182 8.507937e-02
R39688 n3_5021_11182 n3_5021_11204 1.396825e-02
R39689 n3_5021_11204 n3_5021_11231 1.714286e-02
R39690 n3_5021_11231 n3_5021_11264 2.095238e-02
R39691 n3_5021_11264 n3_5021_11447 1.161905e-01
R39692 n3_5021_11447 n3_5021_11480 2.095238e-02
R39693 n3_5021_11480 n3_5021_11663 1.161905e-01
R39694 n3_5021_11663 n3_5021_11674 6.984127e-03
R39695 n3_5021_11674 n3_5021_11696 1.396825e-02
R39696 n3_5021_11770 n3_5021_11879 6.920635e-02
R39697 n3_5021_11879 n3_5021_11912 2.095238e-02
R39698 n3_5021_11912 n3_5021_12095 1.161905e-01
R39699 n3_5021_12095 n3_5021_12128 2.095238e-02
R39700 n3_5021_12128 n3_5021_12284 9.904762e-02
R39701 n3_5021_12284 n3_5021_12311 1.714286e-02
R39702 n3_5021_12311 n3_5021_12344 2.095238e-02
R39703 n3_5021_12344 n3_5021_12527 1.161905e-01
R39704 n3_5021_12527 n3_5021_12560 2.095238e-02
R39705 n3_5021_12560 n3_5021_12743 1.161905e-01
R39706 n3_5021_12743 n3_5021_12776 2.095238e-02
R39707 n3_5021_12776 n3_5021_12959 1.161905e-01
R39708 n3_5021_12959 n3_5021_12992 2.095238e-02
R39709 n3_5021_12992 n3_5021_13175 1.161905e-01
R39710 n3_5021_13175 n3_5021_13208 2.095238e-02
R39711 n3_5021_13208 n3_5021_13391 1.161905e-01
R39712 n3_5021_13391 n3_5021_13424 2.095238e-02
R39713 n3_5021_13424 n3_5021_13580 9.904762e-02
R39714 n3_5021_13580 n3_5021_13607 1.714286e-02
R39715 n3_5021_13607 n3_5021_13640 2.095238e-02
R39716 n3_5021_13640 n3_5021_13823 1.161905e-01
R39717 n3_5021_13823 n3_5021_13856 2.095238e-02
R39718 n3_5021_13856 n3_5021_13924 4.317460e-02
R39719 n3_5021_14020 n3_5021_14039 1.206349e-02
R39720 n3_5021_14039 n3_5021_14072 2.095238e-02
R39721 n3_5021_14072 n3_5021_14206 8.507937e-02
R39722 n3_5021_14206 n3_5021_14255 3.111111e-02
R39723 n3_5021_14255 n3_5021_14288 2.095238e-02
R39724 n3_5021_14288 n3_5021_14471 1.161905e-01
R39725 n3_5021_14471 n3_5021_14504 2.095238e-02
R39726 n3_5021_14504 n3_5021_14687 1.161905e-01
R39727 n3_5021_14687 n3_5021_14720 2.095238e-02
R39728 n3_5021_14720 n3_5021_14903 1.161905e-01
R39729 n3_5021_14903 n3_5021_14936 2.095238e-02
R39730 n3_5021_14936 n3_5021_15119 1.161905e-01
R39731 n3_5021_15119 n3_5021_15152 2.095238e-02
R39732 n3_5021_15152 n3_5021_15335 1.161905e-01
R39733 n3_5021_15335 n3_5021_15368 2.095238e-02
R39734 n3_5021_15368 n3_5021_15524 9.904762e-02
R39735 n3_5021_15524 n3_5021_15551 1.714286e-02
R39736 n3_5021_15551 n3_5021_15584 2.095238e-02
R39737 n3_5021_15584 n3_5021_15740 9.904762e-02
R39738 n3_5021_15740 n3_5021_15767 1.714286e-02
R39739 n3_5021_15767 n3_5021_15800 2.095238e-02
R39740 n3_5021_15800 n3_5021_15983 1.161905e-01
R39741 n3_5021_15983 n3_5021_16016 2.095238e-02
R39742 n3_5021_16016 n3_5021_16172 9.904762e-02
R39743 n3_5021_16172 n3_5021_16174 1.269841e-03
R39744 n3_5021_16174 n3_5021_16199 1.587302e-02
R39745 n3_5021_16270 n3_5021_16415 9.206349e-02
R39746 n3_5021_16415 n3_5021_16448 2.095238e-02
R39747 n3_5021_16448 n3_5021_16631 1.161905e-01
R39748 n3_5021_16631 n3_5021_16664 2.095238e-02
R39749 n3_5021_16664 n3_5021_16847 1.161905e-01
R39750 n3_5021_16847 n3_5021_16880 2.095238e-02
R39751 n3_5021_16880 n3_5021_17036 9.904762e-02
R39752 n3_5021_17036 n3_5021_17063 1.714286e-02
R39753 n3_5021_17063 n3_5021_17096 2.095238e-02
R39754 n3_5021_17096 n3_5021_17252 9.904762e-02
R39755 n3_5021_17252 n3_5021_17279 1.714286e-02
R39756 n3_5021_17279 n3_5021_17312 2.095238e-02
R39757 n3_5021_17312 n3_5021_17446 8.507937e-02
R39758 n3_5021_17446 n3_5021_17468 1.396825e-02
R39759 n3_5021_17468 n3_5021_17495 1.714286e-02
R39760 n3_5021_17495 n3_5021_17528 2.095238e-02
R39761 n3_5021_17528 n3_5021_17684 9.904762e-02
R39762 n3_5021_17684 n3_5021_17711 1.714286e-02
R39763 n3_5021_17711 n3_5021_17744 2.095238e-02
R39764 n3_5021_17744 n3_5021_17927 1.161905e-01
R39765 n3_5021_17927 n3_5021_17960 2.095238e-02
R39766 n3_5021_17960 n3_5021_18143 1.161905e-01
R39767 n3_5021_18143 n3_5021_18176 2.095238e-02
R39768 n3_5021_18176 n3_5021_18359 1.161905e-01
R39769 n3_5021_18359 n3_5021_18392 2.095238e-02
R39770 n3_5021_18392 n3_5021_18424 2.031746e-02
R39771 n3_5021_18520 n3_5021_18527 4.444444e-03
R39772 n3_5021_18527 n3_5021_18548 1.333333e-02
R39773 n3_5021_18548 n3_5021_18575 1.714286e-02
R39774 n3_5021_18575 n3_5021_18608 2.095238e-02
R39775 n3_5021_18608 n3_5021_18764 9.904762e-02
R39776 n3_5021_18764 n3_5021_18791 1.714286e-02
R39777 n3_5021_18791 n3_5021_18824 2.095238e-02
R39778 n3_5021_18824 n3_5021_18980 9.904762e-02
R39779 n3_5021_18980 n3_5021_19007 1.714286e-02
R39780 n3_5021_19007 n3_5021_19040 2.095238e-02
R39781 n3_5021_19040 n3_5021_19196 9.904762e-02
R39782 n3_5021_19196 n3_5021_19223 1.714286e-02
R39783 n3_5021_19223 n3_5021_19256 2.095238e-02
R39784 n3_5021_19256 n3_5021_19439 1.161905e-01
R39785 n3_5021_19439 n3_5021_19472 2.095238e-02
R39786 n3_5021_19472 n3_5021_19628 9.904762e-02
R39787 n3_5021_19628 n3_5021_19655 1.714286e-02
R39788 n3_5021_19655 n3_5021_19688 2.095238e-02
R39789 n3_5021_19688 n3_5021_19871 1.161905e-01
R39790 n3_5021_19871 n3_5021_19904 2.095238e-02
R39791 n3_5021_19904 n3_5021_20087 1.161905e-01
R39792 n3_5021_20087 n3_5021_20120 2.095238e-02
R39793 n3_5021_20120 n3_5021_20303 1.161905e-01
R39794 n3_5021_20303 n3_5021_20336 2.095238e-02
R39795 n3_5021_20336 n3_5021_20519 1.161905e-01
R39796 n3_5021_20519 n3_5021_20552 2.095238e-02
R39797 n3_5021_20552 n3_5021_20674 7.746032e-02
R39798 n3_5021_20674 n3_5021_20687 8.253968e-03
R39799 n3_5021_20768 n3_5021_20770 1.269841e-03
R39800 n3_5021_20770 n3_5021_20951 1.149206e-01
R39801 n3_5021_20951 n3_5021_20984 2.095238e-02
R39802 n3_5114_215 n3_5114_248 2.095238e-02
R39803 n3_5114_248 n3_5114_431 1.161905e-01
R39804 n3_5114_431 n3_5114_464 2.095238e-02
R39805 n3_5114_464 n3_5114_513 3.111111e-02
R39806 n3_5114_513 n3_5114_647 8.507937e-02
R39807 n3_5114_647 n3_5114_680 2.095238e-02
R39808 n3_5114_680 n3_5114_863 1.161905e-01
R39809 n3_5114_863 n3_5114_896 2.095238e-02
R39810 n3_5114_896 n3_5114_945 3.111111e-02
R39811 n3_5114_945 n3_5114_1079 8.507937e-02
R39812 n3_5114_1079 n3_5114_1112 2.095238e-02
R39813 n3_5114_1112 n3_5114_1295 1.161905e-01
R39814 n3_5114_1295 n3_5114_1328 2.095238e-02
R39815 n3_5114_1328 n3_5114_1511 1.161905e-01
R39816 n3_5114_1511 n3_5114_1544 2.095238e-02
R39817 n3_5114_1544 n3_5114_1727 1.161905e-01
R39818 n3_5114_1727 n3_5114_1760 2.095238e-02
R39819 n3_5114_1760 n3_5114_1916 9.904762e-02
R39820 n3_5114_1916 n3_5114_1943 1.714286e-02
R39821 n3_5114_1943 n3_5114_1976 2.095238e-02
R39822 n3_5114_1976 n3_5114_2159 1.161905e-01
R39823 n3_5114_2159 n3_5114_2192 2.095238e-02
R39824 n3_5114_2192 n3_5114_2375 1.161905e-01
R39825 n3_5114_2375 n3_5114_2408 2.095238e-02
R39826 n3_5114_2408 n3_5114_2543 8.571429e-02
R39827 n3_5114_2543 n3_5114_2564 1.333333e-02
R39828 n3_5114_2564 n3_5114_2591 1.714286e-02
R39829 n3_5114_2591 n3_5114_2624 2.095238e-02
R39830 n3_5114_18527 n3_5114_18548 1.333333e-02
R39831 n3_5114_18548 n3_5114_18575 1.714286e-02
R39832 n3_5114_18575 n3_5114_18608 2.095238e-02
R39833 n3_5114_18608 n3_5114_18764 9.904762e-02
R39834 n3_5114_18764 n3_5114_18791 1.714286e-02
R39835 n3_5114_18791 n3_5114_18824 2.095238e-02
R39836 n3_5114_18824 n3_5114_18980 9.904762e-02
R39837 n3_5114_18980 n3_5114_19007 1.714286e-02
R39838 n3_5114_19007 n3_5114_19040 2.095238e-02
R39839 n3_5114_19040 n3_5114_19196 9.904762e-02
R39840 n3_5114_19196 n3_5114_19223 1.714286e-02
R39841 n3_5114_19223 n3_5114_19256 2.095238e-02
R39842 n3_5114_19256 n3_5114_19439 1.161905e-01
R39843 n3_5114_19439 n3_5114_19472 2.095238e-02
R39844 n3_5114_19472 n3_5114_19628 9.904762e-02
R39845 n3_5114_19628 n3_5114_19655 1.714286e-02
R39846 n3_5114_19655 n3_5114_19688 2.095238e-02
R39847 n3_5114_19688 n3_5114_19871 1.161905e-01
R39848 n3_5114_19871 n3_5114_19904 2.095238e-02
R39849 n3_5114_19904 n3_5114_20087 1.161905e-01
R39850 n3_5114_20087 n3_5114_20120 2.095238e-02
R39851 n3_5114_20120 n3_5114_20303 1.161905e-01
R39852 n3_5114_20303 n3_5114_20336 2.095238e-02
R39853 n3_5114_20336 n3_5114_20519 1.161905e-01
R39854 n3_5114_20519 n3_5114_20552 2.095238e-02
R39855 n3_5114_20552 n3_5114_20687 8.571429e-02
R39856 n3_5114_20687 n3_5114_20735 3.047619e-02
R39857 n3_5114_20735 n3_5114_20768 2.095238e-02
R39858 n3_5114_20768 n3_5114_20951 1.161905e-01
R39859 n3_5114_20951 n3_5114_20984 2.095238e-02
R39860 n3_6900_215 n3_6900_248 2.095238e-02
R39861 n3_6900_248 n3_6900_383 8.571429e-02
R39862 n3_6900_383 n3_6900_431 3.047619e-02
R39863 n3_6900_431 n3_6900_464 2.095238e-02
R39864 n3_6900_464 n3_6900_647 1.161905e-01
R39865 n3_6900_647 n3_6900_680 2.095238e-02
R39866 n3_6900_680 n3_6900_863 1.161905e-01
R39867 n3_6900_863 n3_6900_896 2.095238e-02
R39868 n3_6900_896 n3_6900_1079 1.161905e-01
R39869 n3_6900_1079 n3_6900_1112 2.095238e-02
R39870 n3_6900_1112 n3_6900_1295 1.161905e-01
R39871 n3_6900_1295 n3_6900_1328 2.095238e-02
R39872 n3_6900_1328 n3_6900_1511 1.161905e-01
R39873 n3_6900_1511 n3_6900_1544 2.095238e-02
R39874 n3_6900_1544 n3_6900_1727 1.161905e-01
R39875 n3_6900_1727 n3_6900_1760 2.095238e-02
R39876 n3_6900_1760 n3_6900_1916 9.904762e-02
R39877 n3_6900_1916 n3_6900_1943 1.714286e-02
R39878 n3_6900_1943 n3_6900_1976 2.095238e-02
R39879 n3_6900_1976 n3_6900_2159 1.161905e-01
R39880 n3_6900_2159 n3_6900_2192 2.095238e-02
R39881 n3_6900_2192 n3_6900_2375 1.161905e-01
R39882 n3_6900_2375 n3_6900_2408 2.095238e-02
R39883 n3_6900_2408 n3_6900_2543 8.571429e-02
R39884 n3_6900_2543 n3_6900_2564 1.333333e-02
R39885 n3_6900_2564 n3_6900_2591 1.714286e-02
R39886 n3_6900_2591 n3_6900_2624 2.095238e-02
R39887 n3_6900_18527 n3_6900_18548 1.333333e-02
R39888 n3_6900_18548 n3_6900_18575 1.714286e-02
R39889 n3_6900_18575 n3_6900_18608 2.095238e-02
R39890 n3_6900_18608 n3_6900_18764 9.904762e-02
R39891 n3_6900_18764 n3_6900_18791 1.714286e-02
R39892 n3_6900_18791 n3_6900_18824 2.095238e-02
R39893 n3_6900_18824 n3_6900_19007 1.161905e-01
R39894 n3_6900_19007 n3_6900_19040 2.095238e-02
R39895 n3_6900_19040 n3_6900_19196 9.904762e-02
R39896 n3_6900_19196 n3_6900_19223 1.714286e-02
R39897 n3_6900_19223 n3_6900_19256 2.095238e-02
R39898 n3_6900_19256 n3_6900_19439 1.161905e-01
R39899 n3_6900_19439 n3_6900_19472 2.095238e-02
R39900 n3_6900_19472 n3_6900_19655 1.161905e-01
R39901 n3_6900_19655 n3_6900_19688 2.095238e-02
R39902 n3_6900_19688 n3_6900_19871 1.161905e-01
R39903 n3_6900_19871 n3_6900_19904 2.095238e-02
R39904 n3_6900_19904 n3_6900_20087 1.161905e-01
R39905 n3_6900_20087 n3_6900_20120 2.095238e-02
R39906 n3_6900_20120 n3_6900_20303 1.161905e-01
R39907 n3_6900_20303 n3_6900_20336 2.095238e-02
R39908 n3_6900_20336 n3_6900_20519 1.161905e-01
R39909 n3_6900_20519 n3_6900_20552 2.095238e-02
R39910 n3_6900_20552 n3_6900_20687 8.571429e-02
R39911 n3_6900_20687 n3_6900_20735 3.047619e-02
R39912 n3_6900_20735 n3_6900_20768 2.095238e-02
R39913 n3_6900_20768 n3_6900_20951 1.161905e-01
R39914 n3_6900_20951 n3_6900_20984 2.095238e-02
R39915 n3_7083_424 n3_7130_424 2.984127e-02
R39916 n3_7130_424 n3_7271_424 8.952381e-02
R39917 n3_7083_520 n3_7130_520 2.984127e-02
R39918 n3_7130_520 n3_7271_520 8.952381e-02
R39919 n3_7083_2674 n3_7130_2674 2.984127e-02
R39920 n3_7130_2674 n3_7271_2674 8.952381e-02
R39921 n3_7083_2770 n3_7130_2770 2.984127e-02
R39922 n3_7130_2770 n3_7271_2770 8.952381e-02
R39923 n3_7083_4924 n3_7130_4924 2.984127e-02
R39924 n3_7130_4924 n3_7271_4924 8.952381e-02
R39925 n3_7083_5020 n3_7130_5020 2.984127e-02
R39926 n3_7130_5020 n3_7271_5020 8.952381e-02
R39927 n3_7083_7174 n3_7130_7174 2.984127e-02
R39928 n3_7130_7174 n3_7271_7174 8.952381e-02
R39929 n3_7083_7270 n3_7130_7270 2.984127e-02
R39930 n3_7130_7270 n3_7271_7270 8.952381e-02
R39931 n3_7083_9424 n3_7130_9424 2.984127e-02
R39932 n3_7130_9424 n3_7271_9424 8.952381e-02
R39933 n3_7083_9520 n3_7130_9520 2.984127e-02
R39934 n3_7130_9520 n3_7271_9520 8.952381e-02
R39935 n3_7083_11674 n3_7130_11674 2.984127e-02
R39936 n3_7130_11674 n3_7271_11674 8.952381e-02
R39937 n3_7083_11770 n3_7130_11770 2.984127e-02
R39938 n3_7130_11770 n3_7271_11770 8.952381e-02
R39939 n3_7083_13924 n3_7130_13924 2.984127e-02
R39940 n3_7130_13924 n3_7271_13924 8.952381e-02
R39941 n3_7083_14020 n3_7130_14020 2.984127e-02
R39942 n3_7130_14020 n3_7271_14020 8.952381e-02
R39943 n3_7083_16174 n3_7130_16174 2.984127e-02
R39944 n3_7130_16174 n3_7271_16174 8.952381e-02
R39945 n3_7083_16270 n3_7130_16270 2.984127e-02
R39946 n3_7130_16270 n3_7271_16270 8.952381e-02
R39947 n3_7083_18424 n3_7130_18424 2.984127e-02
R39948 n3_7130_18424 n3_7271_18424 8.952381e-02
R39949 n3_7083_18520 n3_7130_18520 2.984127e-02
R39950 n3_7130_18520 n3_7271_18520 8.952381e-02
R39951 n3_7083_20674 n3_7130_20674 2.984127e-02
R39952 n3_7130_20674 n3_7271_20674 8.952381e-02
R39953 n3_7083_20770 n3_7130_20770 2.984127e-02
R39954 n3_7130_20770 n3_7271_20770 8.952381e-02
R39955 n3_7083_215 n3_7083_248 2.095238e-02
R39956 n3_7083_248 n3_7083_383 8.571429e-02
R39957 n3_7083_383 n3_7083_424 2.603175e-02
R39958 n3_7083_424 n3_7083_431 4.444444e-03
R39959 n3_7083_431 n3_7083_464 2.095238e-02
R39960 n3_7083_464 n3_7083_520 3.555556e-02
R39961 n3_7083_520 n3_7083_647 8.063492e-02
R39962 n3_7083_647 n3_7083_680 2.095238e-02
R39963 n3_7083_680 n3_7083_863 1.161905e-01
R39964 n3_7083_863 n3_7083_896 2.095238e-02
R39965 n3_7083_896 n3_7083_1079 1.161905e-01
R39966 n3_7083_1079 n3_7083_1112 2.095238e-02
R39967 n3_7083_1112 n3_7083_1295 1.161905e-01
R39968 n3_7083_1295 n3_7083_1328 2.095238e-02
R39969 n3_7083_1727 n3_7083_1760 2.095238e-02
R39970 n3_7083_1760 n3_7083_1916 9.904762e-02
R39971 n3_7083_1916 n3_7083_1943 1.714286e-02
R39972 n3_7083_1943 n3_7083_1976 2.095238e-02
R39973 n3_7083_1976 n3_7083_2159 1.161905e-01
R39974 n3_7083_2159 n3_7083_2192 2.095238e-02
R39975 n3_7083_2192 n3_7083_2375 1.161905e-01
R39976 n3_7083_2375 n3_7083_2408 2.095238e-02
R39977 n3_7083_2408 n3_7083_2543 8.571429e-02
R39978 n3_7083_2543 n3_7083_2564 1.333333e-02
R39979 n3_7083_2564 n3_7083_2591 1.714286e-02
R39980 n3_7083_2591 n3_7083_2624 2.095238e-02
R39981 n3_7083_2624 n3_7083_2674 3.174603e-02
R39982 n3_7083_2674 n3_7083_2770 6.095238e-02
R39983 n3_7083_2770 n3_7083_2807 2.349206e-02
R39984 n3_7083_2807 n3_7083_2840 2.095238e-02
R39985 n3_7083_2840 n3_7083_2974 8.507937e-02
R39986 n3_7083_2974 n3_7083_2996 1.396825e-02
R39987 n3_7083_2996 n3_7083_3023 1.714286e-02
R39988 n3_7083_3023 n3_7083_3056 2.095238e-02
R39989 n3_7083_3056 n3_7083_3239 1.161905e-01
R39990 n3_7083_3239 n3_7083_3272 2.095238e-02
R39991 n3_7083_3272 n3_7083_3455 1.161905e-01
R39992 n3_7083_3455 n3_7083_3488 2.095238e-02
R39993 n3_7083_3488 n3_7083_3644 9.904762e-02
R39994 n3_7083_3644 n3_7083_3671 1.714286e-02
R39995 n3_7083_3671 n3_7083_3704 2.095238e-02
R39996 n3_7083_4103 n3_7083_4136 2.095238e-02
R39997 n3_7083_4136 n3_7083_4292 9.904762e-02
R39998 n3_7083_4292 n3_7083_4319 1.714286e-02
R39999 n3_7083_4319 n3_7083_4352 2.095238e-02
R40000 n3_7083_4352 n3_7083_4535 1.161905e-01
R40001 n3_7083_4535 n3_7083_4568 2.095238e-02
R40002 n3_7083_4568 n3_7083_4724 9.904762e-02
R40003 n3_7083_4724 n3_7083_4751 1.714286e-02
R40004 n3_7083_4751 n3_7083_4784 2.095238e-02
R40005 n3_7083_4784 n3_7083_4924 8.888889e-02
R40006 n3_7083_4924 n3_7083_4967 2.730159e-02
R40007 n3_7083_4967 n3_7083_5000 2.095238e-02
R40008 n3_7083_5000 n3_7083_5020 1.269841e-02
R40009 n3_7083_5020 n3_7083_5183 1.034921e-01
R40010 n3_7083_5183 n3_7083_5216 2.095238e-02
R40011 n3_7083_5216 n3_7083_5372 9.904762e-02
R40012 n3_7083_5372 n3_7083_5399 1.714286e-02
R40013 n3_7083_5399 n3_7083_5432 2.095238e-02
R40014 n3_7083_5432 n3_7083_5566 8.507937e-02
R40015 n3_7083_5566 n3_7083_5588 1.396825e-02
R40016 n3_7083_5588 n3_7083_5615 1.714286e-02
R40017 n3_7083_5615 n3_7083_5648 2.095238e-02
R40018 n3_7083_5648 n3_7083_5831 1.161905e-01
R40019 n3_7083_5831 n3_7083_5864 2.095238e-02
R40020 n3_7083_6263 n3_7083_6296 2.095238e-02
R40021 n3_7083_6296 n3_7083_6479 1.161905e-01
R40022 n3_7083_6479 n3_7083_6512 2.095238e-02
R40023 n3_7083_6512 n3_7083_6646 8.507937e-02
R40024 n3_7083_6646 n3_7083_6695 3.111111e-02
R40025 n3_7083_6695 n3_7083_6728 2.095238e-02
R40026 n3_7083_6728 n3_7083_6911 1.161905e-01
R40027 n3_7083_6911 n3_7083_6944 2.095238e-02
R40028 n3_7083_6944 n3_7083_7127 1.161905e-01
R40029 n3_7083_7127 n3_7083_7160 2.095238e-02
R40030 n3_7083_7160 n3_7083_7174 8.888889e-03
R40031 n3_7083_7174 n3_7083_7270 6.095238e-02
R40032 n3_7083_7270 n3_7083_7343 4.634921e-02
R40033 n3_7083_7343 n3_7083_7376 2.095238e-02
R40034 n3_7083_7376 n3_7083_7559 1.161905e-01
R40035 n3_7083_7559 n3_7083_7592 2.095238e-02
R40036 n3_7083_7592 n3_7083_7775 1.161905e-01
R40037 n3_7083_7775 n3_7083_7808 2.095238e-02
R40038 n3_7083_7808 n3_7083_7822 8.888889e-03
R40039 n3_7083_7822 n3_7083_7964 9.015873e-02
R40040 n3_7083_7964 n3_7083_7991 1.714286e-02
R40041 n3_7083_7991 n3_7083_8024 2.095238e-02
R40042 n3_7083_8024 n3_7083_8207 1.161905e-01
R40043 n3_7083_8207 n3_7083_8240 2.095238e-02
R40044 n3_7083_8456 n3_7083_8639 1.161905e-01
R40045 n3_7083_8639 n3_7083_8672 2.095238e-02
R40046 n3_7083_8672 n3_7083_8855 1.161905e-01
R40047 n3_7083_8855 n3_7083_8888 2.095238e-02
R40048 n3_7083_8888 n3_7083_8902 8.888889e-03
R40049 n3_7083_8902 n3_7083_9044 9.015873e-02
R40050 n3_7083_9044 n3_7083_9071 1.714286e-02
R40051 n3_7083_9071 n3_7083_9104 2.095238e-02
R40052 n3_7083_9104 n3_7083_9287 1.161905e-01
R40053 n3_7083_9287 n3_7083_9320 2.095238e-02
R40054 n3_7083_9320 n3_7083_9424 6.603175e-02
R40055 n3_7083_9424 n3_7083_9503 5.015873e-02
R40056 n3_7083_9503 n3_7083_9520 1.079365e-02
R40057 n3_7083_9520 n3_7083_9536 1.015873e-02
R40058 n3_7083_9536 n3_7083_9719 1.161905e-01
R40059 n3_7083_9719 n3_7083_9752 2.095238e-02
R40060 n3_7083_9752 n3_7083_9935 1.161905e-01
R40061 n3_7083_9935 n3_7083_9968 2.095238e-02
R40062 n3_7083_9968 n3_7083_9982 8.888889e-03
R40063 n3_7083_9982 n3_7083_10124 9.015873e-02
R40064 n3_7083_10124 n3_7083_10151 1.714286e-02
R40065 n3_7083_10151 n3_7083_10184 2.095238e-02
R40066 n3_7083_10184 n3_7083_10367 1.161905e-01
R40067 n3_7083_10367 n3_7083_10400 2.095238e-02
R40068 n3_7083_10799 n3_7083_10832 2.095238e-02
R40069 n3_7083_10832 n3_7083_11015 1.161905e-01
R40070 n3_7083_11015 n3_7083_11048 2.095238e-02
R40071 n3_7083_11048 n3_7083_11204 9.904762e-02
R40072 n3_7083_11204 n3_7083_11231 1.714286e-02
R40073 n3_7083_11231 n3_7083_11264 2.095238e-02
R40074 n3_7083_11264 n3_7083_11447 1.161905e-01
R40075 n3_7083_11447 n3_7083_11480 2.095238e-02
R40076 n3_7083_11480 n3_7083_11663 1.161905e-01
R40077 n3_7083_11663 n3_7083_11674 6.984127e-03
R40078 n3_7083_11674 n3_7083_11696 1.396825e-02
R40079 n3_7083_11696 n3_7083_11770 4.698413e-02
R40080 n3_7083_11770 n3_7083_11879 6.920635e-02
R40081 n3_7083_11879 n3_7083_11912 2.095238e-02
R40082 n3_7083_11912 n3_7083_12095 1.161905e-01
R40083 n3_7083_12095 n3_7083_12128 2.095238e-02
R40084 n3_7083_12128 n3_7083_12284 9.904762e-02
R40085 n3_7083_12284 n3_7083_12311 1.714286e-02
R40086 n3_7083_12311 n3_7083_12344 2.095238e-02
R40087 n3_7083_12344 n3_7083_12527 1.161905e-01
R40088 n3_7083_12527 n3_7083_12560 2.095238e-02
R40089 n3_7083_12560 n3_7083_12743 1.161905e-01
R40090 n3_7083_12959 n3_7083_12992 2.095238e-02
R40091 n3_7083_12992 n3_7083_13175 1.161905e-01
R40092 n3_7083_13175 n3_7083_13208 2.095238e-02
R40093 n3_7083_13208 n3_7083_13391 1.161905e-01
R40094 n3_7083_13391 n3_7083_13424 2.095238e-02
R40095 n3_7083_13424 n3_7083_13580 9.904762e-02
R40096 n3_7083_13580 n3_7083_13607 1.714286e-02
R40097 n3_7083_13607 n3_7083_13640 2.095238e-02
R40098 n3_7083_13640 n3_7083_13823 1.161905e-01
R40099 n3_7083_13823 n3_7083_13856 2.095238e-02
R40100 n3_7083_13856 n3_7083_13924 4.317460e-02
R40101 n3_7083_13924 n3_7083_14020 6.095238e-02
R40102 n3_7083_14020 n3_7083_14039 1.206349e-02
R40103 n3_7083_14039 n3_7083_14072 2.095238e-02
R40104 n3_7083_14072 n3_7083_14255 1.161905e-01
R40105 n3_7083_14255 n3_7083_14288 2.095238e-02
R40106 n3_7083_14288 n3_7083_14471 1.161905e-01
R40107 n3_7083_14471 n3_7083_14504 2.095238e-02
R40108 n3_7083_14504 n3_7083_14553 3.111111e-02
R40109 n3_7083_14553 n3_7083_14687 8.507937e-02
R40110 n3_7083_14687 n3_7083_14720 2.095238e-02
R40111 n3_7083_14720 n3_7083_14903 1.161905e-01
R40112 n3_7083_14903 n3_7083_14936 2.095238e-02
R40113 n3_7083_15335 n3_7083_15368 2.095238e-02
R40114 n3_7083_15368 n3_7083_15551 1.161905e-01
R40115 n3_7083_15551 n3_7083_15584 2.095238e-02
R40116 n3_7083_15584 n3_7083_15740 9.904762e-02
R40117 n3_7083_15740 n3_7083_15767 1.714286e-02
R40118 n3_7083_15767 n3_7083_15800 2.095238e-02
R40119 n3_7083_15800 n3_7083_15956 9.904762e-02
R40120 n3_7083_15956 n3_7083_15983 1.714286e-02
R40121 n3_7083_15983 n3_7083_16016 2.095238e-02
R40122 n3_7083_16016 n3_7083_16172 9.904762e-02
R40123 n3_7083_16172 n3_7083_16174 1.269841e-03
R40124 n3_7083_16174 n3_7083_16199 1.587302e-02
R40125 n3_7083_16199 n3_7083_16232 2.095238e-02
R40126 n3_7083_16232 n3_7083_16270 2.412698e-02
R40127 n3_7083_16270 n3_7083_16415 9.206349e-02
R40128 n3_7083_16415 n3_7083_16448 2.095238e-02
R40129 n3_7083_16448 n3_7083_16631 1.161905e-01
R40130 n3_7083_16631 n3_7083_16664 2.095238e-02
R40131 n3_7083_16664 n3_7083_16847 1.161905e-01
R40132 n3_7083_16847 n3_7083_16880 2.095238e-02
R40133 n3_7083_16880 n3_7083_17063 1.161905e-01
R40134 n3_7083_17063 n3_7083_17096 2.095238e-02
R40135 n3_7083_17096 n3_7083_17230 8.507937e-02
R40136 n3_7083_17468 n3_7083_17495 1.714286e-02
R40137 n3_7083_17495 n3_7083_17528 2.095238e-02
R40138 n3_7083_17528 n3_7083_17711 1.161905e-01
R40139 n3_7083_17711 n3_7083_17744 2.095238e-02
R40140 n3_7083_17744 n3_7083_17927 1.161905e-01
R40141 n3_7083_17927 n3_7083_17960 2.095238e-02
R40142 n3_7083_17960 n3_7083_18143 1.161905e-01
R40143 n3_7083_18143 n3_7083_18176 2.095238e-02
R40144 n3_7083_18176 n3_7083_18359 1.161905e-01
R40145 n3_7083_18359 n3_7083_18392 2.095238e-02
R40146 n3_7083_18392 n3_7083_18424 2.031746e-02
R40147 n3_7083_18424 n3_7083_18520 6.095238e-02
R40148 n3_7083_18520 n3_7083_18526 3.809524e-03
R40149 n3_7083_18526 n3_7083_18527 6.349206e-04
R40150 n3_7083_18527 n3_7083_18548 1.333333e-02
R40151 n3_7083_18548 n3_7083_18575 1.714286e-02
R40152 n3_7083_18575 n3_7083_18608 2.095238e-02
R40153 n3_7083_18608 n3_7083_18764 9.904762e-02
R40154 n3_7083_18764 n3_7083_18791 1.714286e-02
R40155 n3_7083_18791 n3_7083_18824 2.095238e-02
R40156 n3_7083_18824 n3_7083_19007 1.161905e-01
R40157 n3_7083_19007 n3_7083_19040 2.095238e-02
R40158 n3_7083_19040 n3_7083_19196 9.904762e-02
R40159 n3_7083_19196 n3_7083_19223 1.714286e-02
R40160 n3_7083_19223 n3_7083_19256 2.095238e-02
R40161 n3_7083_19256 n3_7083_19390 8.507937e-02
R40162 n3_7083_19390 n3_7083_19439 3.111111e-02
R40163 n3_7083_19439 n3_7083_19472 2.095238e-02
R40164 n3_7083_19871 n3_7083_19904 2.095238e-02
R40165 n3_7083_19904 n3_7083_20087 1.161905e-01
R40166 n3_7083_20087 n3_7083_20120 2.095238e-02
R40167 n3_7083_20120 n3_7083_20303 1.161905e-01
R40168 n3_7083_20303 n3_7083_20336 2.095238e-02
R40169 n3_7083_20336 n3_7083_20519 1.161905e-01
R40170 n3_7083_20519 n3_7083_20552 2.095238e-02
R40171 n3_7083_20552 n3_7083_20674 7.746032e-02
R40172 n3_7083_20674 n3_7083_20687 8.253968e-03
R40173 n3_7083_20687 n3_7083_20735 3.047619e-02
R40174 n3_7083_20735 n3_7083_20768 2.095238e-02
R40175 n3_7083_20768 n3_7083_20770 1.269841e-03
R40176 n3_7083_20770 n3_7083_20951 1.149206e-01
R40177 n3_7083_20951 n3_7083_20984 2.095238e-02
R40178 n3_7271_215 n3_7271_248 2.095238e-02
R40179 n3_7271_248 n3_7271_383 8.571429e-02
R40180 n3_7271_383 n3_7271_424 2.603175e-02
R40181 n3_7271_424 n3_7271_431 4.444444e-03
R40182 n3_7271_520 n3_7271_647 8.063492e-02
R40183 n3_7271_647 n3_7271_680 2.095238e-02
R40184 n3_7271_680 n3_7271_863 1.161905e-01
R40185 n3_7271_863 n3_7271_896 2.095238e-02
R40186 n3_7271_896 n3_7271_1079 1.161905e-01
R40187 n3_7271_1079 n3_7271_1112 2.095238e-02
R40188 n3_7271_1112 n3_7271_1295 1.161905e-01
R40189 n3_7271_1295 n3_7271_1328 2.095238e-02
R40190 n3_7271_1328 n3_7271_1511 1.161905e-01
R40191 n3_7271_1511 n3_7271_1544 2.095238e-02
R40192 n3_7271_1544 n3_7271_1727 1.161905e-01
R40193 n3_7271_1727 n3_7271_1760 2.095238e-02
R40194 n3_7271_1760 n3_7271_1916 9.904762e-02
R40195 n3_7271_1916 n3_7271_1943 1.714286e-02
R40196 n3_7271_1943 n3_7271_1976 2.095238e-02
R40197 n3_7271_1976 n3_7271_2159 1.161905e-01
R40198 n3_7271_2159 n3_7271_2192 2.095238e-02
R40199 n3_7271_2192 n3_7271_2375 1.161905e-01
R40200 n3_7271_2375 n3_7271_2408 2.095238e-02
R40201 n3_7271_2408 n3_7271_2543 8.571429e-02
R40202 n3_7271_2543 n3_7271_2564 1.333333e-02
R40203 n3_7271_2564 n3_7271_2591 1.714286e-02
R40204 n3_7271_2591 n3_7271_2624 2.095238e-02
R40205 n3_7271_2624 n3_7271_2674 3.174603e-02
R40206 n3_7271_2770 n3_7271_2807 2.349206e-02
R40207 n3_7271_2807 n3_7271_2840 2.095238e-02
R40208 n3_7271_2840 n3_7271_2974 8.507937e-02
R40209 n3_7271_2974 n3_7271_2996 1.396825e-02
R40210 n3_7271_2996 n3_7271_3023 1.714286e-02
R40211 n3_7271_3023 n3_7271_3056 2.095238e-02
R40212 n3_7271_3056 n3_7271_3239 1.161905e-01
R40213 n3_7271_3239 n3_7271_3272 2.095238e-02
R40214 n3_7271_3272 n3_7271_3455 1.161905e-01
R40215 n3_7271_3455 n3_7271_3488 2.095238e-02
R40216 n3_7271_3488 n3_7271_3644 9.904762e-02
R40217 n3_7271_3644 n3_7271_3671 1.714286e-02
R40218 n3_7271_3671 n3_7271_3704 2.095238e-02
R40219 n3_7271_3704 n3_7271_3887 1.161905e-01
R40220 n3_7271_3887 n3_7271_3920 2.095238e-02
R40221 n3_7271_3920 n3_7271_4103 1.161905e-01
R40222 n3_7271_4103 n3_7271_4136 2.095238e-02
R40223 n3_7271_4136 n3_7271_4292 9.904762e-02
R40224 n3_7271_4292 n3_7271_4319 1.714286e-02
R40225 n3_7271_4319 n3_7271_4352 2.095238e-02
R40226 n3_7271_4352 n3_7271_4535 1.161905e-01
R40227 n3_7271_4535 n3_7271_4568 2.095238e-02
R40228 n3_7271_4568 n3_7271_4724 9.904762e-02
R40229 n3_7271_4724 n3_7271_4751 1.714286e-02
R40230 n3_7271_4751 n3_7271_4784 2.095238e-02
R40231 n3_7271_4784 n3_7271_4924 8.888889e-02
R40232 n3_7271_5000 n3_7271_5020 1.269841e-02
R40233 n3_7271_5020 n3_7271_5183 1.034921e-01
R40234 n3_7271_5183 n3_7271_5216 2.095238e-02
R40235 n3_7271_5216 n3_7271_5372 9.904762e-02
R40236 n3_7271_5372 n3_7271_5399 1.714286e-02
R40237 n3_7271_5399 n3_7271_5432 2.095238e-02
R40238 n3_7271_5432 n3_7271_5566 8.507937e-02
R40239 n3_7271_5566 n3_7271_5588 1.396825e-02
R40240 n3_7271_5588 n3_7271_5615 1.714286e-02
R40241 n3_7271_5615 n3_7271_5648 2.095238e-02
R40242 n3_7271_5648 n3_7271_5831 1.161905e-01
R40243 n3_7271_5831 n3_7271_5864 2.095238e-02
R40244 n3_7271_5864 n3_7271_6047 1.161905e-01
R40245 n3_7271_6047 n3_7271_6080 2.095238e-02
R40246 n3_7271_6080 n3_7271_6263 1.161905e-01
R40247 n3_7271_6263 n3_7271_6296 2.095238e-02
R40248 n3_7271_6296 n3_7271_6479 1.161905e-01
R40249 n3_7271_6479 n3_7271_6512 2.095238e-02
R40250 n3_7271_6512 n3_7271_6646 8.507937e-02
R40251 n3_7271_6646 n3_7271_6695 3.111111e-02
R40252 n3_7271_6695 n3_7271_6728 2.095238e-02
R40253 n3_7271_6728 n3_7271_6911 1.161905e-01
R40254 n3_7271_6911 n3_7271_6944 2.095238e-02
R40255 n3_7271_6944 n3_7271_7127 1.161905e-01
R40256 n3_7271_7127 n3_7271_7160 2.095238e-02
R40257 n3_7271_7160 n3_7271_7174 8.888889e-03
R40258 n3_7271_7270 n3_7271_7343 4.634921e-02
R40259 n3_7271_7343 n3_7271_7376 2.095238e-02
R40260 n3_7271_7376 n3_7271_7559 1.161905e-01
R40261 n3_7271_7559 n3_7271_7592 2.095238e-02
R40262 n3_7271_7592 n3_7271_7775 1.161905e-01
R40263 n3_7271_7775 n3_7271_7808 2.095238e-02
R40264 n3_7271_7808 n3_7271_7822 8.888889e-03
R40265 n3_7271_7822 n3_7271_7964 9.015873e-02
R40266 n3_7271_7964 n3_7271_7991 1.714286e-02
R40267 n3_7271_7991 n3_7271_8024 2.095238e-02
R40268 n3_7271_8024 n3_7271_8207 1.161905e-01
R40269 n3_7271_8207 n3_7271_8240 2.095238e-02
R40270 n3_7271_8240 n3_7271_8423 1.161905e-01
R40271 n3_7271_8423 n3_7271_8456 2.095238e-02
R40272 n3_7271_8456 n3_7271_8639 1.161905e-01
R40273 n3_7271_8639 n3_7271_8672 2.095238e-02
R40274 n3_7271_8672 n3_7271_8855 1.161905e-01
R40275 n3_7271_8855 n3_7271_8888 2.095238e-02
R40276 n3_7271_8888 n3_7271_8902 8.888889e-03
R40277 n3_7271_8902 n3_7271_9044 9.015873e-02
R40278 n3_7271_9044 n3_7271_9071 1.714286e-02
R40279 n3_7271_9071 n3_7271_9104 2.095238e-02
R40280 n3_7271_9104 n3_7271_9287 1.161905e-01
R40281 n3_7271_9287 n3_7271_9320 2.095238e-02
R40282 n3_7271_9320 n3_7271_9424 6.603175e-02
R40283 n3_7271_9503 n3_7271_9520 1.079365e-02
R40284 n3_7271_9520 n3_7271_9536 1.015873e-02
R40285 n3_7271_9536 n3_7271_9719 1.161905e-01
R40286 n3_7271_9719 n3_7271_9752 2.095238e-02
R40287 n3_7271_9752 n3_7271_9935 1.161905e-01
R40288 n3_7271_9935 n3_7271_9968 2.095238e-02
R40289 n3_7271_9968 n3_7271_9982 8.888889e-03
R40290 n3_7271_9982 n3_7271_10124 9.015873e-02
R40291 n3_7271_10124 n3_7271_10151 1.714286e-02
R40292 n3_7271_10151 n3_7271_10184 2.095238e-02
R40293 n3_7271_10184 n3_7271_10367 1.161905e-01
R40294 n3_7271_10367 n3_7271_10400 2.095238e-02
R40295 n3_7271_10616 n3_7271_10799 1.161905e-01
R40296 n3_7271_10799 n3_7271_10832 2.095238e-02
R40297 n3_7271_10832 n3_7271_11015 1.161905e-01
R40298 n3_7271_11015 n3_7271_11048 2.095238e-02
R40299 n3_7271_11048 n3_7271_11204 9.904762e-02
R40300 n3_7271_11204 n3_7271_11231 1.714286e-02
R40301 n3_7271_11231 n3_7271_11264 2.095238e-02
R40302 n3_7271_11264 n3_7271_11447 1.161905e-01
R40303 n3_7271_11447 n3_7271_11480 2.095238e-02
R40304 n3_7271_11480 n3_7271_11663 1.161905e-01
R40305 n3_7271_11663 n3_7271_11674 6.984127e-03
R40306 n3_7271_11674 n3_7271_11696 1.396825e-02
R40307 n3_7271_11770 n3_7271_11879 6.920635e-02
R40308 n3_7271_11879 n3_7271_11912 2.095238e-02
R40309 n3_7271_11912 n3_7271_12095 1.161905e-01
R40310 n3_7271_12095 n3_7271_12128 2.095238e-02
R40311 n3_7271_12128 n3_7271_12284 9.904762e-02
R40312 n3_7271_12284 n3_7271_12311 1.714286e-02
R40313 n3_7271_12311 n3_7271_12344 2.095238e-02
R40314 n3_7271_12344 n3_7271_12527 1.161905e-01
R40315 n3_7271_12527 n3_7271_12560 2.095238e-02
R40316 n3_7271_12560 n3_7271_12743 1.161905e-01
R40317 n3_7271_12743 n3_7271_12776 2.095238e-02
R40318 n3_7271_12776 n3_7271_12959 1.161905e-01
R40319 n3_7271_12959 n3_7271_12992 2.095238e-02
R40320 n3_7271_12992 n3_7271_13175 1.161905e-01
R40321 n3_7271_13175 n3_7271_13208 2.095238e-02
R40322 n3_7271_13208 n3_7271_13391 1.161905e-01
R40323 n3_7271_13391 n3_7271_13424 2.095238e-02
R40324 n3_7271_13424 n3_7271_13580 9.904762e-02
R40325 n3_7271_13580 n3_7271_13607 1.714286e-02
R40326 n3_7271_13607 n3_7271_13640 2.095238e-02
R40327 n3_7271_13640 n3_7271_13823 1.161905e-01
R40328 n3_7271_13823 n3_7271_13856 2.095238e-02
R40329 n3_7271_13856 n3_7271_13924 4.317460e-02
R40330 n3_7271_14020 n3_7271_14039 1.206349e-02
R40331 n3_7271_14039 n3_7271_14072 2.095238e-02
R40332 n3_7271_14072 n3_7271_14255 1.161905e-01
R40333 n3_7271_14255 n3_7271_14288 2.095238e-02
R40334 n3_7271_14288 n3_7271_14471 1.161905e-01
R40335 n3_7271_14471 n3_7271_14504 2.095238e-02
R40336 n3_7271_14504 n3_7271_14553 3.111111e-02
R40337 n3_7271_14553 n3_7271_14687 8.507937e-02
R40338 n3_7271_14687 n3_7271_14720 2.095238e-02
R40339 n3_7271_14720 n3_7271_14903 1.161905e-01
R40340 n3_7271_14903 n3_7271_14936 2.095238e-02
R40341 n3_7271_14936 n3_7271_15119 1.161905e-01
R40342 n3_7271_15119 n3_7271_15152 2.095238e-02
R40343 n3_7271_15152 n3_7271_15335 1.161905e-01
R40344 n3_7271_15335 n3_7271_15368 2.095238e-02
R40345 n3_7271_15368 n3_7271_15551 1.161905e-01
R40346 n3_7271_15551 n3_7271_15584 2.095238e-02
R40347 n3_7271_15584 n3_7271_15740 9.904762e-02
R40348 n3_7271_15740 n3_7271_15767 1.714286e-02
R40349 n3_7271_15767 n3_7271_15800 2.095238e-02
R40350 n3_7271_15800 n3_7271_15956 9.904762e-02
R40351 n3_7271_15956 n3_7271_15983 1.714286e-02
R40352 n3_7271_15983 n3_7271_16016 2.095238e-02
R40353 n3_7271_16016 n3_7271_16172 9.904762e-02
R40354 n3_7271_16172 n3_7271_16174 1.269841e-03
R40355 n3_7271_16174 n3_7271_16199 1.587302e-02
R40356 n3_7271_16270 n3_7271_16415 9.206349e-02
R40357 n3_7271_16415 n3_7271_16448 2.095238e-02
R40358 n3_7271_16448 n3_7271_16631 1.161905e-01
R40359 n3_7271_16631 n3_7271_16664 2.095238e-02
R40360 n3_7271_16664 n3_7271_16847 1.161905e-01
R40361 n3_7271_16847 n3_7271_16880 2.095238e-02
R40362 n3_7271_16880 n3_7271_17063 1.161905e-01
R40363 n3_7271_17063 n3_7271_17096 2.095238e-02
R40364 n3_7271_17096 n3_7271_17230 8.507937e-02
R40365 n3_7271_17230 n3_7271_17252 1.396825e-02
R40366 n3_7271_17252 n3_7271_17279 1.714286e-02
R40367 n3_7271_17279 n3_7271_17312 2.095238e-02
R40368 n3_7271_17312 n3_7271_17468 9.904762e-02
R40369 n3_7271_17468 n3_7271_17495 1.714286e-02
R40370 n3_7271_17495 n3_7271_17528 2.095238e-02
R40371 n3_7271_17528 n3_7271_17711 1.161905e-01
R40372 n3_7271_17711 n3_7271_17744 2.095238e-02
R40373 n3_7271_17744 n3_7271_17927 1.161905e-01
R40374 n3_7271_17927 n3_7271_17960 2.095238e-02
R40375 n3_7271_17960 n3_7271_18143 1.161905e-01
R40376 n3_7271_18143 n3_7271_18176 2.095238e-02
R40377 n3_7271_18176 n3_7271_18359 1.161905e-01
R40378 n3_7271_18359 n3_7271_18392 2.095238e-02
R40379 n3_7271_18392 n3_7271_18424 2.031746e-02
R40380 n3_7271_18520 n3_7271_18526 3.809524e-03
R40381 n3_7271_18526 n3_7271_18527 6.349206e-04
R40382 n3_7271_18527 n3_7271_18548 1.333333e-02
R40383 n3_7271_18548 n3_7271_18575 1.714286e-02
R40384 n3_7271_18575 n3_7271_18608 2.095238e-02
R40385 n3_7271_18608 n3_7271_18764 9.904762e-02
R40386 n3_7271_18764 n3_7271_18791 1.714286e-02
R40387 n3_7271_18791 n3_7271_18824 2.095238e-02
R40388 n3_7271_18824 n3_7271_19007 1.161905e-01
R40389 n3_7271_19007 n3_7271_19040 2.095238e-02
R40390 n3_7271_19040 n3_7271_19196 9.904762e-02
R40391 n3_7271_19196 n3_7271_19223 1.714286e-02
R40392 n3_7271_19223 n3_7271_19256 2.095238e-02
R40393 n3_7271_19256 n3_7271_19390 8.507937e-02
R40394 n3_7271_19390 n3_7271_19439 3.111111e-02
R40395 n3_7271_19439 n3_7271_19472 2.095238e-02
R40396 n3_7271_19472 n3_7271_19655 1.161905e-01
R40397 n3_7271_19655 n3_7271_19688 2.095238e-02
R40398 n3_7271_19688 n3_7271_19871 1.161905e-01
R40399 n3_7271_19871 n3_7271_19904 2.095238e-02
R40400 n3_7271_19904 n3_7271_20087 1.161905e-01
R40401 n3_7271_20087 n3_7271_20120 2.095238e-02
R40402 n3_7271_20120 n3_7271_20303 1.161905e-01
R40403 n3_7271_20303 n3_7271_20336 2.095238e-02
R40404 n3_7271_20336 n3_7271_20519 1.161905e-01
R40405 n3_7271_20519 n3_7271_20552 2.095238e-02
R40406 n3_7271_20552 n3_7271_20674 7.746032e-02
R40407 n3_7271_20674 n3_7271_20687 8.253968e-03
R40408 n3_7271_20768 n3_7271_20770 1.269841e-03
R40409 n3_7271_20770 n3_7271_20951 1.149206e-01
R40410 n3_7271_20951 n3_7271_20984 2.095238e-02
R40411 n3_7364_215 n3_7364_248 2.095238e-02
R40412 n3_7364_248 n3_7364_383 8.571429e-02
R40413 n3_7364_383 n3_7364_431 3.047619e-02
R40414 n3_7364_431 n3_7364_464 2.095238e-02
R40415 n3_7364_464 n3_7364_647 1.161905e-01
R40416 n3_7364_647 n3_7364_680 2.095238e-02
R40417 n3_7364_680 n3_7364_863 1.161905e-01
R40418 n3_7364_863 n3_7364_896 2.095238e-02
R40419 n3_7364_896 n3_7364_1079 1.161905e-01
R40420 n3_7364_1079 n3_7364_1112 2.095238e-02
R40421 n3_7364_1112 n3_7364_1295 1.161905e-01
R40422 n3_7364_1295 n3_7364_1328 2.095238e-02
R40423 n3_7364_1328 n3_7364_1511 1.161905e-01
R40424 n3_7364_1511 n3_7364_1544 2.095238e-02
R40425 n3_7364_1544 n3_7364_1727 1.161905e-01
R40426 n3_7364_1727 n3_7364_1760 2.095238e-02
R40427 n3_7364_1760 n3_7364_1916 9.904762e-02
R40428 n3_7364_1916 n3_7364_1943 1.714286e-02
R40429 n3_7364_1943 n3_7364_1976 2.095238e-02
R40430 n3_7364_1976 n3_7364_2159 1.161905e-01
R40431 n3_7364_2159 n3_7364_2192 2.095238e-02
R40432 n3_7364_2192 n3_7364_2375 1.161905e-01
R40433 n3_7364_2375 n3_7364_2408 2.095238e-02
R40434 n3_7364_2408 n3_7364_2543 8.571429e-02
R40435 n3_7364_2543 n3_7364_2564 1.333333e-02
R40436 n3_7364_2564 n3_7364_2591 1.714286e-02
R40437 n3_7364_2591 n3_7364_2624 2.095238e-02
R40438 n3_7364_18526 n3_7364_18527 6.349206e-04
R40439 n3_7364_18527 n3_7364_18575 3.047619e-02
R40440 n3_7364_18575 n3_7364_18608 2.095238e-02
R40441 n3_7364_18608 n3_7364_18764 9.904762e-02
R40442 n3_7364_18764 n3_7364_18791 1.714286e-02
R40443 n3_7364_18791 n3_7364_18824 2.095238e-02
R40444 n3_7364_18824 n3_7364_19007 1.161905e-01
R40445 n3_7364_19007 n3_7364_19040 2.095238e-02
R40446 n3_7364_19040 n3_7364_19223 1.161905e-01
R40447 n3_7364_19223 n3_7364_19256 2.095238e-02
R40448 n3_7364_19256 n3_7364_19390 8.507937e-02
R40449 n3_7364_19390 n3_7364_19439 3.111111e-02
R40450 n3_7364_19439 n3_7364_19472 2.095238e-02
R40451 n3_7364_19472 n3_7364_19655 1.161905e-01
R40452 n3_7364_19655 n3_7364_19688 2.095238e-02
R40453 n3_7364_19688 n3_7364_19871 1.161905e-01
R40454 n3_7364_19871 n3_7364_19904 2.095238e-02
R40455 n3_7364_19904 n3_7364_20087 1.161905e-01
R40456 n3_7364_20087 n3_7364_20120 2.095238e-02
R40457 n3_7364_20120 n3_7364_20303 1.161905e-01
R40458 n3_7364_20303 n3_7364_20336 2.095238e-02
R40459 n3_7364_20336 n3_7364_20519 1.161905e-01
R40460 n3_7364_20519 n3_7364_20552 2.095238e-02
R40461 n3_7364_20552 n3_7364_20687 8.571429e-02
R40462 n3_7364_20687 n3_7364_20735 3.047619e-02
R40463 n3_7364_20735 n3_7364_20768 2.095238e-02
R40464 n3_7364_20768 n3_7364_20951 1.161905e-01
R40465 n3_7364_20951 n3_7364_20984 2.095238e-02
R40466 n3_9150_215 n3_9150_248 2.095238e-02
R40467 n3_9150_248 n3_9150_383 8.571429e-02
R40468 n3_9150_383 n3_9150_431 3.047619e-02
R40469 n3_9150_431 n3_9150_464 2.095238e-02
R40470 n3_9150_464 n3_9150_647 1.161905e-01
R40471 n3_9150_647 n3_9150_680 2.095238e-02
R40472 n3_9150_680 n3_9150_863 1.161905e-01
R40473 n3_9150_863 n3_9150_896 2.095238e-02
R40474 n3_9150_896 n3_9150_1079 1.161905e-01
R40475 n3_9150_1079 n3_9150_1112 2.095238e-02
R40476 n3_9150_1112 n3_9150_1295 1.161905e-01
R40477 n3_9150_1295 n3_9150_1328 2.095238e-02
R40478 n3_9150_1328 n3_9150_1511 1.161905e-01
R40479 n3_9150_1511 n3_9150_1544 2.095238e-02
R40480 n3_9150_1544 n3_9150_1727 1.161905e-01
R40481 n3_9150_1727 n3_9150_1760 2.095238e-02
R40482 n3_9150_1760 n3_9150_1894 8.507937e-02
R40483 n3_9150_1894 n3_9150_1943 3.111111e-02
R40484 n3_9150_1943 n3_9150_1976 2.095238e-02
R40485 n3_9150_1976 n3_9150_2159 1.161905e-01
R40486 n3_9150_2159 n3_9150_2192 2.095238e-02
R40487 n3_9150_2192 n3_9150_2375 1.161905e-01
R40488 n3_9150_2375 n3_9150_2408 2.095238e-02
R40489 n3_9150_2408 n3_9150_2543 8.571429e-02
R40490 n3_9150_2543 n3_9150_2564 1.333333e-02
R40491 n3_9150_2564 n3_9150_2591 1.714286e-02
R40492 n3_9150_2591 n3_9150_2624 2.095238e-02
R40493 n3_9150_18527 n3_9150_18548 1.333333e-02
R40494 n3_9150_18548 n3_9150_18575 1.714286e-02
R40495 n3_9150_18575 n3_9150_18608 2.095238e-02
R40496 n3_9150_18608 n3_9150_18764 9.904762e-02
R40497 n3_9150_18764 n3_9150_18791 1.714286e-02
R40498 n3_9150_18791 n3_9150_18824 2.095238e-02
R40499 n3_9150_18824 n3_9150_19007 1.161905e-01
R40500 n3_9150_19007 n3_9150_19040 2.095238e-02
R40501 n3_9150_19040 n3_9150_19223 1.161905e-01
R40502 n3_9150_19223 n3_9150_19256 2.095238e-02
R40503 n3_9150_19256 n3_9150_19412 9.904762e-02
R40504 n3_9150_19412 n3_9150_19439 1.714286e-02
R40505 n3_9150_19439 n3_9150_19472 2.095238e-02
R40506 n3_9150_19472 n3_9150_19655 1.161905e-01
R40507 n3_9150_19655 n3_9150_19688 2.095238e-02
R40508 n3_9150_19688 n3_9150_19871 1.161905e-01
R40509 n3_9150_19871 n3_9150_19904 2.095238e-02
R40510 n3_9150_19904 n3_9150_20087 1.161905e-01
R40511 n3_9150_20087 n3_9150_20120 2.095238e-02
R40512 n3_9150_20120 n3_9150_20303 1.161905e-01
R40513 n3_9150_20303 n3_9150_20336 2.095238e-02
R40514 n3_9150_20336 n3_9150_20519 1.161905e-01
R40515 n3_9150_20519 n3_9150_20552 2.095238e-02
R40516 n3_9150_20552 n3_9150_20687 8.571429e-02
R40517 n3_9150_20687 n3_9150_20735 3.047619e-02
R40518 n3_9150_20735 n3_9150_20768 2.095238e-02
R40519 n3_9150_20768 n3_9150_20951 1.161905e-01
R40520 n3_9150_20951 n3_9150_20984 2.095238e-02
R40521 n3_9333_424 n3_9380_424 2.984127e-02
R40522 n3_9380_424 n3_9521_424 8.952381e-02
R40523 n3_9333_520 n3_9380_520 2.984127e-02
R40524 n3_9380_520 n3_9521_520 8.952381e-02
R40525 n3_9333_2674 n3_9380_2674 2.984127e-02
R40526 n3_9380_2674 n3_9521_2674 8.952381e-02
R40527 n3_9333_2770 n3_9380_2770 2.984127e-02
R40528 n3_9380_2770 n3_9521_2770 8.952381e-02
R40529 n3_9333_4924 n3_9380_4924 2.984127e-02
R40530 n3_9380_4924 n3_9521_4924 8.952381e-02
R40531 n3_9333_5020 n3_9380_5020 2.984127e-02
R40532 n3_9380_5020 n3_9521_5020 8.952381e-02
R40533 n3_9333_7174 n3_9380_7174 2.984127e-02
R40534 n3_9380_7174 n3_9521_7174 8.952381e-02
R40535 n3_9333_7270 n3_9380_7270 2.984127e-02
R40536 n3_9380_7270 n3_9521_7270 8.952381e-02
R40537 n3_9333_9424 n3_9380_9424 2.984127e-02
R40538 n3_9380_9424 n3_9521_9424 8.952381e-02
R40539 n3_9333_9520 n3_9380_9520 2.984127e-02
R40540 n3_9380_9520 n3_9521_9520 8.952381e-02
R40541 n3_9333_11674 n3_9380_11674 2.984127e-02
R40542 n3_9380_11674 n3_9521_11674 8.952381e-02
R40543 n3_9333_11770 n3_9380_11770 2.984127e-02
R40544 n3_9380_11770 n3_9521_11770 8.952381e-02
R40545 n3_9333_13924 n3_9380_13924 2.984127e-02
R40546 n3_9380_13924 n3_9521_13924 8.952381e-02
R40547 n3_9333_14020 n3_9380_14020 2.984127e-02
R40548 n3_9380_14020 n3_9521_14020 8.952381e-02
R40549 n3_9333_16174 n3_9380_16174 2.984127e-02
R40550 n3_9380_16174 n3_9521_16174 8.952381e-02
R40551 n3_9333_16270 n3_9380_16270 2.984127e-02
R40552 n3_9380_16270 n3_9521_16270 8.952381e-02
R40553 n3_9333_18424 n3_9380_18424 2.984127e-02
R40554 n3_9380_18424 n3_9521_18424 8.952381e-02
R40555 n3_9333_18520 n3_9380_18520 2.984127e-02
R40556 n3_9380_18520 n3_9521_18520 8.952381e-02
R40557 n3_9333_20674 n3_9380_20674 2.984127e-02
R40558 n3_9380_20674 n3_9521_20674 8.952381e-02
R40559 n3_9333_20770 n3_9380_20770 2.984127e-02
R40560 n3_9380_20770 n3_9521_20770 8.952381e-02
R40561 n3_9333_215 n3_9333_248 2.095238e-02
R40562 n3_9333_248 n3_9333_383 8.571429e-02
R40563 n3_9333_383 n3_9333_424 2.603175e-02
R40564 n3_9333_424 n3_9333_431 4.444444e-03
R40565 n3_9333_431 n3_9333_464 2.095238e-02
R40566 n3_9333_464 n3_9333_520 3.555556e-02
R40567 n3_9333_520 n3_9333_647 8.063492e-02
R40568 n3_9333_647 n3_9333_680 2.095238e-02
R40569 n3_9333_680 n3_9333_863 1.161905e-01
R40570 n3_9333_863 n3_9333_896 2.095238e-02
R40571 n3_9333_896 n3_9333_1079 1.161905e-01
R40572 n3_9333_1079 n3_9333_1112 2.095238e-02
R40573 n3_9333_1112 n3_9333_1295 1.161905e-01
R40574 n3_9333_1295 n3_9333_1328 2.095238e-02
R40575 n3_9333_1727 n3_9333_1760 2.095238e-02
R40576 n3_9333_1760 n3_9333_1894 8.507937e-02
R40577 n3_9333_1894 n3_9333_1916 1.396825e-02
R40578 n3_9333_1916 n3_9333_1943 1.714286e-02
R40579 n3_9333_1943 n3_9333_1976 2.095238e-02
R40580 n3_9333_1976 n3_9333_2159 1.161905e-01
R40581 n3_9333_2159 n3_9333_2192 2.095238e-02
R40582 n3_9333_2192 n3_9333_2375 1.161905e-01
R40583 n3_9333_2375 n3_9333_2408 2.095238e-02
R40584 n3_9333_2408 n3_9333_2543 8.571429e-02
R40585 n3_9333_2543 n3_9333_2564 1.333333e-02
R40586 n3_9333_2564 n3_9333_2591 1.714286e-02
R40587 n3_9333_2591 n3_9333_2624 2.095238e-02
R40588 n3_9333_2624 n3_9333_2674 3.174603e-02
R40589 n3_9333_2674 n3_9333_2770 6.095238e-02
R40590 n3_9333_2770 n3_9333_2807 2.349206e-02
R40591 n3_9333_2807 n3_9333_2840 2.095238e-02
R40592 n3_9333_2840 n3_9333_2996 9.904762e-02
R40593 n3_9333_2996 n3_9333_3023 1.714286e-02
R40594 n3_9333_3023 n3_9333_3056 2.095238e-02
R40595 n3_9333_3056 n3_9333_3239 1.161905e-01
R40596 n3_9333_3239 n3_9333_3272 2.095238e-02
R40597 n3_9333_3272 n3_9333_3455 1.161905e-01
R40598 n3_9333_3455 n3_9333_3488 2.095238e-02
R40599 n3_9333_3488 n3_9333_3644 9.904762e-02
R40600 n3_9333_3644 n3_9333_3671 1.714286e-02
R40601 n3_9333_3671 n3_9333_3704 2.095238e-02
R40602 n3_9333_4103 n3_9333_4136 2.095238e-02
R40603 n3_9333_4136 n3_9333_4292 9.904762e-02
R40604 n3_9333_4292 n3_9333_4319 1.714286e-02
R40605 n3_9333_4319 n3_9333_4352 2.095238e-02
R40606 n3_9333_4352 n3_9333_4535 1.161905e-01
R40607 n3_9333_4535 n3_9333_4568 2.095238e-02
R40608 n3_9333_4568 n3_9333_4724 9.904762e-02
R40609 n3_9333_4724 n3_9333_4751 1.714286e-02
R40610 n3_9333_4751 n3_9333_4784 2.095238e-02
R40611 n3_9333_4784 n3_9333_4924 8.888889e-02
R40612 n3_9333_4924 n3_9333_4967 2.730159e-02
R40613 n3_9333_4967 n3_9333_5000 2.095238e-02
R40614 n3_9333_5000 n3_9333_5020 1.269841e-02
R40615 n3_9333_5020 n3_9333_5183 1.034921e-01
R40616 n3_9333_5183 n3_9333_5216 2.095238e-02
R40617 n3_9333_5216 n3_9333_5350 8.507937e-02
R40618 n3_9333_5350 n3_9333_5372 1.396825e-02
R40619 n3_9333_5372 n3_9333_5399 1.714286e-02
R40620 n3_9333_5399 n3_9333_5432 2.095238e-02
R40621 n3_9333_5432 n3_9333_5588 9.904762e-02
R40622 n3_9333_5588 n3_9333_5615 1.714286e-02
R40623 n3_9333_5615 n3_9333_5648 2.095238e-02
R40624 n3_9333_5648 n3_9333_5831 1.161905e-01
R40625 n3_9333_5831 n3_9333_5864 2.095238e-02
R40626 n3_9333_6263 n3_9333_6296 2.095238e-02
R40627 n3_9333_6296 n3_9333_6479 1.161905e-01
R40628 n3_9333_6479 n3_9333_6512 2.095238e-02
R40629 n3_9333_6512 n3_9333_6668 9.904762e-02
R40630 n3_9333_6668 n3_9333_6695 1.714286e-02
R40631 n3_9333_6695 n3_9333_6728 2.095238e-02
R40632 n3_9333_6728 n3_9333_6911 1.161905e-01
R40633 n3_9333_6911 n3_9333_6944 2.095238e-02
R40634 n3_9333_6944 n3_9333_7100 9.904762e-02
R40635 n3_9333_7100 n3_9333_7127 1.714286e-02
R40636 n3_9333_7127 n3_9333_7160 2.095238e-02
R40637 n3_9333_7160 n3_9333_7174 8.888889e-03
R40638 n3_9333_7174 n3_9333_7270 6.095238e-02
R40639 n3_9333_7270 n3_9333_7316 2.920635e-02
R40640 n3_9333_7316 n3_9333_7343 1.714286e-02
R40641 n3_9333_7343 n3_9333_7376 2.095238e-02
R40642 n3_9333_7376 n3_9333_7532 9.904762e-02
R40643 n3_9333_7532 n3_9333_7559 1.714286e-02
R40644 n3_9333_7559 n3_9333_7592 2.095238e-02
R40645 n3_9333_7592 n3_9333_7775 1.161905e-01
R40646 n3_9333_7775 n3_9333_7808 2.095238e-02
R40647 n3_9333_7808 n3_9333_7991 1.161905e-01
R40648 n3_9333_7991 n3_9333_8024 2.095238e-02
R40649 n3_9333_8024 n3_9333_8207 1.161905e-01
R40650 n3_9333_8207 n3_9333_8240 2.095238e-02
R40651 n3_9333_8456 n3_9333_8639 1.161905e-01
R40652 n3_9333_8639 n3_9333_8672 2.095238e-02
R40653 n3_9333_8672 n3_9333_8855 1.161905e-01
R40654 n3_9333_8855 n3_9333_8888 2.095238e-02
R40655 n3_9333_8888 n3_9333_9071 1.161905e-01
R40656 n3_9333_9071 n3_9333_9104 2.095238e-02
R40657 n3_9333_9104 n3_9333_9287 1.161905e-01
R40658 n3_9333_9287 n3_9333_9320 2.095238e-02
R40659 n3_9333_9320 n3_9333_9424 6.603175e-02
R40660 n3_9333_9424 n3_9333_9503 5.015873e-02
R40661 n3_9333_9503 n3_9333_9520 1.079365e-02
R40662 n3_9333_9520 n3_9333_9536 1.015873e-02
R40663 n3_9333_9536 n3_9333_9719 1.161905e-01
R40664 n3_9333_9719 n3_9333_9752 2.095238e-02
R40665 n3_9333_9752 n3_9333_9935 1.161905e-01
R40666 n3_9333_9935 n3_9333_9968 2.095238e-02
R40667 n3_9333_9968 n3_9333_10151 1.161905e-01
R40668 n3_9333_10151 n3_9333_10184 2.095238e-02
R40669 n3_9333_10184 n3_9333_10367 1.161905e-01
R40670 n3_9333_10367 n3_9333_10400 2.095238e-02
R40671 n3_9333_10799 n3_9333_10832 2.095238e-02
R40672 n3_9333_10832 n3_9333_11015 1.161905e-01
R40673 n3_9333_11015 n3_9333_11048 2.095238e-02
R40674 n3_9333_11048 n3_9333_11231 1.161905e-01
R40675 n3_9333_11231 n3_9333_11264 2.095238e-02
R40676 n3_9333_11264 n3_9333_11447 1.161905e-01
R40677 n3_9333_11447 n3_9333_11480 2.095238e-02
R40678 n3_9333_11480 n3_9333_11663 1.161905e-01
R40679 n3_9333_11663 n3_9333_11674 6.984127e-03
R40680 n3_9333_11674 n3_9333_11696 1.396825e-02
R40681 n3_9333_11696 n3_9333_11770 4.698413e-02
R40682 n3_9333_11770 n3_9333_11879 6.920635e-02
R40683 n3_9333_11879 n3_9333_11912 2.095238e-02
R40684 n3_9333_11912 n3_9333_12095 1.161905e-01
R40685 n3_9333_12095 n3_9333_12128 2.095238e-02
R40686 n3_9333_12128 n3_9333_12311 1.161905e-01
R40687 n3_9333_12311 n3_9333_12344 2.095238e-02
R40688 n3_9333_12344 n3_9333_12527 1.161905e-01
R40689 n3_9333_12527 n3_9333_12560 2.095238e-02
R40690 n3_9333_12560 n3_9333_12743 1.161905e-01
R40691 n3_9333_12959 n3_9333_12992 2.095238e-02
R40692 n3_9333_12992 n3_9333_13175 1.161905e-01
R40693 n3_9333_13175 n3_9333_13208 2.095238e-02
R40694 n3_9333_13208 n3_9333_13391 1.161905e-01
R40695 n3_9333_13391 n3_9333_13424 2.095238e-02
R40696 n3_9333_13424 n3_9333_13607 1.161905e-01
R40697 n3_9333_13607 n3_9333_13640 2.095238e-02
R40698 n3_9333_13640 n3_9333_13796 9.904762e-02
R40699 n3_9333_13796 n3_9333_13823 1.714286e-02
R40700 n3_9333_13823 n3_9333_13856 2.095238e-02
R40701 n3_9333_13856 n3_9333_13924 4.317460e-02
R40702 n3_9333_13924 n3_9333_13990 4.190476e-02
R40703 n3_9333_13990 n3_9333_14012 1.396825e-02
R40704 n3_9333_14012 n3_9333_14020 5.079365e-03
R40705 n3_9333_14020 n3_9333_14039 1.206349e-02
R40706 n3_9333_14039 n3_9333_14072 2.095238e-02
R40707 n3_9333_14072 n3_9333_14228 9.904762e-02
R40708 n3_9333_14228 n3_9333_14255 1.714286e-02
R40709 n3_9333_14255 n3_9333_14288 2.095238e-02
R40710 n3_9333_14288 n3_9333_14471 1.161905e-01
R40711 n3_9333_14471 n3_9333_14504 2.095238e-02
R40712 n3_9333_14504 n3_9333_14660 9.904762e-02
R40713 n3_9333_14660 n3_9333_14687 1.714286e-02
R40714 n3_9333_14687 n3_9333_14720 2.095238e-02
R40715 n3_9333_14720 n3_9333_14903 1.161905e-01
R40716 n3_9333_14903 n3_9333_14936 2.095238e-02
R40717 n3_9333_15335 n3_9333_15368 2.095238e-02
R40718 n3_9333_15368 n3_9333_15551 1.161905e-01
R40719 n3_9333_15551 n3_9333_15584 2.095238e-02
R40720 n3_9333_15584 n3_9333_15740 9.904762e-02
R40721 n3_9333_15740 n3_9333_15767 1.714286e-02
R40722 n3_9333_15767 n3_9333_15800 2.095238e-02
R40723 n3_9333_15800 n3_9333_15934 8.507937e-02
R40724 n3_9333_15934 n3_9333_15956 1.396825e-02
R40725 n3_9333_15956 n3_9333_15983 1.714286e-02
R40726 n3_9333_15983 n3_9333_16016 2.095238e-02
R40727 n3_9333_16016 n3_9333_16172 9.904762e-02
R40728 n3_9333_16172 n3_9333_16174 1.269841e-03
R40729 n3_9333_16174 n3_9333_16199 1.587302e-02
R40730 n3_9333_16199 n3_9333_16232 2.095238e-02
R40731 n3_9333_16232 n3_9333_16270 2.412698e-02
R40732 n3_9333_16270 n3_9333_16415 9.206349e-02
R40733 n3_9333_16415 n3_9333_16448 2.095238e-02
R40734 n3_9333_16448 n3_9333_16631 1.161905e-01
R40735 n3_9333_16631 n3_9333_16664 2.095238e-02
R40736 n3_9333_16664 n3_9333_16847 1.161905e-01
R40737 n3_9333_16847 n3_9333_16880 2.095238e-02
R40738 n3_9333_16880 n3_9333_17063 1.161905e-01
R40739 n3_9333_17063 n3_9333_17096 2.095238e-02
R40740 n3_9333_17096 n3_9333_17230 8.507937e-02
R40741 n3_9333_17468 n3_9333_17495 1.714286e-02
R40742 n3_9333_17495 n3_9333_17528 2.095238e-02
R40743 n3_9333_17528 n3_9333_17711 1.161905e-01
R40744 n3_9333_17711 n3_9333_17744 2.095238e-02
R40745 n3_9333_17744 n3_9333_17927 1.161905e-01
R40746 n3_9333_17927 n3_9333_17960 2.095238e-02
R40747 n3_9333_17960 n3_9333_18143 1.161905e-01
R40748 n3_9333_18143 n3_9333_18176 2.095238e-02
R40749 n3_9333_18176 n3_9333_18359 1.161905e-01
R40750 n3_9333_18359 n3_9333_18392 2.095238e-02
R40751 n3_9333_18392 n3_9333_18424 2.031746e-02
R40752 n3_9333_18424 n3_9333_18520 6.095238e-02
R40753 n3_9333_18520 n3_9333_18527 4.444444e-03
R40754 n3_9333_18527 n3_9333_18548 1.333333e-02
R40755 n3_9333_18548 n3_9333_18575 1.714286e-02
R40756 n3_9333_18575 n3_9333_18608 2.095238e-02
R40757 n3_9333_18608 n3_9333_18764 9.904762e-02
R40758 n3_9333_18764 n3_9333_18791 1.714286e-02
R40759 n3_9333_18791 n3_9333_18824 2.095238e-02
R40760 n3_9333_18824 n3_9333_19007 1.161905e-01
R40761 n3_9333_19007 n3_9333_19040 2.095238e-02
R40762 n3_9333_19040 n3_9333_19223 1.161905e-01
R40763 n3_9333_19223 n3_9333_19256 2.095238e-02
R40764 n3_9333_19256 n3_9333_19412 9.904762e-02
R40765 n3_9333_19412 n3_9333_19439 1.714286e-02
R40766 n3_9333_19439 n3_9333_19472 2.095238e-02
R40767 n3_9333_19871 n3_9333_19904 2.095238e-02
R40768 n3_9333_19904 n3_9333_20087 1.161905e-01
R40769 n3_9333_20087 n3_9333_20120 2.095238e-02
R40770 n3_9333_20120 n3_9333_20303 1.161905e-01
R40771 n3_9333_20303 n3_9333_20336 2.095238e-02
R40772 n3_9333_20336 n3_9333_20519 1.161905e-01
R40773 n3_9333_20519 n3_9333_20552 2.095238e-02
R40774 n3_9333_20552 n3_9333_20674 7.746032e-02
R40775 n3_9333_20674 n3_9333_20687 8.253968e-03
R40776 n3_9333_20687 n3_9333_20735 3.047619e-02
R40777 n3_9333_20735 n3_9333_20768 2.095238e-02
R40778 n3_9333_20768 n3_9333_20770 1.269841e-03
R40779 n3_9333_20770 n3_9333_20951 1.149206e-01
R40780 n3_9333_20951 n3_9333_20984 2.095238e-02
R40781 n3_9521_215 n3_9521_248 2.095238e-02
R40782 n3_9521_248 n3_9521_383 8.571429e-02
R40783 n3_9521_383 n3_9521_424 2.603175e-02
R40784 n3_9521_424 n3_9521_431 4.444444e-03
R40785 n3_9521_520 n3_9521_647 8.063492e-02
R40786 n3_9521_647 n3_9521_680 2.095238e-02
R40787 n3_9521_680 n3_9521_863 1.161905e-01
R40788 n3_9521_863 n3_9521_896 2.095238e-02
R40789 n3_9521_896 n3_9521_1079 1.161905e-01
R40790 n3_9521_1079 n3_9521_1112 2.095238e-02
R40791 n3_9521_1112 n3_9521_1295 1.161905e-01
R40792 n3_9521_1295 n3_9521_1328 2.095238e-02
R40793 n3_9521_1328 n3_9521_1511 1.161905e-01
R40794 n3_9521_1511 n3_9521_1544 2.095238e-02
R40795 n3_9521_1544 n3_9521_1727 1.161905e-01
R40796 n3_9521_1727 n3_9521_1760 2.095238e-02
R40797 n3_9521_1760 n3_9521_1894 8.507937e-02
R40798 n3_9521_1894 n3_9521_1916 1.396825e-02
R40799 n3_9521_1916 n3_9521_1943 1.714286e-02
R40800 n3_9521_1943 n3_9521_1976 2.095238e-02
R40801 n3_9521_1976 n3_9521_2159 1.161905e-01
R40802 n3_9521_2159 n3_9521_2192 2.095238e-02
R40803 n3_9521_2192 n3_9521_2375 1.161905e-01
R40804 n3_9521_2375 n3_9521_2408 2.095238e-02
R40805 n3_9521_2408 n3_9521_2543 8.571429e-02
R40806 n3_9521_2543 n3_9521_2564 1.333333e-02
R40807 n3_9521_2564 n3_9521_2591 1.714286e-02
R40808 n3_9521_2591 n3_9521_2624 2.095238e-02
R40809 n3_9521_2624 n3_9521_2674 3.174603e-02
R40810 n3_9521_2770 n3_9521_2807 2.349206e-02
R40811 n3_9521_2807 n3_9521_2840 2.095238e-02
R40812 n3_9521_2840 n3_9521_2996 9.904762e-02
R40813 n3_9521_2996 n3_9521_3023 1.714286e-02
R40814 n3_9521_3023 n3_9521_3056 2.095238e-02
R40815 n3_9521_3056 n3_9521_3239 1.161905e-01
R40816 n3_9521_3239 n3_9521_3272 2.095238e-02
R40817 n3_9521_3272 n3_9521_3455 1.161905e-01
R40818 n3_9521_3455 n3_9521_3488 2.095238e-02
R40819 n3_9521_3488 n3_9521_3644 9.904762e-02
R40820 n3_9521_3644 n3_9521_3671 1.714286e-02
R40821 n3_9521_3671 n3_9521_3704 2.095238e-02
R40822 n3_9521_3704 n3_9521_3887 1.161905e-01
R40823 n3_9521_3887 n3_9521_3920 2.095238e-02
R40824 n3_9521_3920 n3_9521_4103 1.161905e-01
R40825 n3_9521_4103 n3_9521_4136 2.095238e-02
R40826 n3_9521_4136 n3_9521_4292 9.904762e-02
R40827 n3_9521_4292 n3_9521_4319 1.714286e-02
R40828 n3_9521_4319 n3_9521_4352 2.095238e-02
R40829 n3_9521_4352 n3_9521_4535 1.161905e-01
R40830 n3_9521_4535 n3_9521_4568 2.095238e-02
R40831 n3_9521_4568 n3_9521_4724 9.904762e-02
R40832 n3_9521_4724 n3_9521_4751 1.714286e-02
R40833 n3_9521_4751 n3_9521_4784 2.095238e-02
R40834 n3_9521_4784 n3_9521_4924 8.888889e-02
R40835 n3_9521_5000 n3_9521_5020 1.269841e-02
R40836 n3_9521_5020 n3_9521_5183 1.034921e-01
R40837 n3_9521_5183 n3_9521_5216 2.095238e-02
R40838 n3_9521_5216 n3_9521_5350 8.507937e-02
R40839 n3_9521_5350 n3_9521_5372 1.396825e-02
R40840 n3_9521_5372 n3_9521_5399 1.714286e-02
R40841 n3_9521_5399 n3_9521_5432 2.095238e-02
R40842 n3_9521_5432 n3_9521_5588 9.904762e-02
R40843 n3_9521_5588 n3_9521_5615 1.714286e-02
R40844 n3_9521_5615 n3_9521_5648 2.095238e-02
R40845 n3_9521_5648 n3_9521_5831 1.161905e-01
R40846 n3_9521_5831 n3_9521_5864 2.095238e-02
R40847 n3_9521_5864 n3_9521_6047 1.161905e-01
R40848 n3_9521_6047 n3_9521_6080 2.095238e-02
R40849 n3_9521_6080 n3_9521_6263 1.161905e-01
R40850 n3_9521_6263 n3_9521_6296 2.095238e-02
R40851 n3_9521_6296 n3_9521_6479 1.161905e-01
R40852 n3_9521_6479 n3_9521_6512 2.095238e-02
R40853 n3_9521_6512 n3_9521_6668 9.904762e-02
R40854 n3_9521_6668 n3_9521_6695 1.714286e-02
R40855 n3_9521_6695 n3_9521_6728 2.095238e-02
R40856 n3_9521_6728 n3_9521_6911 1.161905e-01
R40857 n3_9521_6911 n3_9521_6944 2.095238e-02
R40858 n3_9521_6944 n3_9521_7100 9.904762e-02
R40859 n3_9521_7100 n3_9521_7127 1.714286e-02
R40860 n3_9521_7127 n3_9521_7160 2.095238e-02
R40861 n3_9521_7160 n3_9521_7174 8.888889e-03
R40862 n3_9521_7270 n3_9521_7316 2.920635e-02
R40863 n3_9521_7316 n3_9521_7343 1.714286e-02
R40864 n3_9521_7343 n3_9521_7376 2.095238e-02
R40865 n3_9521_7376 n3_9521_7532 9.904762e-02
R40866 n3_9521_7532 n3_9521_7559 1.714286e-02
R40867 n3_9521_7559 n3_9521_7592 2.095238e-02
R40868 n3_9521_7592 n3_9521_7775 1.161905e-01
R40869 n3_9521_7775 n3_9521_7808 2.095238e-02
R40870 n3_9521_7808 n3_9521_7991 1.161905e-01
R40871 n3_9521_7991 n3_9521_8024 2.095238e-02
R40872 n3_9521_8024 n3_9521_8207 1.161905e-01
R40873 n3_9521_8207 n3_9521_8240 2.095238e-02
R40874 n3_9521_8240 n3_9521_8423 1.161905e-01
R40875 n3_9521_8423 n3_9521_8456 2.095238e-02
R40876 n3_9521_8456 n3_9521_8639 1.161905e-01
R40877 n3_9521_8639 n3_9521_8672 2.095238e-02
R40878 n3_9521_8672 n3_9521_8855 1.161905e-01
R40879 n3_9521_8855 n3_9521_8888 2.095238e-02
R40880 n3_9521_8888 n3_9521_9071 1.161905e-01
R40881 n3_9521_9071 n3_9521_9104 2.095238e-02
R40882 n3_9521_9104 n3_9521_9287 1.161905e-01
R40883 n3_9521_9287 n3_9521_9320 2.095238e-02
R40884 n3_9521_9320 n3_9521_9424 6.603175e-02
R40885 n3_9521_9503 n3_9521_9520 1.079365e-02
R40886 n3_9521_9520 n3_9521_9536 1.015873e-02
R40887 n3_9521_9536 n3_9521_9719 1.161905e-01
R40888 n3_9521_9719 n3_9521_9752 2.095238e-02
R40889 n3_9521_9752 n3_9521_9935 1.161905e-01
R40890 n3_9521_9935 n3_9521_9968 2.095238e-02
R40891 n3_9521_9968 n3_9521_10151 1.161905e-01
R40892 n3_9521_10151 n3_9521_10184 2.095238e-02
R40893 n3_9521_10184 n3_9521_10367 1.161905e-01
R40894 n3_9521_10367 n3_9521_10400 2.095238e-02
R40895 n3_9521_10616 n3_9521_10799 1.161905e-01
R40896 n3_9521_10799 n3_9521_10832 2.095238e-02
R40897 n3_9521_10832 n3_9521_11015 1.161905e-01
R40898 n3_9521_11015 n3_9521_11048 2.095238e-02
R40899 n3_9521_11048 n3_9521_11231 1.161905e-01
R40900 n3_9521_11231 n3_9521_11264 2.095238e-02
R40901 n3_9521_11264 n3_9521_11447 1.161905e-01
R40902 n3_9521_11447 n3_9521_11480 2.095238e-02
R40903 n3_9521_11480 n3_9521_11663 1.161905e-01
R40904 n3_9521_11663 n3_9521_11674 6.984127e-03
R40905 n3_9521_11674 n3_9521_11696 1.396825e-02
R40906 n3_9521_11770 n3_9521_11879 6.920635e-02
R40907 n3_9521_11879 n3_9521_11912 2.095238e-02
R40908 n3_9521_11912 n3_9521_12095 1.161905e-01
R40909 n3_9521_12095 n3_9521_12128 2.095238e-02
R40910 n3_9521_12128 n3_9521_12311 1.161905e-01
R40911 n3_9521_12311 n3_9521_12344 2.095238e-02
R40912 n3_9521_12344 n3_9521_12527 1.161905e-01
R40913 n3_9521_12527 n3_9521_12560 2.095238e-02
R40914 n3_9521_12560 n3_9521_12743 1.161905e-01
R40915 n3_9521_12743 n3_9521_12776 2.095238e-02
R40916 n3_9521_12776 n3_9521_12959 1.161905e-01
R40917 n3_9521_12959 n3_9521_12992 2.095238e-02
R40918 n3_9521_12992 n3_9521_13175 1.161905e-01
R40919 n3_9521_13175 n3_9521_13208 2.095238e-02
R40920 n3_9521_13208 n3_9521_13391 1.161905e-01
R40921 n3_9521_13391 n3_9521_13424 2.095238e-02
R40922 n3_9521_13424 n3_9521_13607 1.161905e-01
R40923 n3_9521_13607 n3_9521_13640 2.095238e-02
R40924 n3_9521_13640 n3_9521_13796 9.904762e-02
R40925 n3_9521_13796 n3_9521_13823 1.714286e-02
R40926 n3_9521_13823 n3_9521_13856 2.095238e-02
R40927 n3_9521_13856 n3_9521_13924 4.317460e-02
R40928 n3_9521_13990 n3_9521_14012 1.396825e-02
R40929 n3_9521_14012 n3_9521_14020 5.079365e-03
R40930 n3_9521_14020 n3_9521_14039 1.206349e-02
R40931 n3_9521_14039 n3_9521_14072 2.095238e-02
R40932 n3_9521_14072 n3_9521_14228 9.904762e-02
R40933 n3_9521_14228 n3_9521_14255 1.714286e-02
R40934 n3_9521_14255 n3_9521_14288 2.095238e-02
R40935 n3_9521_14288 n3_9521_14471 1.161905e-01
R40936 n3_9521_14471 n3_9521_14504 2.095238e-02
R40937 n3_9521_14504 n3_9521_14660 9.904762e-02
R40938 n3_9521_14660 n3_9521_14687 1.714286e-02
R40939 n3_9521_14687 n3_9521_14720 2.095238e-02
R40940 n3_9521_14720 n3_9521_14903 1.161905e-01
R40941 n3_9521_14903 n3_9521_14936 2.095238e-02
R40942 n3_9521_14936 n3_9521_15119 1.161905e-01
R40943 n3_9521_15119 n3_9521_15152 2.095238e-02
R40944 n3_9521_15152 n3_9521_15335 1.161905e-01
R40945 n3_9521_15335 n3_9521_15368 2.095238e-02
R40946 n3_9521_15368 n3_9521_15551 1.161905e-01
R40947 n3_9521_15551 n3_9521_15584 2.095238e-02
R40948 n3_9521_15584 n3_9521_15740 9.904762e-02
R40949 n3_9521_15740 n3_9521_15767 1.714286e-02
R40950 n3_9521_15767 n3_9521_15800 2.095238e-02
R40951 n3_9521_15800 n3_9521_15934 8.507937e-02
R40952 n3_9521_15934 n3_9521_15956 1.396825e-02
R40953 n3_9521_15956 n3_9521_15983 1.714286e-02
R40954 n3_9521_15983 n3_9521_16016 2.095238e-02
R40955 n3_9521_16016 n3_9521_16172 9.904762e-02
R40956 n3_9521_16172 n3_9521_16174 1.269841e-03
R40957 n3_9521_16174 n3_9521_16199 1.587302e-02
R40958 n3_9521_16270 n3_9521_16415 9.206349e-02
R40959 n3_9521_16415 n3_9521_16448 2.095238e-02
R40960 n3_9521_16448 n3_9521_16631 1.161905e-01
R40961 n3_9521_16631 n3_9521_16664 2.095238e-02
R40962 n3_9521_16664 n3_9521_16847 1.161905e-01
R40963 n3_9521_16847 n3_9521_16880 2.095238e-02
R40964 n3_9521_16880 n3_9521_17063 1.161905e-01
R40965 n3_9521_17063 n3_9521_17096 2.095238e-02
R40966 n3_9521_17096 n3_9521_17230 8.507937e-02
R40967 n3_9521_17230 n3_9521_17252 1.396825e-02
R40968 n3_9521_17252 n3_9521_17279 1.714286e-02
R40969 n3_9521_17279 n3_9521_17312 2.095238e-02
R40970 n3_9521_17312 n3_9521_17468 9.904762e-02
R40971 n3_9521_17468 n3_9521_17495 1.714286e-02
R40972 n3_9521_17495 n3_9521_17528 2.095238e-02
R40973 n3_9521_17528 n3_9521_17711 1.161905e-01
R40974 n3_9521_17711 n3_9521_17744 2.095238e-02
R40975 n3_9521_17744 n3_9521_17927 1.161905e-01
R40976 n3_9521_17927 n3_9521_17960 2.095238e-02
R40977 n3_9521_17960 n3_9521_18143 1.161905e-01
R40978 n3_9521_18143 n3_9521_18176 2.095238e-02
R40979 n3_9521_18176 n3_9521_18359 1.161905e-01
R40980 n3_9521_18359 n3_9521_18392 2.095238e-02
R40981 n3_9521_18392 n3_9521_18424 2.031746e-02
R40982 n3_9521_18520 n3_9521_18527 4.444444e-03
R40983 n3_9521_18527 n3_9521_18548 1.333333e-02
R40984 n3_9521_18548 n3_9521_18575 1.714286e-02
R40985 n3_9521_18575 n3_9521_18608 2.095238e-02
R40986 n3_9521_18608 n3_9521_18764 9.904762e-02
R40987 n3_9521_18764 n3_9521_18791 1.714286e-02
R40988 n3_9521_18791 n3_9521_18824 2.095238e-02
R40989 n3_9521_18824 n3_9521_19007 1.161905e-01
R40990 n3_9521_19007 n3_9521_19040 2.095238e-02
R40991 n3_9521_19040 n3_9521_19223 1.161905e-01
R40992 n3_9521_19223 n3_9521_19256 2.095238e-02
R40993 n3_9521_19256 n3_9521_19412 9.904762e-02
R40994 n3_9521_19412 n3_9521_19439 1.714286e-02
R40995 n3_9521_19439 n3_9521_19472 2.095238e-02
R40996 n3_9521_19472 n3_9521_19655 1.161905e-01
R40997 n3_9521_19655 n3_9521_19688 2.095238e-02
R40998 n3_9521_19688 n3_9521_19871 1.161905e-01
R40999 n3_9521_19871 n3_9521_19904 2.095238e-02
R41000 n3_9521_19904 n3_9521_20087 1.161905e-01
R41001 n3_9521_20087 n3_9521_20120 2.095238e-02
R41002 n3_9521_20120 n3_9521_20303 1.161905e-01
R41003 n3_9521_20303 n3_9521_20336 2.095238e-02
R41004 n3_9521_20336 n3_9521_20519 1.161905e-01
R41005 n3_9521_20519 n3_9521_20552 2.095238e-02
R41006 n3_9521_20552 n3_9521_20674 7.746032e-02
R41007 n3_9521_20674 n3_9521_20687 8.253968e-03
R41008 n3_9521_20768 n3_9521_20770 1.269841e-03
R41009 n3_9521_20770 n3_9521_20951 1.149206e-01
R41010 n3_9521_20951 n3_9521_20984 2.095238e-02
R41011 n3_9614_215 n3_9614_248 2.095238e-02
R41012 n3_9614_248 n3_9614_383 8.571429e-02
R41013 n3_9614_383 n3_9614_431 3.047619e-02
R41014 n3_9614_431 n3_9614_464 2.095238e-02
R41015 n3_9614_464 n3_9614_647 1.161905e-01
R41016 n3_9614_647 n3_9614_680 2.095238e-02
R41017 n3_9614_680 n3_9614_863 1.161905e-01
R41018 n3_9614_863 n3_9614_896 2.095238e-02
R41019 n3_9614_896 n3_9614_1079 1.161905e-01
R41020 n3_9614_1079 n3_9614_1112 2.095238e-02
R41021 n3_9614_1112 n3_9614_1295 1.161905e-01
R41022 n3_9614_1295 n3_9614_1328 2.095238e-02
R41023 n3_9614_1328 n3_9614_1511 1.161905e-01
R41024 n3_9614_1511 n3_9614_1544 2.095238e-02
R41025 n3_9614_1544 n3_9614_1727 1.161905e-01
R41026 n3_9614_1727 n3_9614_1760 2.095238e-02
R41027 n3_9614_1760 n3_9614_1916 9.904762e-02
R41028 n3_9614_1916 n3_9614_1943 1.714286e-02
R41029 n3_9614_1943 n3_9614_1976 2.095238e-02
R41030 n3_9614_1976 n3_9614_2159 1.161905e-01
R41031 n3_9614_2159 n3_9614_2192 2.095238e-02
R41032 n3_9614_2192 n3_9614_2375 1.161905e-01
R41033 n3_9614_2375 n3_9614_2408 2.095238e-02
R41034 n3_9614_2408 n3_9614_2543 8.571429e-02
R41035 n3_9614_2543 n3_9614_2564 1.333333e-02
R41036 n3_9614_2564 n3_9614_2591 1.714286e-02
R41037 n3_9614_2591 n3_9614_2624 2.095238e-02
R41038 n3_9614_18527 n3_9614_18548 1.333333e-02
R41039 n3_9614_18548 n3_9614_18575 1.714286e-02
R41040 n3_9614_18575 n3_9614_18608 2.095238e-02
R41041 n3_9614_18608 n3_9614_18764 9.904762e-02
R41042 n3_9614_18764 n3_9614_18791 1.714286e-02
R41043 n3_9614_18791 n3_9614_18824 2.095238e-02
R41044 n3_9614_18824 n3_9614_19007 1.161905e-01
R41045 n3_9614_19007 n3_9614_19040 2.095238e-02
R41046 n3_9614_19040 n3_9614_19223 1.161905e-01
R41047 n3_9614_19223 n3_9614_19256 2.095238e-02
R41048 n3_9614_19256 n3_9614_19412 9.904762e-02
R41049 n3_9614_19412 n3_9614_19439 1.714286e-02
R41050 n3_9614_19439 n3_9614_19472 2.095238e-02
R41051 n3_9614_19472 n3_9614_19655 1.161905e-01
R41052 n3_9614_19655 n3_9614_19688 2.095238e-02
R41053 n3_9614_19688 n3_9614_19871 1.161905e-01
R41054 n3_9614_19871 n3_9614_19904 2.095238e-02
R41055 n3_9614_19904 n3_9614_20087 1.161905e-01
R41056 n3_9614_20087 n3_9614_20120 2.095238e-02
R41057 n3_9614_20120 n3_9614_20303 1.161905e-01
R41058 n3_9614_20303 n3_9614_20336 2.095238e-02
R41059 n3_9614_20336 n3_9614_20519 1.161905e-01
R41060 n3_9614_20519 n3_9614_20552 2.095238e-02
R41061 n3_9614_20552 n3_9614_20687 8.571429e-02
R41062 n3_9614_20687 n3_9614_20735 3.047619e-02
R41063 n3_9614_20735 n3_9614_20768 2.095238e-02
R41064 n3_9614_20768 n3_9614_20951 1.161905e-01
R41065 n3_9614_20951 n3_9614_20984 2.095238e-02
R41066 n3_11400_215 n3_11400_248 2.095238e-02
R41067 n3_11400_248 n3_11400_383 8.571429e-02
R41068 n3_11400_383 n3_11400_431 3.047619e-02
R41069 n3_11400_431 n3_11400_464 2.095238e-02
R41070 n3_11400_464 n3_11400_647 1.161905e-01
R41071 n3_11400_647 n3_11400_680 2.095238e-02
R41072 n3_11400_680 n3_11400_863 1.161905e-01
R41073 n3_11400_863 n3_11400_896 2.095238e-02
R41074 n3_11400_896 n3_11400_1079 1.161905e-01
R41075 n3_11400_1079 n3_11400_1112 2.095238e-02
R41076 n3_11400_1112 n3_11400_1295 1.161905e-01
R41077 n3_11400_1295 n3_11400_1328 2.095238e-02
R41078 n3_11400_1328 n3_11400_1511 1.161905e-01
R41079 n3_11400_1511 n3_11400_1544 2.095238e-02
R41080 n3_11400_1544 n3_11400_1727 1.161905e-01
R41081 n3_11400_1727 n3_11400_1760 2.095238e-02
R41082 n3_11400_1760 n3_11400_1894 8.507937e-02
R41083 n3_11400_1894 n3_11400_1943 3.111111e-02
R41084 n3_11400_1943 n3_11400_1976 2.095238e-02
R41085 n3_11400_1976 n3_11400_2159 1.161905e-01
R41086 n3_11400_2159 n3_11400_2192 2.095238e-02
R41087 n3_11400_2192 n3_11400_2375 1.161905e-01
R41088 n3_11400_2375 n3_11400_2408 2.095238e-02
R41089 n3_11400_2408 n3_11400_2543 8.571429e-02
R41090 n3_11400_2543 n3_11400_2591 3.047619e-02
R41091 n3_11400_2591 n3_11400_2624 2.095238e-02
R41092 n3_11400_18527 n3_11400_18548 1.333333e-02
R41093 n3_11400_18548 n3_11400_18575 1.714286e-02
R41094 n3_11400_18575 n3_11400_18608 2.095238e-02
R41095 n3_11400_18608 n3_11400_18764 9.904762e-02
R41096 n3_11400_18764 n3_11400_18791 1.714286e-02
R41097 n3_11400_18791 n3_11400_18824 2.095238e-02
R41098 n3_11400_18824 n3_11400_19007 1.161905e-01
R41099 n3_11400_19007 n3_11400_19040 2.095238e-02
R41100 n3_11400_19040 n3_11400_19223 1.161905e-01
R41101 n3_11400_19223 n3_11400_19256 2.095238e-02
R41102 n3_11400_19256 n3_11400_19412 9.904762e-02
R41103 n3_11400_19412 n3_11400_19439 1.714286e-02
R41104 n3_11400_19439 n3_11400_19472 2.095238e-02
R41105 n3_11400_19472 n3_11400_19655 1.161905e-01
R41106 n3_11400_19655 n3_11400_19688 2.095238e-02
R41107 n3_11400_19688 n3_11400_19871 1.161905e-01
R41108 n3_11400_19871 n3_11400_19904 2.095238e-02
R41109 n3_11400_19904 n3_11400_20087 1.161905e-01
R41110 n3_11400_20087 n3_11400_20120 2.095238e-02
R41111 n3_11400_20120 n3_11400_20303 1.161905e-01
R41112 n3_11400_20303 n3_11400_20336 2.095238e-02
R41113 n3_11400_20336 n3_11400_20519 1.161905e-01
R41114 n3_11400_20519 n3_11400_20552 2.095238e-02
R41115 n3_11400_20552 n3_11400_20687 8.571429e-02
R41116 n3_11400_20687 n3_11400_20735 3.047619e-02
R41117 n3_11400_20735 n3_11400_20768 2.095238e-02
R41118 n3_11400_20768 n3_11400_20951 1.161905e-01
R41119 n3_11400_20951 n3_11400_20984 2.095238e-02
R41120 n3_11583_424 n3_11630_424 2.984127e-02
R41121 n3_11630_424 n3_11771_424 8.952381e-02
R41122 n3_11583_520 n3_11630_520 2.984127e-02
R41123 n3_11630_520 n3_11771_520 8.952381e-02
R41124 n3_11583_2674 n3_11630_2674 2.984127e-02
R41125 n3_11630_2674 n3_11771_2674 8.952381e-02
R41126 n3_11583_2770 n3_11630_2770 2.984127e-02
R41127 n3_11630_2770 n3_11771_2770 8.952381e-02
R41128 n3_11583_4924 n3_11630_4924 2.984127e-02
R41129 n3_11630_4924 n3_11771_4924 8.952381e-02
R41130 n3_11583_5020 n3_11630_5020 2.984127e-02
R41131 n3_11630_5020 n3_11771_5020 8.952381e-02
R41132 n3_11583_7174 n3_11630_7174 2.984127e-02
R41133 n3_11630_7174 n3_11771_7174 8.952381e-02
R41134 n3_11583_7270 n3_11630_7270 2.984127e-02
R41135 n3_11630_7270 n3_11771_7270 8.952381e-02
R41136 n3_11583_9424 n3_11630_9424 2.984127e-02
R41137 n3_11630_9424 n3_11771_9424 8.952381e-02
R41138 n3_11583_9520 n3_11630_9520 2.984127e-02
R41139 n3_11630_9520 n3_11771_9520 8.952381e-02
R41140 n3_11583_11674 n3_11630_11674 2.984127e-02
R41141 n3_11630_11674 n3_11771_11674 8.952381e-02
R41142 n3_11583_11770 n3_11630_11770 2.984127e-02
R41143 n3_11630_11770 n3_11771_11770 8.952381e-02
R41144 n3_11583_13924 n3_11630_13924 2.984127e-02
R41145 n3_11630_13924 n3_11771_13924 8.952381e-02
R41146 n3_11583_14020 n3_11630_14020 2.984127e-02
R41147 n3_11630_14020 n3_11771_14020 8.952381e-02
R41148 n3_11583_16174 n3_11630_16174 2.984127e-02
R41149 n3_11630_16174 n3_11771_16174 8.952381e-02
R41150 n3_11583_16270 n3_11630_16270 2.984127e-02
R41151 n3_11630_16270 n3_11771_16270 8.952381e-02
R41152 n3_11583_18424 n3_11630_18424 2.984127e-02
R41153 n3_11630_18424 n3_11771_18424 8.952381e-02
R41154 n3_11583_18520 n3_11630_18520 2.984127e-02
R41155 n3_11630_18520 n3_11771_18520 8.952381e-02
R41156 n3_11583_20674 n3_11630_20674 2.984127e-02
R41157 n3_11630_20674 n3_11771_20674 8.952381e-02
R41158 n3_11583_20770 n3_11630_20770 2.984127e-02
R41159 n3_11630_20770 n3_11771_20770 8.952381e-02
R41160 n3_11583_215 n3_11583_248 2.095238e-02
R41161 n3_11583_248 n3_11583_383 8.571429e-02
R41162 n3_11583_383 n3_11583_424 2.603175e-02
R41163 n3_11583_424 n3_11583_431 4.444444e-03
R41164 n3_11583_431 n3_11583_464 2.095238e-02
R41165 n3_11583_464 n3_11583_520 3.555556e-02
R41166 n3_11583_520 n3_11583_647 8.063492e-02
R41167 n3_11583_647 n3_11583_680 2.095238e-02
R41168 n3_11583_680 n3_11583_863 1.161905e-01
R41169 n3_11583_863 n3_11583_896 2.095238e-02
R41170 n3_11583_896 n3_11583_1079 1.161905e-01
R41171 n3_11583_1079 n3_11583_1112 2.095238e-02
R41172 n3_11583_1112 n3_11583_1295 1.161905e-01
R41173 n3_11583_1295 n3_11583_1328 2.095238e-02
R41174 n3_11583_1727 n3_11583_1760 2.095238e-02
R41175 n3_11583_1760 n3_11583_1894 8.507937e-02
R41176 n3_11583_1894 n3_11583_1943 3.111111e-02
R41177 n3_11583_1943 n3_11583_1976 2.095238e-02
R41178 n3_11583_1976 n3_11583_2159 1.161905e-01
R41179 n3_11583_2159 n3_11583_2192 2.095238e-02
R41180 n3_11583_2192 n3_11583_2375 1.161905e-01
R41181 n3_11583_2375 n3_11583_2408 2.095238e-02
R41182 n3_11583_2408 n3_11583_2542 8.507937e-02
R41183 n3_11583_2542 n3_11583_2543 6.349206e-04
R41184 n3_11583_2543 n3_11583_2591 3.047619e-02
R41185 n3_11583_2591 n3_11583_2624 2.095238e-02
R41186 n3_11583_2624 n3_11583_2674 3.174603e-02
R41187 n3_11583_2674 n3_11583_2760 5.460317e-02
R41188 n3_11583_2760 n3_11583_2770 6.349206e-03
R41189 n3_11583_2770 n3_11583_2807 2.349206e-02
R41190 n3_11583_2807 n3_11583_2840 2.095238e-02
R41191 n3_11583_2840 n3_11583_2974 8.507937e-02
R41192 n3_11583_2974 n3_11583_3023 3.111111e-02
R41193 n3_11583_3023 n3_11583_3056 2.095238e-02
R41194 n3_11583_3056 n3_11583_3239 1.161905e-01
R41195 n3_11583_3239 n3_11583_3272 2.095238e-02
R41196 n3_11583_3272 n3_11583_3455 1.161905e-01
R41197 n3_11583_3455 n3_11583_3488 2.095238e-02
R41198 n3_11583_3488 n3_11583_3622 8.507937e-02
R41199 n3_11583_3622 n3_11583_3671 3.111111e-02
R41200 n3_11583_3671 n3_11583_3704 2.095238e-02
R41201 n3_11583_4103 n3_11583_4136 2.095238e-02
R41202 n3_11583_4136 n3_11583_4270 8.507937e-02
R41203 n3_11583_4270 n3_11583_4319 3.111111e-02
R41204 n3_11583_4319 n3_11583_4352 2.095238e-02
R41205 n3_11583_4352 n3_11583_4535 1.161905e-01
R41206 n3_11583_4535 n3_11583_4568 2.095238e-02
R41207 n3_11583_4568 n3_11583_4702 8.507937e-02
R41208 n3_11583_4702 n3_11583_4751 3.111111e-02
R41209 n3_11583_4751 n3_11583_4784 2.095238e-02
R41210 n3_11583_4784 n3_11583_4924 8.888889e-02
R41211 n3_11583_4924 n3_11583_4967 2.730159e-02
R41212 n3_11583_4967 n3_11583_5000 2.095238e-02
R41213 n3_11583_5000 n3_11583_5020 1.269841e-02
R41214 n3_11583_5020 n3_11583_5183 1.034921e-01
R41215 n3_11583_5183 n3_11583_5216 2.095238e-02
R41216 n3_11583_5216 n3_11583_5350 8.507937e-02
R41217 n3_11583_5350 n3_11583_5399 3.111111e-02
R41218 n3_11583_5399 n3_11583_5432 2.095238e-02
R41219 n3_11583_5432 n3_11583_5566 8.507937e-02
R41220 n3_11583_5566 n3_11583_5615 3.111111e-02
R41221 n3_11583_5615 n3_11583_5648 2.095238e-02
R41222 n3_11583_5648 n3_11583_5782 8.507937e-02
R41223 n3_11583_5782 n3_11583_5831 3.111111e-02
R41224 n3_11583_5831 n3_11583_5864 2.095238e-02
R41225 n3_11583_6263 n3_11583_6296 2.095238e-02
R41226 n3_11583_6296 n3_11583_6430 8.507937e-02
R41227 n3_11583_6430 n3_11583_6479 3.111111e-02
R41228 n3_11583_6479 n3_11583_6512 2.095238e-02
R41229 n3_11583_6512 n3_11583_6646 8.507937e-02
R41230 n3_11583_6646 n3_11583_6695 3.111111e-02
R41231 n3_11583_6695 n3_11583_6728 2.095238e-02
R41232 n3_11583_6728 n3_11583_6862 8.507937e-02
R41233 n3_11583_6862 n3_11583_6911 3.111111e-02
R41234 n3_11583_6911 n3_11583_6944 2.095238e-02
R41235 n3_11583_6944 n3_11583_7078 8.507937e-02
R41236 n3_11583_7078 n3_11583_7127 3.111111e-02
R41237 n3_11583_7127 n3_11583_7160 2.095238e-02
R41238 n3_11583_7160 n3_11583_7174 8.888889e-03
R41239 n3_11583_7174 n3_11583_7270 6.095238e-02
R41240 n3_11583_7270 n3_11583_7294 1.523810e-02
R41241 n3_11583_7294 n3_11583_7343 3.111111e-02
R41242 n3_11583_7343 n3_11583_7376 2.095238e-02
R41243 n3_11583_7376 n3_11583_7510 8.507937e-02
R41244 n3_11583_7510 n3_11583_7559 3.111111e-02
R41245 n3_11583_7559 n3_11583_7592 2.095238e-02
R41246 n3_11583_7592 n3_11583_7775 1.161905e-01
R41247 n3_11583_7775 n3_11583_7808 2.095238e-02
R41248 n3_11583_7808 n3_11583_7991 1.161905e-01
R41249 n3_11583_7991 n3_11583_8024 2.095238e-02
R41250 n3_11583_8024 n3_11583_8207 1.161905e-01
R41251 n3_11583_8207 n3_11583_8240 2.095238e-02
R41252 n3_11583_8456 n3_11583_8639 1.161905e-01
R41253 n3_11583_8639 n3_11583_8672 2.095238e-02
R41254 n3_11583_8672 n3_11583_8855 1.161905e-01
R41255 n3_11583_8855 n3_11583_8888 2.095238e-02
R41256 n3_11583_8888 n3_11583_9071 1.161905e-01
R41257 n3_11583_9071 n3_11583_9104 2.095238e-02
R41258 n3_11583_9104 n3_11583_9287 1.161905e-01
R41259 n3_11583_9287 n3_11583_9320 2.095238e-02
R41260 n3_11583_9320 n3_11583_9424 6.603175e-02
R41261 n3_11583_9424 n3_11583_9503 5.015873e-02
R41262 n3_11583_9503 n3_11583_9520 1.079365e-02
R41263 n3_11583_9520 n3_11583_9536 1.015873e-02
R41264 n3_11583_9536 n3_11583_9719 1.161905e-01
R41265 n3_11583_9719 n3_11583_9752 2.095238e-02
R41266 n3_11583_9752 n3_11583_9935 1.161905e-01
R41267 n3_11583_9935 n3_11583_9968 2.095238e-02
R41268 n3_11583_9968 n3_11583_10151 1.161905e-01
R41269 n3_11583_10151 n3_11583_10184 2.095238e-02
R41270 n3_11583_10184 n3_11583_10367 1.161905e-01
R41271 n3_11583_10367 n3_11583_10400 2.095238e-02
R41272 n3_11583_10799 n3_11583_10832 2.095238e-02
R41273 n3_11583_10832 n3_11583_11015 1.161905e-01
R41274 n3_11583_11015 n3_11583_11048 2.095238e-02
R41275 n3_11583_11048 n3_11583_11231 1.161905e-01
R41276 n3_11583_11231 n3_11583_11264 2.095238e-02
R41277 n3_11583_11264 n3_11583_11447 1.161905e-01
R41278 n3_11583_11447 n3_11583_11480 2.095238e-02
R41279 n3_11583_11480 n3_11583_11663 1.161905e-01
R41280 n3_11583_11663 n3_11583_11674 6.984127e-03
R41281 n3_11583_11674 n3_11583_11696 1.396825e-02
R41282 n3_11583_11696 n3_11583_11770 4.698413e-02
R41283 n3_11583_11770 n3_11583_11879 6.920635e-02
R41284 n3_11583_11879 n3_11583_11912 2.095238e-02
R41285 n3_11583_11912 n3_11583_12095 1.161905e-01
R41286 n3_11583_12095 n3_11583_12128 2.095238e-02
R41287 n3_11583_12128 n3_11583_12311 1.161905e-01
R41288 n3_11583_12311 n3_11583_12344 2.095238e-02
R41289 n3_11583_12344 n3_11583_12527 1.161905e-01
R41290 n3_11583_12527 n3_11583_12560 2.095238e-02
R41291 n3_11583_12560 n3_11583_12743 1.161905e-01
R41292 n3_11583_12959 n3_11583_12992 2.095238e-02
R41293 n3_11583_12992 n3_11583_13175 1.161905e-01
R41294 n3_11583_13175 n3_11583_13208 2.095238e-02
R41295 n3_11583_13208 n3_11583_13391 1.161905e-01
R41296 n3_11583_13391 n3_11583_13424 2.095238e-02
R41297 n3_11583_13424 n3_11583_13607 1.161905e-01
R41298 n3_11583_13607 n3_11583_13640 2.095238e-02
R41299 n3_11583_13640 n3_11583_13774 8.507937e-02
R41300 n3_11583_13774 n3_11583_13823 3.111111e-02
R41301 n3_11583_13823 n3_11583_13856 2.095238e-02
R41302 n3_11583_13856 n3_11583_13924 4.317460e-02
R41303 n3_11583_13924 n3_11583_14012 5.587302e-02
R41304 n3_11583_14012 n3_11583_14020 5.079365e-03
R41305 n3_11583_14020 n3_11583_14039 1.206349e-02
R41306 n3_11583_14039 n3_11583_14072 2.095238e-02
R41307 n3_11583_14072 n3_11583_14220 9.396825e-02
R41308 n3_11583_14220 n3_11583_14255 2.222222e-02
R41309 n3_11583_14255 n3_11583_14288 2.095238e-02
R41310 n3_11583_14288 n3_11583_14471 1.161905e-01
R41311 n3_11583_14471 n3_11583_14504 2.095238e-02
R41312 n3_11583_14504 n3_11583_14660 9.904762e-02
R41313 n3_11583_14660 n3_11583_14687 1.714286e-02
R41314 n3_11583_14687 n3_11583_14720 2.095238e-02
R41315 n3_11583_14720 n3_11583_14903 1.161905e-01
R41316 n3_11583_14903 n3_11583_14936 2.095238e-02
R41317 n3_11583_15335 n3_11583_15368 2.095238e-02
R41318 n3_11583_15368 n3_11583_15551 1.161905e-01
R41319 n3_11583_15551 n3_11583_15584 2.095238e-02
R41320 n3_11583_15584 n3_11583_15740 9.904762e-02
R41321 n3_11583_15740 n3_11583_15767 1.714286e-02
R41322 n3_11583_15767 n3_11583_15800 2.095238e-02
R41323 n3_11583_15800 n3_11583_15948 9.396825e-02
R41324 n3_11583_15948 n3_11583_15956 5.079365e-03
R41325 n3_11583_15956 n3_11583_15983 1.714286e-02
R41326 n3_11583_15983 n3_11583_16016 2.095238e-02
R41327 n3_11583_16016 n3_11583_16172 9.904762e-02
R41328 n3_11583_16172 n3_11583_16174 1.269841e-03
R41329 n3_11583_16174 n3_11583_16199 1.587302e-02
R41330 n3_11583_16199 n3_11583_16232 2.095238e-02
R41331 n3_11583_16232 n3_11583_16270 2.412698e-02
R41332 n3_11583_16270 n3_11583_16415 9.206349e-02
R41333 n3_11583_16415 n3_11583_16448 2.095238e-02
R41334 n3_11583_16448 n3_11583_16604 9.904762e-02
R41335 n3_11583_16604 n3_11583_16631 1.714286e-02
R41336 n3_11583_16631 n3_11583_16664 2.095238e-02
R41337 n3_11583_16664 n3_11583_16847 1.161905e-01
R41338 n3_11583_16847 n3_11583_16880 2.095238e-02
R41339 n3_11583_16880 n3_11583_17063 1.161905e-01
R41340 n3_11583_17063 n3_11583_17096 2.095238e-02
R41341 n3_11583_17096 n3_11583_17244 9.396825e-02
R41342 n3_11583_17468 n3_11583_17495 1.714286e-02
R41343 n3_11583_17495 n3_11583_17528 2.095238e-02
R41344 n3_11583_17528 n3_11583_17684 9.904762e-02
R41345 n3_11583_17684 n3_11583_17711 1.714286e-02
R41346 n3_11583_17711 n3_11583_17744 2.095238e-02
R41347 n3_11583_17744 n3_11583_17927 1.161905e-01
R41348 n3_11583_17927 n3_11583_17960 2.095238e-02
R41349 n3_11583_17960 n3_11583_18143 1.161905e-01
R41350 n3_11583_18143 n3_11583_18176 2.095238e-02
R41351 n3_11583_18176 n3_11583_18332 9.904762e-02
R41352 n3_11583_18332 n3_11583_18359 1.714286e-02
R41353 n3_11583_18359 n3_11583_18392 2.095238e-02
R41354 n3_11583_18392 n3_11583_18424 2.031746e-02
R41355 n3_11583_18424 n3_11583_18520 6.095238e-02
R41356 n3_11583_18520 n3_11583_18527 4.444444e-03
R41357 n3_11583_18527 n3_11583_18548 1.333333e-02
R41358 n3_11583_18548 n3_11583_18575 1.714286e-02
R41359 n3_11583_18575 n3_11583_18608 2.095238e-02
R41360 n3_11583_18608 n3_11583_18764 9.904762e-02
R41361 n3_11583_18764 n3_11583_18791 1.714286e-02
R41362 n3_11583_18791 n3_11583_18824 2.095238e-02
R41363 n3_11583_18824 n3_11583_19007 1.161905e-01
R41364 n3_11583_19007 n3_11583_19040 2.095238e-02
R41365 n3_11583_19040 n3_11583_19223 1.161905e-01
R41366 n3_11583_19223 n3_11583_19256 2.095238e-02
R41367 n3_11583_19256 n3_11583_19404 9.396825e-02
R41368 n3_11583_19404 n3_11583_19412 5.079365e-03
R41369 n3_11583_19412 n3_11583_19439 1.714286e-02
R41370 n3_11583_19439 n3_11583_19472 2.095238e-02
R41371 n3_11583_19871 n3_11583_19904 2.095238e-02
R41372 n3_11583_19904 n3_11583_20087 1.161905e-01
R41373 n3_11583_20087 n3_11583_20120 2.095238e-02
R41374 n3_11583_20120 n3_11583_20303 1.161905e-01
R41375 n3_11583_20303 n3_11583_20336 2.095238e-02
R41376 n3_11583_20336 n3_11583_20519 1.161905e-01
R41377 n3_11583_20519 n3_11583_20552 2.095238e-02
R41378 n3_11583_20552 n3_11583_20674 7.746032e-02
R41379 n3_11583_20674 n3_11583_20687 8.253968e-03
R41380 n3_11583_20687 n3_11583_20735 3.047619e-02
R41381 n3_11583_20735 n3_11583_20768 2.095238e-02
R41382 n3_11583_20768 n3_11583_20770 1.269841e-03
R41383 n3_11583_20770 n3_11583_20951 1.149206e-01
R41384 n3_11583_20951 n3_11583_20984 2.095238e-02
R41385 n3_11771_215 n3_11771_248 2.095238e-02
R41386 n3_11771_248 n3_11771_383 8.571429e-02
R41387 n3_11771_383 n3_11771_424 2.603175e-02
R41388 n3_11771_424 n3_11771_431 4.444444e-03
R41389 n3_11771_520 n3_11771_647 8.063492e-02
R41390 n3_11771_647 n3_11771_680 2.095238e-02
R41391 n3_11771_680 n3_11771_863 1.161905e-01
R41392 n3_11771_863 n3_11771_896 2.095238e-02
R41393 n3_11771_896 n3_11771_1079 1.161905e-01
R41394 n3_11771_1079 n3_11771_1112 2.095238e-02
R41395 n3_11771_1112 n3_11771_1295 1.161905e-01
R41396 n3_11771_1295 n3_11771_1328 2.095238e-02
R41397 n3_11771_1328 n3_11771_1511 1.161905e-01
R41398 n3_11771_1511 n3_11771_1544 2.095238e-02
R41399 n3_11771_1544 n3_11771_1727 1.161905e-01
R41400 n3_11771_1727 n3_11771_1760 2.095238e-02
R41401 n3_11771_1760 n3_11771_1894 8.507937e-02
R41402 n3_11771_1894 n3_11771_1943 3.111111e-02
R41403 n3_11771_1943 n3_11771_1976 2.095238e-02
R41404 n3_11771_1976 n3_11771_2159 1.161905e-01
R41405 n3_11771_2159 n3_11771_2192 2.095238e-02
R41406 n3_11771_2192 n3_11771_2375 1.161905e-01
R41407 n3_11771_2375 n3_11771_2408 2.095238e-02
R41408 n3_11771_2408 n3_11771_2542 8.507937e-02
R41409 n3_11771_2542 n3_11771_2543 6.349206e-04
R41410 n3_11771_2543 n3_11771_2591 3.047619e-02
R41411 n3_11771_2591 n3_11771_2624 2.095238e-02
R41412 n3_11771_2624 n3_11771_2674 3.174603e-02
R41413 n3_11771_2760 n3_11771_2770 6.349206e-03
R41414 n3_11771_2770 n3_11771_2807 2.349206e-02
R41415 n3_11771_2807 n3_11771_2840 2.095238e-02
R41416 n3_11771_2840 n3_11771_2974 8.507937e-02
R41417 n3_11771_2974 n3_11771_3023 3.111111e-02
R41418 n3_11771_3023 n3_11771_3056 2.095238e-02
R41419 n3_11771_3056 n3_11771_3239 1.161905e-01
R41420 n3_11771_3239 n3_11771_3272 2.095238e-02
R41421 n3_11771_3272 n3_11771_3455 1.161905e-01
R41422 n3_11771_3455 n3_11771_3488 2.095238e-02
R41423 n3_11771_3488 n3_11771_3622 8.507937e-02
R41424 n3_11771_3622 n3_11771_3671 3.111111e-02
R41425 n3_11771_3671 n3_11771_3704 2.095238e-02
R41426 n3_11771_3704 n3_11771_3887 1.161905e-01
R41427 n3_11771_3887 n3_11771_3920 2.095238e-02
R41428 n3_11771_3920 n3_11771_4103 1.161905e-01
R41429 n3_11771_4103 n3_11771_4136 2.095238e-02
R41430 n3_11771_4136 n3_11771_4270 8.507937e-02
R41431 n3_11771_4270 n3_11771_4319 3.111111e-02
R41432 n3_11771_4319 n3_11771_4352 2.095238e-02
R41433 n3_11771_4352 n3_11771_4535 1.161905e-01
R41434 n3_11771_4535 n3_11771_4568 2.095238e-02
R41435 n3_11771_4568 n3_11771_4702 8.507937e-02
R41436 n3_11771_4702 n3_11771_4751 3.111111e-02
R41437 n3_11771_4751 n3_11771_4784 2.095238e-02
R41438 n3_11771_4784 n3_11771_4924 8.888889e-02
R41439 n3_11771_5000 n3_11771_5020 1.269841e-02
R41440 n3_11771_5020 n3_11771_5183 1.034921e-01
R41441 n3_11771_5183 n3_11771_5216 2.095238e-02
R41442 n3_11771_5216 n3_11771_5350 8.507937e-02
R41443 n3_11771_5350 n3_11771_5399 3.111111e-02
R41444 n3_11771_5399 n3_11771_5432 2.095238e-02
R41445 n3_11771_5432 n3_11771_5566 8.507937e-02
R41446 n3_11771_5566 n3_11771_5615 3.111111e-02
R41447 n3_11771_5615 n3_11771_5648 2.095238e-02
R41448 n3_11771_5648 n3_11771_5782 8.507937e-02
R41449 n3_11771_5782 n3_11771_5831 3.111111e-02
R41450 n3_11771_5831 n3_11771_5864 2.095238e-02
R41451 n3_11771_5864 n3_11771_6047 1.161905e-01
R41452 n3_11771_6047 n3_11771_6080 2.095238e-02
R41453 n3_11771_6080 n3_11771_6263 1.161905e-01
R41454 n3_11771_6263 n3_11771_6296 2.095238e-02
R41455 n3_11771_6296 n3_11771_6430 8.507937e-02
R41456 n3_11771_6430 n3_11771_6479 3.111111e-02
R41457 n3_11771_6479 n3_11771_6512 2.095238e-02
R41458 n3_11771_6512 n3_11771_6646 8.507937e-02
R41459 n3_11771_6646 n3_11771_6695 3.111111e-02
R41460 n3_11771_6695 n3_11771_6728 2.095238e-02
R41461 n3_11771_6728 n3_11771_6862 8.507937e-02
R41462 n3_11771_6862 n3_11771_6911 3.111111e-02
R41463 n3_11771_6911 n3_11771_6944 2.095238e-02
R41464 n3_11771_6944 n3_11771_7078 8.507937e-02
R41465 n3_11771_7078 n3_11771_7127 3.111111e-02
R41466 n3_11771_7127 n3_11771_7160 2.095238e-02
R41467 n3_11771_7160 n3_11771_7174 8.888889e-03
R41468 n3_11771_7270 n3_11771_7294 1.523810e-02
R41469 n3_11771_7294 n3_11771_7343 3.111111e-02
R41470 n3_11771_7343 n3_11771_7376 2.095238e-02
R41471 n3_11771_7376 n3_11771_7510 8.507937e-02
R41472 n3_11771_7510 n3_11771_7559 3.111111e-02
R41473 n3_11771_7559 n3_11771_7592 2.095238e-02
R41474 n3_11771_7592 n3_11771_7775 1.161905e-01
R41475 n3_11771_7775 n3_11771_7808 2.095238e-02
R41476 n3_11771_7808 n3_11771_7991 1.161905e-01
R41477 n3_11771_7991 n3_11771_8024 2.095238e-02
R41478 n3_11771_8024 n3_11771_8207 1.161905e-01
R41479 n3_11771_8207 n3_11771_8240 2.095238e-02
R41480 n3_11771_8240 n3_11771_8423 1.161905e-01
R41481 n3_11771_8423 n3_11771_8456 2.095238e-02
R41482 n3_11771_8456 n3_11771_8639 1.161905e-01
R41483 n3_11771_8639 n3_11771_8672 2.095238e-02
R41484 n3_11771_8672 n3_11771_8855 1.161905e-01
R41485 n3_11771_8855 n3_11771_8888 2.095238e-02
R41486 n3_11771_8888 n3_11771_9071 1.161905e-01
R41487 n3_11771_9071 n3_11771_9104 2.095238e-02
R41488 n3_11771_9104 n3_11771_9287 1.161905e-01
R41489 n3_11771_9287 n3_11771_9320 2.095238e-02
R41490 n3_11771_9320 n3_11771_9424 6.603175e-02
R41491 n3_11771_9503 n3_11771_9520 1.079365e-02
R41492 n3_11771_9520 n3_11771_9536 1.015873e-02
R41493 n3_11771_9536 n3_11771_9719 1.161905e-01
R41494 n3_11771_9719 n3_11771_9752 2.095238e-02
R41495 n3_11771_9752 n3_11771_9935 1.161905e-01
R41496 n3_11771_9935 n3_11771_9968 2.095238e-02
R41497 n3_11771_9968 n3_11771_10151 1.161905e-01
R41498 n3_11771_10151 n3_11771_10184 2.095238e-02
R41499 n3_11771_10184 n3_11771_10367 1.161905e-01
R41500 n3_11771_10367 n3_11771_10400 2.095238e-02
R41501 n3_11771_10616 n3_11771_10799 1.161905e-01
R41502 n3_11771_10799 n3_11771_10832 2.095238e-02
R41503 n3_11771_10832 n3_11771_11015 1.161905e-01
R41504 n3_11771_11015 n3_11771_11048 2.095238e-02
R41505 n3_11771_11048 n3_11771_11231 1.161905e-01
R41506 n3_11771_11231 n3_11771_11264 2.095238e-02
R41507 n3_11771_11264 n3_11771_11447 1.161905e-01
R41508 n3_11771_11447 n3_11771_11480 2.095238e-02
R41509 n3_11771_11480 n3_11771_11663 1.161905e-01
R41510 n3_11771_11663 n3_11771_11674 6.984127e-03
R41511 n3_11771_11674 n3_11771_11696 1.396825e-02
R41512 n3_11771_11770 n3_11771_11879 6.920635e-02
R41513 n3_11771_11879 n3_11771_11912 2.095238e-02
R41514 n3_11771_11912 n3_11771_12095 1.161905e-01
R41515 n3_11771_12095 n3_11771_12128 2.095238e-02
R41516 n3_11771_12128 n3_11771_12311 1.161905e-01
R41517 n3_11771_12311 n3_11771_12344 2.095238e-02
R41518 n3_11771_12344 n3_11771_12527 1.161905e-01
R41519 n3_11771_12527 n3_11771_12560 2.095238e-02
R41520 n3_11771_12560 n3_11771_12743 1.161905e-01
R41521 n3_11771_12743 n3_11771_12776 2.095238e-02
R41522 n3_11771_12776 n3_11771_12959 1.161905e-01
R41523 n3_11771_12959 n3_11771_12992 2.095238e-02
R41524 n3_11771_12992 n3_11771_13175 1.161905e-01
R41525 n3_11771_13175 n3_11771_13208 2.095238e-02
R41526 n3_11771_13208 n3_11771_13391 1.161905e-01
R41527 n3_11771_13391 n3_11771_13424 2.095238e-02
R41528 n3_11771_13424 n3_11771_13607 1.161905e-01
R41529 n3_11771_13607 n3_11771_13640 2.095238e-02
R41530 n3_11771_13640 n3_11771_13774 8.507937e-02
R41531 n3_11771_13774 n3_11771_13823 3.111111e-02
R41532 n3_11771_13823 n3_11771_13856 2.095238e-02
R41533 n3_11771_13856 n3_11771_13924 4.317460e-02
R41534 n3_11771_14012 n3_11771_14020 5.079365e-03
R41535 n3_11771_14020 n3_11771_14039 1.206349e-02
R41536 n3_11771_14039 n3_11771_14072 2.095238e-02
R41537 n3_11771_14072 n3_11771_14220 9.396825e-02
R41538 n3_11771_14220 n3_11771_14255 2.222222e-02
R41539 n3_11771_14255 n3_11771_14288 2.095238e-02
R41540 n3_11771_14288 n3_11771_14471 1.161905e-01
R41541 n3_11771_14471 n3_11771_14504 2.095238e-02
R41542 n3_11771_14504 n3_11771_14660 9.904762e-02
R41543 n3_11771_14660 n3_11771_14687 1.714286e-02
R41544 n3_11771_14687 n3_11771_14720 2.095238e-02
R41545 n3_11771_14720 n3_11771_14903 1.161905e-01
R41546 n3_11771_14903 n3_11771_14936 2.095238e-02
R41547 n3_11771_14936 n3_11771_15119 1.161905e-01
R41548 n3_11771_15119 n3_11771_15152 2.095238e-02
R41549 n3_11771_15152 n3_11771_15335 1.161905e-01
R41550 n3_11771_15335 n3_11771_15368 2.095238e-02
R41551 n3_11771_15368 n3_11771_15551 1.161905e-01
R41552 n3_11771_15551 n3_11771_15584 2.095238e-02
R41553 n3_11771_15584 n3_11771_15740 9.904762e-02
R41554 n3_11771_15740 n3_11771_15767 1.714286e-02
R41555 n3_11771_15767 n3_11771_15800 2.095238e-02
R41556 n3_11771_15800 n3_11771_15948 9.396825e-02
R41557 n3_11771_15948 n3_11771_15956 5.079365e-03
R41558 n3_11771_15956 n3_11771_15983 1.714286e-02
R41559 n3_11771_15983 n3_11771_16016 2.095238e-02
R41560 n3_11771_16016 n3_11771_16172 9.904762e-02
R41561 n3_11771_16172 n3_11771_16174 1.269841e-03
R41562 n3_11771_16174 n3_11771_16199 1.587302e-02
R41563 n3_11771_16270 n3_11771_16415 9.206349e-02
R41564 n3_11771_16415 n3_11771_16448 2.095238e-02
R41565 n3_11771_16448 n3_11771_16604 9.904762e-02
R41566 n3_11771_16604 n3_11771_16631 1.714286e-02
R41567 n3_11771_16631 n3_11771_16664 2.095238e-02
R41568 n3_11771_16664 n3_11771_16847 1.161905e-01
R41569 n3_11771_16847 n3_11771_16880 2.095238e-02
R41570 n3_11771_16880 n3_11771_17063 1.161905e-01
R41571 n3_11771_17063 n3_11771_17096 2.095238e-02
R41572 n3_11771_17096 n3_11771_17244 9.396825e-02
R41573 n3_11771_17244 n3_11771_17279 2.222222e-02
R41574 n3_11771_17279 n3_11771_17312 2.095238e-02
R41575 n3_11771_17312 n3_11771_17468 9.904762e-02
R41576 n3_11771_17468 n3_11771_17495 1.714286e-02
R41577 n3_11771_17495 n3_11771_17528 2.095238e-02
R41578 n3_11771_17528 n3_11771_17684 9.904762e-02
R41579 n3_11771_17684 n3_11771_17711 1.714286e-02
R41580 n3_11771_17711 n3_11771_17744 2.095238e-02
R41581 n3_11771_17744 n3_11771_17927 1.161905e-01
R41582 n3_11771_17927 n3_11771_17960 2.095238e-02
R41583 n3_11771_17960 n3_11771_18143 1.161905e-01
R41584 n3_11771_18143 n3_11771_18176 2.095238e-02
R41585 n3_11771_18176 n3_11771_18332 9.904762e-02
R41586 n3_11771_18332 n3_11771_18359 1.714286e-02
R41587 n3_11771_18359 n3_11771_18392 2.095238e-02
R41588 n3_11771_18392 n3_11771_18424 2.031746e-02
R41589 n3_11771_18520 n3_11771_18527 4.444444e-03
R41590 n3_11771_18527 n3_11771_18548 1.333333e-02
R41591 n3_11771_18548 n3_11771_18575 1.714286e-02
R41592 n3_11771_18575 n3_11771_18608 2.095238e-02
R41593 n3_11771_18608 n3_11771_18764 9.904762e-02
R41594 n3_11771_18764 n3_11771_18791 1.714286e-02
R41595 n3_11771_18791 n3_11771_18824 2.095238e-02
R41596 n3_11771_18824 n3_11771_19007 1.161905e-01
R41597 n3_11771_19007 n3_11771_19040 2.095238e-02
R41598 n3_11771_19040 n3_11771_19223 1.161905e-01
R41599 n3_11771_19223 n3_11771_19256 2.095238e-02
R41600 n3_11771_19256 n3_11771_19404 9.396825e-02
R41601 n3_11771_19404 n3_11771_19412 5.079365e-03
R41602 n3_11771_19412 n3_11771_19439 1.714286e-02
R41603 n3_11771_19439 n3_11771_19472 2.095238e-02
R41604 n3_11771_19472 n3_11771_19655 1.161905e-01
R41605 n3_11771_19655 n3_11771_19688 2.095238e-02
R41606 n3_11771_19688 n3_11771_19871 1.161905e-01
R41607 n3_11771_19871 n3_11771_19904 2.095238e-02
R41608 n3_11771_19904 n3_11771_20087 1.161905e-01
R41609 n3_11771_20087 n3_11771_20120 2.095238e-02
R41610 n3_11771_20120 n3_11771_20303 1.161905e-01
R41611 n3_11771_20303 n3_11771_20336 2.095238e-02
R41612 n3_11771_20336 n3_11771_20519 1.161905e-01
R41613 n3_11771_20519 n3_11771_20552 2.095238e-02
R41614 n3_11771_20552 n3_11771_20674 7.746032e-02
R41615 n3_11771_20674 n3_11771_20687 8.253968e-03
R41616 n3_11771_20768 n3_11771_20770 1.269841e-03
R41617 n3_11771_20770 n3_11771_20951 1.149206e-01
R41618 n3_11771_20951 n3_11771_20984 2.095238e-02
R41619 n3_11864_215 n3_11864_248 2.095238e-02
R41620 n3_11864_248 n3_11864_383 8.571429e-02
R41621 n3_11864_383 n3_11864_431 3.047619e-02
R41622 n3_11864_431 n3_11864_464 2.095238e-02
R41623 n3_11864_464 n3_11864_647 1.161905e-01
R41624 n3_11864_647 n3_11864_680 2.095238e-02
R41625 n3_11864_680 n3_11864_863 1.161905e-01
R41626 n3_11864_863 n3_11864_896 2.095238e-02
R41627 n3_11864_896 n3_11864_1079 1.161905e-01
R41628 n3_11864_1079 n3_11864_1112 2.095238e-02
R41629 n3_11864_1112 n3_11864_1295 1.161905e-01
R41630 n3_11864_1295 n3_11864_1328 2.095238e-02
R41631 n3_11864_1328 n3_11864_1511 1.161905e-01
R41632 n3_11864_1511 n3_11864_1544 2.095238e-02
R41633 n3_11864_1544 n3_11864_1727 1.161905e-01
R41634 n3_11864_1727 n3_11864_1760 2.095238e-02
R41635 n3_11864_1760 n3_11864_1894 8.507937e-02
R41636 n3_11864_1894 n3_11864_1943 3.111111e-02
R41637 n3_11864_1943 n3_11864_1976 2.095238e-02
R41638 n3_11864_1976 n3_11864_2159 1.161905e-01
R41639 n3_11864_2159 n3_11864_2192 2.095238e-02
R41640 n3_11864_2192 n3_11864_2375 1.161905e-01
R41641 n3_11864_2375 n3_11864_2408 2.095238e-02
R41642 n3_11864_2408 n3_11864_2542 8.507937e-02
R41643 n3_11864_2542 n3_11864_2543 6.349206e-04
R41644 n3_11864_2543 n3_11864_2591 3.047619e-02
R41645 n3_11864_2591 n3_11864_2624 2.095238e-02
R41646 n3_11864_18527 n3_11864_18575 3.047619e-02
R41647 n3_11864_18575 n3_11864_18608 2.095238e-02
R41648 n3_11864_18608 n3_11864_18764 9.904762e-02
R41649 n3_11864_18764 n3_11864_18791 1.714286e-02
R41650 n3_11864_18791 n3_11864_18824 2.095238e-02
R41651 n3_11864_18824 n3_11864_19007 1.161905e-01
R41652 n3_11864_19007 n3_11864_19040 2.095238e-02
R41653 n3_11864_19040 n3_11864_19223 1.161905e-01
R41654 n3_11864_19223 n3_11864_19256 2.095238e-02
R41655 n3_11864_19256 n3_11864_19404 9.396825e-02
R41656 n3_11864_19404 n3_11864_19439 2.222222e-02
R41657 n3_11864_19439 n3_11864_19472 2.095238e-02
R41658 n3_11864_19472 n3_11864_19655 1.161905e-01
R41659 n3_11864_19655 n3_11864_19688 2.095238e-02
R41660 n3_11864_19688 n3_11864_19871 1.161905e-01
R41661 n3_11864_19871 n3_11864_19904 2.095238e-02
R41662 n3_11864_19904 n3_11864_20087 1.161905e-01
R41663 n3_11864_20087 n3_11864_20120 2.095238e-02
R41664 n3_11864_20120 n3_11864_20303 1.161905e-01
R41665 n3_11864_20303 n3_11864_20336 2.095238e-02
R41666 n3_11864_20336 n3_11864_20519 1.161905e-01
R41667 n3_11864_20519 n3_11864_20552 2.095238e-02
R41668 n3_11864_20552 n3_11864_20687 8.571429e-02
R41669 n3_11864_20687 n3_11864_20735 3.047619e-02
R41670 n3_11864_20735 n3_11864_20768 2.095238e-02
R41671 n3_11864_20768 n3_11864_20951 1.161905e-01
R41672 n3_11864_20951 n3_11864_20984 2.095238e-02
R41673 n3_13650_215 n3_13650_248 2.095238e-02
R41674 n3_13650_248 n3_13650_383 8.571429e-02
R41675 n3_13650_383 n3_13650_431 3.047619e-02
R41676 n3_13650_431 n3_13650_464 2.095238e-02
R41677 n3_13650_464 n3_13650_647 1.161905e-01
R41678 n3_13650_647 n3_13650_680 2.095238e-02
R41679 n3_13650_680 n3_13650_863 1.161905e-01
R41680 n3_13650_863 n3_13650_896 2.095238e-02
R41681 n3_13650_896 n3_13650_1079 1.161905e-01
R41682 n3_13650_1079 n3_13650_1112 2.095238e-02
R41683 n3_13650_1112 n3_13650_1295 1.161905e-01
R41684 n3_13650_1295 n3_13650_1328 2.095238e-02
R41685 n3_13650_1328 n3_13650_1511 1.161905e-01
R41686 n3_13650_1511 n3_13650_1544 2.095238e-02
R41687 n3_13650_1544 n3_13650_1727 1.161905e-01
R41688 n3_13650_1727 n3_13650_1760 2.095238e-02
R41689 n3_13650_1760 n3_13650_1894 8.507937e-02
R41690 n3_13650_1894 n3_13650_1943 3.111111e-02
R41691 n3_13650_1943 n3_13650_1976 2.095238e-02
R41692 n3_13650_1976 n3_13650_2159 1.161905e-01
R41693 n3_13650_2159 n3_13650_2192 2.095238e-02
R41694 n3_13650_2192 n3_13650_2375 1.161905e-01
R41695 n3_13650_2375 n3_13650_2408 2.095238e-02
R41696 n3_13650_2408 n3_13650_2445 2.349206e-02
R41697 n3_13650_2445 n3_13650_2542 6.158730e-02
R41698 n3_13650_2542 n3_13650_2543 6.349206e-04
R41699 n3_13650_2543 n3_13650_2591 3.047619e-02
R41700 n3_13650_2591 n3_13650_2624 2.095238e-02
R41701 n3_13650_18527 n3_13650_18575 3.047619e-02
R41702 n3_13650_18575 n3_13650_18608 2.095238e-02
R41703 n3_13650_18608 n3_13650_18764 9.904762e-02
R41704 n3_13650_18764 n3_13650_18791 1.714286e-02
R41705 n3_13650_18791 n3_13650_18824 2.095238e-02
R41706 n3_13650_18824 n3_13650_19007 1.161905e-01
R41707 n3_13650_19007 n3_13650_19040 2.095238e-02
R41708 n3_13650_19040 n3_13650_19223 1.161905e-01
R41709 n3_13650_19223 n3_13650_19256 2.095238e-02
R41710 n3_13650_19256 n3_13650_19412 9.904762e-02
R41711 n3_13650_19412 n3_13650_19439 1.714286e-02
R41712 n3_13650_19439 n3_13650_19472 2.095238e-02
R41713 n3_13650_19472 n3_13650_19655 1.161905e-01
R41714 n3_13650_19655 n3_13650_19688 2.095238e-02
R41715 n3_13650_19688 n3_13650_19871 1.161905e-01
R41716 n3_13650_19871 n3_13650_19904 2.095238e-02
R41717 n3_13650_19904 n3_13650_20087 1.161905e-01
R41718 n3_13650_20087 n3_13650_20120 2.095238e-02
R41719 n3_13650_20120 n3_13650_20303 1.161905e-01
R41720 n3_13650_20303 n3_13650_20336 2.095238e-02
R41721 n3_13650_20336 n3_13650_20519 1.161905e-01
R41722 n3_13650_20519 n3_13650_20552 2.095238e-02
R41723 n3_13650_20552 n3_13650_20687 8.571429e-02
R41724 n3_13650_20687 n3_13650_20735 3.047619e-02
R41725 n3_13650_20735 n3_13650_20768 2.095238e-02
R41726 n3_13650_20768 n3_13650_20951 1.161905e-01
R41727 n3_13650_20951 n3_13650_20984 2.095238e-02
R41728 n3_13833_424 n3_13880_424 2.984127e-02
R41729 n3_13880_424 n3_14021_424 8.952381e-02
R41730 n3_13833_520 n3_13880_520 2.984127e-02
R41731 n3_13880_520 n3_14021_520 8.952381e-02
R41732 n3_13833_2674 n3_13880_2674 2.984127e-02
R41733 n3_13880_2674 n3_14021_2674 8.952381e-02
R41734 n3_13833_2770 n3_13880_2770 2.984127e-02
R41735 n3_13880_2770 n3_14021_2770 8.952381e-02
R41736 n3_13833_4924 n3_13880_4924 2.984127e-02
R41737 n3_13880_4924 n3_14021_4924 8.952381e-02
R41738 n3_13833_5020 n3_13880_5020 2.984127e-02
R41739 n3_13880_5020 n3_14021_5020 8.952381e-02
R41740 n3_13833_7174 n3_13880_7174 2.984127e-02
R41741 n3_13880_7174 n3_14021_7174 8.952381e-02
R41742 n3_13833_7270 n3_13880_7270 2.984127e-02
R41743 n3_13880_7270 n3_14021_7270 8.952381e-02
R41744 n3_13833_9424 n3_13880_9424 2.984127e-02
R41745 n3_13880_9424 n3_14021_9424 8.952381e-02
R41746 n3_13833_9520 n3_13880_9520 2.984127e-02
R41747 n3_13880_9520 n3_14021_9520 8.952381e-02
R41748 n3_13833_11674 n3_13880_11674 2.984127e-02
R41749 n3_13880_11674 n3_14021_11674 8.952381e-02
R41750 n3_13833_11770 n3_13880_11770 2.984127e-02
R41751 n3_13880_11770 n3_14021_11770 8.952381e-02
R41752 n3_13833_13924 n3_13880_13924 2.984127e-02
R41753 n3_13880_13924 n3_14021_13924 8.952381e-02
R41754 n3_13833_14020 n3_13880_14020 2.984127e-02
R41755 n3_13880_14020 n3_14021_14020 8.952381e-02
R41756 n3_13833_16174 n3_13880_16174 2.984127e-02
R41757 n3_13880_16174 n3_14021_16174 8.952381e-02
R41758 n3_13833_16270 n3_13880_16270 2.984127e-02
R41759 n3_13880_16270 n3_14021_16270 8.952381e-02
R41760 n3_13833_18424 n3_13880_18424 2.984127e-02
R41761 n3_13880_18424 n3_14021_18424 8.952381e-02
R41762 n3_13833_18520 n3_13880_18520 2.984127e-02
R41763 n3_13880_18520 n3_14021_18520 8.952381e-02
R41764 n3_13833_20674 n3_13880_20674 2.984127e-02
R41765 n3_13880_20674 n3_14021_20674 8.952381e-02
R41766 n3_13833_20770 n3_13880_20770 2.984127e-02
R41767 n3_13880_20770 n3_14021_20770 8.952381e-02
R41768 n3_13833_215 n3_13833_248 2.095238e-02
R41769 n3_13833_248 n3_13833_383 8.571429e-02
R41770 n3_13833_383 n3_13833_424 2.603175e-02
R41771 n3_13833_424 n3_13833_431 4.444444e-03
R41772 n3_13833_431 n3_13833_464 2.095238e-02
R41773 n3_13833_464 n3_13833_520 3.555556e-02
R41774 n3_13833_520 n3_13833_647 8.063492e-02
R41775 n3_13833_647 n3_13833_680 2.095238e-02
R41776 n3_13833_680 n3_13833_863 1.161905e-01
R41777 n3_13833_863 n3_13833_896 2.095238e-02
R41778 n3_13833_896 n3_13833_1079 1.161905e-01
R41779 n3_13833_1079 n3_13833_1112 2.095238e-02
R41780 n3_13833_1112 n3_13833_1295 1.161905e-01
R41781 n3_13833_1295 n3_13833_1328 2.095238e-02
R41782 n3_13833_1727 n3_13833_1760 2.095238e-02
R41783 n3_13833_1760 n3_13833_1894 8.507937e-02
R41784 n3_13833_1894 n3_13833_1943 3.111111e-02
R41785 n3_13833_1943 n3_13833_1976 2.095238e-02
R41786 n3_13833_1976 n3_13833_2159 1.161905e-01
R41787 n3_13833_2159 n3_13833_2192 2.095238e-02
R41788 n3_13833_2192 n3_13833_2375 1.161905e-01
R41789 n3_13833_2375 n3_13833_2408 2.095238e-02
R41790 n3_13833_2408 n3_13833_2445 2.349206e-02
R41791 n3_13833_2445 n3_13833_2542 6.158730e-02
R41792 n3_13833_2542 n3_13833_2543 6.349206e-04
R41793 n3_13833_2543 n3_13833_2591 3.047619e-02
R41794 n3_13833_2591 n3_13833_2624 2.095238e-02
R41795 n3_13833_2624 n3_13833_2674 3.174603e-02
R41796 n3_13833_2674 n3_13833_2770 6.095238e-02
R41797 n3_13833_2770 n3_13833_2807 2.349206e-02
R41798 n3_13833_2807 n3_13833_2840 2.095238e-02
R41799 n3_13833_2840 n3_13833_2877 2.349206e-02
R41800 n3_13833_2877 n3_13833_2974 6.158730e-02
R41801 n3_13833_2974 n3_13833_3023 3.111111e-02
R41802 n3_13833_3023 n3_13833_3056 2.095238e-02
R41803 n3_13833_3056 n3_13833_3239 1.161905e-01
R41804 n3_13833_3239 n3_13833_3272 2.095238e-02
R41805 n3_13833_3272 n3_13833_3455 1.161905e-01
R41806 n3_13833_3455 n3_13833_3488 2.095238e-02
R41807 n3_13833_3488 n3_13833_3622 8.507937e-02
R41808 n3_13833_3622 n3_13833_3671 3.111111e-02
R41809 n3_13833_3671 n3_13833_3704 2.095238e-02
R41810 n3_13833_4054 n3_13833_4103 3.111111e-02
R41811 n3_13833_4103 n3_13833_4136 2.095238e-02
R41812 n3_13833_4136 n3_13833_4270 8.507937e-02
R41813 n3_13833_4270 n3_13833_4319 3.111111e-02
R41814 n3_13833_4319 n3_13833_4352 2.095238e-02
R41815 n3_13833_4352 n3_13833_4535 1.161905e-01
R41816 n3_13833_4535 n3_13833_4568 2.095238e-02
R41817 n3_13833_4568 n3_13833_4702 8.507937e-02
R41818 n3_13833_4702 n3_13833_4751 3.111111e-02
R41819 n3_13833_4751 n3_13833_4784 2.095238e-02
R41820 n3_13833_4784 n3_13833_4924 8.888889e-02
R41821 n3_13833_4924 n3_13833_4967 2.730159e-02
R41822 n3_13833_4967 n3_13833_5000 2.095238e-02
R41823 n3_13833_5000 n3_13833_5020 1.269841e-02
R41824 n3_13833_5020 n3_13833_5134 7.238095e-02
R41825 n3_13833_5134 n3_13833_5183 3.111111e-02
R41826 n3_13833_5183 n3_13833_5216 2.095238e-02
R41827 n3_13833_5216 n3_13833_5350 8.507937e-02
R41828 n3_13833_5350 n3_13833_5399 3.111111e-02
R41829 n3_13833_5399 n3_13833_5432 2.095238e-02
R41830 n3_13833_5432 n3_13833_5615 1.161905e-01
R41831 n3_13833_5615 n3_13833_5648 2.095238e-02
R41832 n3_13833_5648 n3_13833_5782 8.507937e-02
R41833 n3_13833_5782 n3_13833_5831 3.111111e-02
R41834 n3_13833_5831 n3_13833_5864 2.095238e-02
R41835 n3_13833_6263 n3_13833_6296 2.095238e-02
R41836 n3_13833_6296 n3_13833_6430 8.507937e-02
R41837 n3_13833_6430 n3_13833_6479 3.111111e-02
R41838 n3_13833_6479 n3_13833_6512 2.095238e-02
R41839 n3_13833_6512 n3_13833_6646 8.507937e-02
R41840 n3_13833_6646 n3_13833_6695 3.111111e-02
R41841 n3_13833_6695 n3_13833_6728 2.095238e-02
R41842 n3_13833_6728 n3_13833_6911 1.161905e-01
R41843 n3_13833_6911 n3_13833_6944 2.095238e-02
R41844 n3_13833_6944 n3_13833_7127 1.161905e-01
R41845 n3_13833_7127 n3_13833_7160 2.095238e-02
R41846 n3_13833_7160 n3_13833_7174 8.888889e-03
R41847 n3_13833_7174 n3_13833_7270 6.095238e-02
R41848 n3_13833_7270 n3_13833_7343 4.634921e-02
R41849 n3_13833_7343 n3_13833_7376 2.095238e-02
R41850 n3_13833_7376 n3_13833_7559 1.161905e-01
R41851 n3_13833_7559 n3_13833_7592 2.095238e-02
R41852 n3_13833_7592 n3_13833_7775 1.161905e-01
R41853 n3_13833_7775 n3_13833_7808 2.095238e-02
R41854 n3_13833_7808 n3_13833_7845 2.349206e-02
R41855 n3_13833_7845 n3_13833_7942 6.158730e-02
R41856 n3_13833_7942 n3_13833_7991 3.111111e-02
R41857 n3_13833_7991 n3_13833_8024 2.095238e-02
R41858 n3_13833_8024 n3_13833_8207 1.161905e-01
R41859 n3_13833_8207 n3_13833_8240 2.095238e-02
R41860 n3_13833_8456 n3_13833_8639 1.161905e-01
R41861 n3_13833_8639 n3_13833_8672 2.095238e-02
R41862 n3_13833_8672 n3_13833_8806 8.507937e-02
R41863 n3_13833_8806 n3_13833_8855 3.111111e-02
R41864 n3_13833_8855 n3_13833_8888 2.095238e-02
R41865 n3_13833_8888 n3_13833_8925 2.349206e-02
R41866 n3_13833_8925 n3_13833_9022 6.158730e-02
R41867 n3_13833_9022 n3_13833_9071 3.111111e-02
R41868 n3_13833_9071 n3_13833_9104 2.095238e-02
R41869 n3_13833_9104 n3_13833_9287 1.161905e-01
R41870 n3_13833_9287 n3_13833_9320 2.095238e-02
R41871 n3_13833_9320 n3_13833_9424 6.603175e-02
R41872 n3_13833_9424 n3_13833_9503 5.015873e-02
R41873 n3_13833_9503 n3_13833_9520 1.079365e-02
R41874 n3_13833_9520 n3_13833_9536 1.015873e-02
R41875 n3_13833_9536 n3_13833_9719 1.161905e-01
R41876 n3_13833_9719 n3_13833_9752 2.095238e-02
R41877 n3_13833_9752 n3_13833_9886 8.507937e-02
R41878 n3_13833_9886 n3_13833_9935 3.111111e-02
R41879 n3_13833_9935 n3_13833_9968 2.095238e-02
R41880 n3_13833_9968 n3_13833_10005 2.349206e-02
R41881 n3_13833_10005 n3_13833_10102 6.158730e-02
R41882 n3_13833_10102 n3_13833_10151 3.111111e-02
R41883 n3_13833_10151 n3_13833_10184 2.095238e-02
R41884 n3_13833_10184 n3_13833_10367 1.161905e-01
R41885 n3_13833_10367 n3_13833_10400 2.095238e-02
R41886 n3_13833_10799 n3_13833_10832 2.095238e-02
R41887 n3_13833_10832 n3_13833_10988 9.904762e-02
R41888 n3_13833_10988 n3_13833_11015 1.714286e-02
R41889 n3_13833_11015 n3_13833_11048 2.095238e-02
R41890 n3_13833_11048 n3_13833_11204 9.904762e-02
R41891 n3_13833_11204 n3_13833_11231 1.714286e-02
R41892 n3_13833_11231 n3_13833_11264 2.095238e-02
R41893 n3_13833_11264 n3_13833_11447 1.161905e-01
R41894 n3_13833_11447 n3_13833_11480 2.095238e-02
R41895 n3_13833_11480 n3_13833_11663 1.161905e-01
R41896 n3_13833_11663 n3_13833_11674 6.984127e-03
R41897 n3_13833_11674 n3_13833_11696 1.396825e-02
R41898 n3_13833_11696 n3_13833_11770 4.698413e-02
R41899 n3_13833_11770 n3_13833_11879 6.920635e-02
R41900 n3_13833_11879 n3_13833_11912 2.095238e-02
R41901 n3_13833_11912 n3_13833_12068 9.904762e-02
R41902 n3_13833_12068 n3_13833_12095 1.714286e-02
R41903 n3_13833_12095 n3_13833_12128 2.095238e-02
R41904 n3_13833_12128 n3_13833_12284 9.904762e-02
R41905 n3_13833_12284 n3_13833_12311 1.714286e-02
R41906 n3_13833_12311 n3_13833_12344 2.095238e-02
R41907 n3_13833_12344 n3_13833_12527 1.161905e-01
R41908 n3_13833_12527 n3_13833_12560 2.095238e-02
R41909 n3_13833_12560 n3_13833_12743 1.161905e-01
R41910 n3_13833_12959 n3_13833_12992 2.095238e-02
R41911 n3_13833_12992 n3_13833_13175 1.161905e-01
R41912 n3_13833_13175 n3_13833_13208 2.095238e-02
R41913 n3_13833_13208 n3_13833_13391 1.161905e-01
R41914 n3_13833_13391 n3_13833_13424 2.095238e-02
R41915 n3_13833_13424 n3_13833_13607 1.161905e-01
R41916 n3_13833_13607 n3_13833_13640 2.095238e-02
R41917 n3_13833_13640 n3_13833_13823 1.161905e-01
R41918 n3_13833_13823 n3_13833_13856 2.095238e-02
R41919 n3_13833_13856 n3_13833_13924 4.317460e-02
R41920 n3_13833_13924 n3_13833_14020 6.095238e-02
R41921 n3_13833_14020 n3_13833_14039 1.206349e-02
R41922 n3_13833_14039 n3_13833_14072 2.095238e-02
R41923 n3_13833_14072 n3_13833_14220 9.396825e-02
R41924 n3_13833_14220 n3_13833_14255 2.222222e-02
R41925 n3_13833_14255 n3_13833_14288 2.095238e-02
R41926 n3_13833_14288 n3_13833_14471 1.161905e-01
R41927 n3_13833_14471 n3_13833_14504 2.095238e-02
R41928 n3_13833_14504 n3_13833_14652 9.396825e-02
R41929 n3_13833_14652 n3_13833_14687 2.222222e-02
R41930 n3_13833_14687 n3_13833_14720 2.095238e-02
R41931 n3_13833_14720 n3_13833_14868 9.396825e-02
R41932 n3_13833_14868 n3_13833_14903 2.222222e-02
R41933 n3_13833_14903 n3_13833_14936 2.095238e-02
R41934 n3_13833_15335 n3_13833_15368 2.095238e-02
R41935 n3_13833_15368 n3_13833_15524 9.904762e-02
R41936 n3_13833_15524 n3_13833_15551 1.714286e-02
R41937 n3_13833_15551 n3_13833_15584 2.095238e-02
R41938 n3_13833_15584 n3_13833_15767 1.161905e-01
R41939 n3_13833_15767 n3_13833_15800 2.095238e-02
R41940 n3_13833_15800 n3_13833_15956 9.904762e-02
R41941 n3_13833_15956 n3_13833_15983 1.714286e-02
R41942 n3_13833_15983 n3_13833_16016 2.095238e-02
R41943 n3_13833_16016 n3_13833_16174 1.003175e-01
R41944 n3_13833_16174 n3_13833_16199 1.587302e-02
R41945 n3_13833_16199 n3_13833_16232 2.095238e-02
R41946 n3_13833_16232 n3_13833_16270 2.412698e-02
R41947 n3_13833_16270 n3_13833_16415 9.206349e-02
R41948 n3_13833_16415 n3_13833_16448 2.095238e-02
R41949 n3_13833_16448 n3_13833_16604 9.904762e-02
R41950 n3_13833_16604 n3_13833_16631 1.714286e-02
R41951 n3_13833_16631 n3_13833_16664 2.095238e-02
R41952 n3_13833_16664 n3_13833_16847 1.161905e-01
R41953 n3_13833_16847 n3_13833_16880 2.095238e-02
R41954 n3_13833_16880 n3_13833_17063 1.161905e-01
R41955 n3_13833_17063 n3_13833_17096 2.095238e-02
R41956 n3_13833_17495 n3_13833_17528 2.095238e-02
R41957 n3_13833_17528 n3_13833_17684 9.904762e-02
R41958 n3_13833_17684 n3_13833_17711 1.714286e-02
R41959 n3_13833_17711 n3_13833_17744 2.095238e-02
R41960 n3_13833_17744 n3_13833_17927 1.161905e-01
R41961 n3_13833_17927 n3_13833_17960 2.095238e-02
R41962 n3_13833_17960 n3_13833_18094 8.507937e-02
R41963 n3_13833_18094 n3_13833_18143 3.111111e-02
R41964 n3_13833_18143 n3_13833_18176 2.095238e-02
R41965 n3_13833_18176 n3_13833_18324 9.396825e-02
R41966 n3_13833_18324 n3_13833_18332 5.079365e-03
R41967 n3_13833_18332 n3_13833_18359 1.714286e-02
R41968 n3_13833_18359 n3_13833_18392 2.095238e-02
R41969 n3_13833_18392 n3_13833_18424 2.031746e-02
R41970 n3_13833_18424 n3_13833_18520 6.095238e-02
R41971 n3_13833_18520 n3_13833_18527 4.444444e-03
R41972 n3_13833_18527 n3_13833_18575 3.047619e-02
R41973 n3_13833_18575 n3_13833_18608 2.095238e-02
R41974 n3_13833_18608 n3_13833_18764 9.904762e-02
R41975 n3_13833_18764 n3_13833_18791 1.714286e-02
R41976 n3_13833_18791 n3_13833_18824 2.095238e-02
R41977 n3_13833_18824 n3_13833_19007 1.161905e-01
R41978 n3_13833_19007 n3_13833_19040 2.095238e-02
R41979 n3_13833_19040 n3_13833_19223 1.161905e-01
R41980 n3_13833_19223 n3_13833_19256 2.095238e-02
R41981 n3_13833_19256 n3_13833_19404 9.396825e-02
R41982 n3_13833_19404 n3_13833_19412 5.079365e-03
R41983 n3_13833_19412 n3_13833_19439 1.714286e-02
R41984 n3_13833_19439 n3_13833_19472 2.095238e-02
R41985 n3_13833_19871 n3_13833_19904 2.095238e-02
R41986 n3_13833_19904 n3_13833_20087 1.161905e-01
R41987 n3_13833_20087 n3_13833_20120 2.095238e-02
R41988 n3_13833_20120 n3_13833_20303 1.161905e-01
R41989 n3_13833_20303 n3_13833_20336 2.095238e-02
R41990 n3_13833_20336 n3_13833_20519 1.161905e-01
R41991 n3_13833_20519 n3_13833_20552 2.095238e-02
R41992 n3_13833_20552 n3_13833_20674 7.746032e-02
R41993 n3_13833_20674 n3_13833_20687 8.253968e-03
R41994 n3_13833_20687 n3_13833_20735 3.047619e-02
R41995 n3_13833_20735 n3_13833_20768 2.095238e-02
R41996 n3_13833_20768 n3_13833_20770 1.269841e-03
R41997 n3_13833_20770 n3_13833_20951 1.149206e-01
R41998 n3_13833_20951 n3_13833_20984 2.095238e-02
R41999 n3_14021_215 n3_14021_248 2.095238e-02
R42000 n3_14021_248 n3_14021_383 8.571429e-02
R42001 n3_14021_383 n3_14021_424 2.603175e-02
R42002 n3_14021_424 n3_14021_431 4.444444e-03
R42003 n3_14021_520 n3_14021_647 8.063492e-02
R42004 n3_14021_647 n3_14021_680 2.095238e-02
R42005 n3_14021_680 n3_14021_863 1.161905e-01
R42006 n3_14021_863 n3_14021_896 2.095238e-02
R42007 n3_14021_896 n3_14021_1079 1.161905e-01
R42008 n3_14021_1079 n3_14021_1112 2.095238e-02
R42009 n3_14021_1112 n3_14021_1295 1.161905e-01
R42010 n3_14021_1295 n3_14021_1328 2.095238e-02
R42011 n3_14021_1328 n3_14021_1511 1.161905e-01
R42012 n3_14021_1511 n3_14021_1544 2.095238e-02
R42013 n3_14021_1544 n3_14021_1727 1.161905e-01
R42014 n3_14021_1727 n3_14021_1760 2.095238e-02
R42015 n3_14021_1760 n3_14021_1894 8.507937e-02
R42016 n3_14021_1894 n3_14021_1943 3.111111e-02
R42017 n3_14021_1943 n3_14021_1976 2.095238e-02
R42018 n3_14021_1976 n3_14021_2159 1.161905e-01
R42019 n3_14021_2159 n3_14021_2192 2.095238e-02
R42020 n3_14021_2192 n3_14021_2375 1.161905e-01
R42021 n3_14021_2375 n3_14021_2408 2.095238e-02
R42022 n3_14021_2408 n3_14021_2445 2.349206e-02
R42023 n3_14021_2445 n3_14021_2542 6.158730e-02
R42024 n3_14021_2542 n3_14021_2543 6.349206e-04
R42025 n3_14021_2543 n3_14021_2591 3.047619e-02
R42026 n3_14021_2591 n3_14021_2624 2.095238e-02
R42027 n3_14021_2624 n3_14021_2674 3.174603e-02
R42028 n3_14021_2770 n3_14021_2807 2.349206e-02
R42029 n3_14021_2807 n3_14021_2840 2.095238e-02
R42030 n3_14021_2840 n3_14021_2877 2.349206e-02
R42031 n3_14021_2877 n3_14021_2974 6.158730e-02
R42032 n3_14021_2974 n3_14021_3023 3.111111e-02
R42033 n3_14021_3023 n3_14021_3056 2.095238e-02
R42034 n3_14021_3056 n3_14021_3239 1.161905e-01
R42035 n3_14021_3239 n3_14021_3272 2.095238e-02
R42036 n3_14021_3272 n3_14021_3455 1.161905e-01
R42037 n3_14021_3455 n3_14021_3488 2.095238e-02
R42038 n3_14021_3488 n3_14021_3622 8.507937e-02
R42039 n3_14021_3622 n3_14021_3671 3.111111e-02
R42040 n3_14021_3671 n3_14021_3704 2.095238e-02
R42041 n3_14021_3704 n3_14021_3887 1.161905e-01
R42042 n3_14021_3887 n3_14021_3920 2.095238e-02
R42043 n3_14021_3920 n3_14021_4054 8.507937e-02
R42044 n3_14021_4054 n3_14021_4103 3.111111e-02
R42045 n3_14021_4103 n3_14021_4136 2.095238e-02
R42046 n3_14021_4136 n3_14021_4270 8.507937e-02
R42047 n3_14021_4270 n3_14021_4319 3.111111e-02
R42048 n3_14021_4319 n3_14021_4352 2.095238e-02
R42049 n3_14021_4352 n3_14021_4535 1.161905e-01
R42050 n3_14021_4535 n3_14021_4568 2.095238e-02
R42051 n3_14021_4568 n3_14021_4702 8.507937e-02
R42052 n3_14021_4702 n3_14021_4751 3.111111e-02
R42053 n3_14021_4751 n3_14021_4784 2.095238e-02
R42054 n3_14021_4784 n3_14021_4924 8.888889e-02
R42055 n3_14021_5000 n3_14021_5020 1.269841e-02
R42056 n3_14021_5020 n3_14021_5134 7.238095e-02
R42057 n3_14021_5134 n3_14021_5183 3.111111e-02
R42058 n3_14021_5183 n3_14021_5216 2.095238e-02
R42059 n3_14021_5216 n3_14021_5350 8.507937e-02
R42060 n3_14021_5350 n3_14021_5399 3.111111e-02
R42061 n3_14021_5399 n3_14021_5432 2.095238e-02
R42062 n3_14021_5432 n3_14021_5615 1.161905e-01
R42063 n3_14021_5615 n3_14021_5648 2.095238e-02
R42064 n3_14021_5648 n3_14021_5782 8.507937e-02
R42065 n3_14021_5782 n3_14021_5831 3.111111e-02
R42066 n3_14021_5831 n3_14021_5864 2.095238e-02
R42067 n3_14021_5864 n3_14021_6047 1.161905e-01
R42068 n3_14021_6047 n3_14021_6080 2.095238e-02
R42069 n3_14021_6080 n3_14021_6263 1.161905e-01
R42070 n3_14021_6263 n3_14021_6296 2.095238e-02
R42071 n3_14021_6296 n3_14021_6430 8.507937e-02
R42072 n3_14021_6430 n3_14021_6479 3.111111e-02
R42073 n3_14021_6479 n3_14021_6512 2.095238e-02
R42074 n3_14021_6512 n3_14021_6646 8.507937e-02
R42075 n3_14021_6646 n3_14021_6695 3.111111e-02
R42076 n3_14021_6695 n3_14021_6728 2.095238e-02
R42077 n3_14021_6728 n3_14021_6911 1.161905e-01
R42078 n3_14021_6911 n3_14021_6944 2.095238e-02
R42079 n3_14021_6944 n3_14021_7127 1.161905e-01
R42080 n3_14021_7127 n3_14021_7160 2.095238e-02
R42081 n3_14021_7160 n3_14021_7174 8.888889e-03
R42082 n3_14021_7270 n3_14021_7343 4.634921e-02
R42083 n3_14021_7343 n3_14021_7376 2.095238e-02
R42084 n3_14021_7376 n3_14021_7559 1.161905e-01
R42085 n3_14021_7559 n3_14021_7592 2.095238e-02
R42086 n3_14021_7592 n3_14021_7775 1.161905e-01
R42087 n3_14021_7775 n3_14021_7808 2.095238e-02
R42088 n3_14021_7808 n3_14021_7845 2.349206e-02
R42089 n3_14021_7845 n3_14021_7942 6.158730e-02
R42090 n3_14021_7942 n3_14021_7991 3.111111e-02
R42091 n3_14021_7991 n3_14021_8024 2.095238e-02
R42092 n3_14021_8024 n3_14021_8207 1.161905e-01
R42093 n3_14021_8207 n3_14021_8240 2.095238e-02
R42094 n3_14021_8240 n3_14021_8423 1.161905e-01
R42095 n3_14021_8423 n3_14021_8456 2.095238e-02
R42096 n3_14021_8456 n3_14021_8639 1.161905e-01
R42097 n3_14021_8639 n3_14021_8672 2.095238e-02
R42098 n3_14021_8672 n3_14021_8806 8.507937e-02
R42099 n3_14021_8806 n3_14021_8855 3.111111e-02
R42100 n3_14021_8855 n3_14021_8888 2.095238e-02
R42101 n3_14021_8888 n3_14021_8925 2.349206e-02
R42102 n3_14021_8925 n3_14021_9022 6.158730e-02
R42103 n3_14021_9022 n3_14021_9071 3.111111e-02
R42104 n3_14021_9071 n3_14021_9104 2.095238e-02
R42105 n3_14021_9104 n3_14021_9287 1.161905e-01
R42106 n3_14021_9287 n3_14021_9320 2.095238e-02
R42107 n3_14021_9320 n3_14021_9424 6.603175e-02
R42108 n3_14021_9503 n3_14021_9520 1.079365e-02
R42109 n3_14021_9520 n3_14021_9536 1.015873e-02
R42110 n3_14021_9536 n3_14021_9719 1.161905e-01
R42111 n3_14021_9719 n3_14021_9752 2.095238e-02
R42112 n3_14021_9752 n3_14021_9886 8.507937e-02
R42113 n3_14021_9886 n3_14021_9935 3.111111e-02
R42114 n3_14021_9935 n3_14021_9968 2.095238e-02
R42115 n3_14021_9968 n3_14021_10005 2.349206e-02
R42116 n3_14021_10005 n3_14021_10102 6.158730e-02
R42117 n3_14021_10102 n3_14021_10151 3.111111e-02
R42118 n3_14021_10151 n3_14021_10184 2.095238e-02
R42119 n3_14021_10184 n3_14021_10367 1.161905e-01
R42120 n3_14021_10367 n3_14021_10400 2.095238e-02
R42121 n3_14021_10616 n3_14021_10799 1.161905e-01
R42122 n3_14021_10799 n3_14021_10832 2.095238e-02
R42123 n3_14021_10832 n3_14021_10988 9.904762e-02
R42124 n3_14021_10988 n3_14021_11015 1.714286e-02
R42125 n3_14021_11015 n3_14021_11048 2.095238e-02
R42126 n3_14021_11048 n3_14021_11204 9.904762e-02
R42127 n3_14021_11204 n3_14021_11231 1.714286e-02
R42128 n3_14021_11231 n3_14021_11264 2.095238e-02
R42129 n3_14021_11264 n3_14021_11447 1.161905e-01
R42130 n3_14021_11447 n3_14021_11480 2.095238e-02
R42131 n3_14021_11480 n3_14021_11663 1.161905e-01
R42132 n3_14021_11663 n3_14021_11674 6.984127e-03
R42133 n3_14021_11674 n3_14021_11696 1.396825e-02
R42134 n3_14021_11770 n3_14021_11879 6.920635e-02
R42135 n3_14021_11879 n3_14021_11912 2.095238e-02
R42136 n3_14021_11912 n3_14021_12068 9.904762e-02
R42137 n3_14021_12068 n3_14021_12095 1.714286e-02
R42138 n3_14021_12095 n3_14021_12128 2.095238e-02
R42139 n3_14021_12128 n3_14021_12284 9.904762e-02
R42140 n3_14021_12284 n3_14021_12311 1.714286e-02
R42141 n3_14021_12311 n3_14021_12344 2.095238e-02
R42142 n3_14021_12344 n3_14021_12527 1.161905e-01
R42143 n3_14021_12527 n3_14021_12560 2.095238e-02
R42144 n3_14021_12560 n3_14021_12743 1.161905e-01
R42145 n3_14021_12743 n3_14021_12776 2.095238e-02
R42146 n3_14021_12776 n3_14021_12959 1.161905e-01
R42147 n3_14021_12959 n3_14021_12992 2.095238e-02
R42148 n3_14021_12992 n3_14021_13175 1.161905e-01
R42149 n3_14021_13175 n3_14021_13208 2.095238e-02
R42150 n3_14021_13208 n3_14021_13391 1.161905e-01
R42151 n3_14021_13391 n3_14021_13424 2.095238e-02
R42152 n3_14021_13424 n3_14021_13607 1.161905e-01
R42153 n3_14021_13607 n3_14021_13640 2.095238e-02
R42154 n3_14021_13640 n3_14021_13823 1.161905e-01
R42155 n3_14021_13823 n3_14021_13856 2.095238e-02
R42156 n3_14021_13856 n3_14021_13924 4.317460e-02
R42157 n3_14021_14020 n3_14021_14039 1.206349e-02
R42158 n3_14021_14039 n3_14021_14072 2.095238e-02
R42159 n3_14021_14072 n3_14021_14220 9.396825e-02
R42160 n3_14021_14220 n3_14021_14255 2.222222e-02
R42161 n3_14021_14255 n3_14021_14288 2.095238e-02
R42162 n3_14021_14288 n3_14021_14471 1.161905e-01
R42163 n3_14021_14471 n3_14021_14504 2.095238e-02
R42164 n3_14021_14504 n3_14021_14652 9.396825e-02
R42165 n3_14021_14652 n3_14021_14687 2.222222e-02
R42166 n3_14021_14687 n3_14021_14720 2.095238e-02
R42167 n3_14021_14720 n3_14021_14868 9.396825e-02
R42168 n3_14021_14868 n3_14021_14903 2.222222e-02
R42169 n3_14021_14903 n3_14021_14936 2.095238e-02
R42170 n3_14021_14936 n3_14021_15119 1.161905e-01
R42171 n3_14021_15119 n3_14021_15152 2.095238e-02
R42172 n3_14021_15152 n3_14021_15335 1.161905e-01
R42173 n3_14021_15335 n3_14021_15368 2.095238e-02
R42174 n3_14021_15368 n3_14021_15524 9.904762e-02
R42175 n3_14021_15524 n3_14021_15551 1.714286e-02
R42176 n3_14021_15551 n3_14021_15584 2.095238e-02
R42177 n3_14021_15584 n3_14021_15767 1.161905e-01
R42178 n3_14021_15767 n3_14021_15800 2.095238e-02
R42179 n3_14021_15800 n3_14021_15956 9.904762e-02
R42180 n3_14021_15956 n3_14021_15983 1.714286e-02
R42181 n3_14021_15983 n3_14021_16016 2.095238e-02
R42182 n3_14021_16016 n3_14021_16174 1.003175e-01
R42183 n3_14021_16174 n3_14021_16199 1.587302e-02
R42184 n3_14021_16270 n3_14021_16415 9.206349e-02
R42185 n3_14021_16415 n3_14021_16448 2.095238e-02
R42186 n3_14021_16448 n3_14021_16604 9.904762e-02
R42187 n3_14021_16604 n3_14021_16631 1.714286e-02
R42188 n3_14021_16631 n3_14021_16664 2.095238e-02
R42189 n3_14021_16664 n3_14021_16847 1.161905e-01
R42190 n3_14021_16847 n3_14021_16880 2.095238e-02
R42191 n3_14021_16880 n3_14021_17063 1.161905e-01
R42192 n3_14021_17063 n3_14021_17096 2.095238e-02
R42193 n3_14021_17096 n3_14021_17252 9.904762e-02
R42194 n3_14021_17252 n3_14021_17279 1.714286e-02
R42195 n3_14021_17279 n3_14021_17312 2.095238e-02
R42196 n3_14021_17312 n3_14021_17495 1.161905e-01
R42197 n3_14021_17495 n3_14021_17528 2.095238e-02
R42198 n3_14021_17528 n3_14021_17684 9.904762e-02
R42199 n3_14021_17684 n3_14021_17711 1.714286e-02
R42200 n3_14021_17711 n3_14021_17744 2.095238e-02
R42201 n3_14021_17744 n3_14021_17927 1.161905e-01
R42202 n3_14021_17927 n3_14021_17960 2.095238e-02
R42203 n3_14021_17960 n3_14021_18094 8.507937e-02
R42204 n3_14021_18094 n3_14021_18143 3.111111e-02
R42205 n3_14021_18143 n3_14021_18176 2.095238e-02
R42206 n3_14021_18176 n3_14021_18324 9.396825e-02
R42207 n3_14021_18324 n3_14021_18332 5.079365e-03
R42208 n3_14021_18332 n3_14021_18359 1.714286e-02
R42209 n3_14021_18359 n3_14021_18392 2.095238e-02
R42210 n3_14021_18392 n3_14021_18424 2.031746e-02
R42211 n3_14021_18520 n3_14021_18527 4.444444e-03
R42212 n3_14021_18527 n3_14021_18575 3.047619e-02
R42213 n3_14021_18575 n3_14021_18608 2.095238e-02
R42214 n3_14021_18608 n3_14021_18764 9.904762e-02
R42215 n3_14021_18764 n3_14021_18791 1.714286e-02
R42216 n3_14021_18791 n3_14021_18824 2.095238e-02
R42217 n3_14021_18824 n3_14021_19007 1.161905e-01
R42218 n3_14021_19007 n3_14021_19040 2.095238e-02
R42219 n3_14021_19040 n3_14021_19223 1.161905e-01
R42220 n3_14021_19223 n3_14021_19256 2.095238e-02
R42221 n3_14021_19256 n3_14021_19404 9.396825e-02
R42222 n3_14021_19404 n3_14021_19412 5.079365e-03
R42223 n3_14021_19412 n3_14021_19439 1.714286e-02
R42224 n3_14021_19439 n3_14021_19472 2.095238e-02
R42225 n3_14021_19472 n3_14021_19655 1.161905e-01
R42226 n3_14021_19655 n3_14021_19688 2.095238e-02
R42227 n3_14021_19688 n3_14021_19871 1.161905e-01
R42228 n3_14021_19871 n3_14021_19904 2.095238e-02
R42229 n3_14021_19904 n3_14021_20087 1.161905e-01
R42230 n3_14021_20087 n3_14021_20120 2.095238e-02
R42231 n3_14021_20120 n3_14021_20303 1.161905e-01
R42232 n3_14021_20303 n3_14021_20336 2.095238e-02
R42233 n3_14021_20336 n3_14021_20519 1.161905e-01
R42234 n3_14021_20519 n3_14021_20552 2.095238e-02
R42235 n3_14021_20552 n3_14021_20674 7.746032e-02
R42236 n3_14021_20674 n3_14021_20687 8.253968e-03
R42237 n3_14021_20768 n3_14021_20770 1.269841e-03
R42238 n3_14021_20770 n3_14021_20951 1.149206e-01
R42239 n3_14021_20951 n3_14021_20984 2.095238e-02
R42240 n3_14114_215 n3_14114_248 2.095238e-02
R42241 n3_14114_248 n3_14114_383 8.571429e-02
R42242 n3_14114_383 n3_14114_431 3.047619e-02
R42243 n3_14114_431 n3_14114_464 2.095238e-02
R42244 n3_14114_464 n3_14114_647 1.161905e-01
R42245 n3_14114_647 n3_14114_680 2.095238e-02
R42246 n3_14114_680 n3_14114_863 1.161905e-01
R42247 n3_14114_863 n3_14114_896 2.095238e-02
R42248 n3_14114_896 n3_14114_1079 1.161905e-01
R42249 n3_14114_1079 n3_14114_1112 2.095238e-02
R42250 n3_14114_1112 n3_14114_1295 1.161905e-01
R42251 n3_14114_1295 n3_14114_1328 2.095238e-02
R42252 n3_14114_1328 n3_14114_1511 1.161905e-01
R42253 n3_14114_1511 n3_14114_1544 2.095238e-02
R42254 n3_14114_1544 n3_14114_1727 1.161905e-01
R42255 n3_14114_1727 n3_14114_1760 2.095238e-02
R42256 n3_14114_1760 n3_14114_1894 8.507937e-02
R42257 n3_14114_1894 n3_14114_1943 3.111111e-02
R42258 n3_14114_1943 n3_14114_1976 2.095238e-02
R42259 n3_14114_1976 n3_14114_2159 1.161905e-01
R42260 n3_14114_2159 n3_14114_2192 2.095238e-02
R42261 n3_14114_2192 n3_14114_2375 1.161905e-01
R42262 n3_14114_2375 n3_14114_2408 2.095238e-02
R42263 n3_14114_2408 n3_14114_2445 2.349206e-02
R42264 n3_14114_2445 n3_14114_2542 6.158730e-02
R42265 n3_14114_2542 n3_14114_2543 6.349206e-04
R42266 n3_14114_2543 n3_14114_2591 3.047619e-02
R42267 n3_14114_2591 n3_14114_2624 2.095238e-02
R42268 n3_14114_18527 n3_14114_18575 3.047619e-02
R42269 n3_14114_18575 n3_14114_18608 2.095238e-02
R42270 n3_14114_18608 n3_14114_18764 9.904762e-02
R42271 n3_14114_18764 n3_14114_18791 1.714286e-02
R42272 n3_14114_18791 n3_14114_18824 2.095238e-02
R42273 n3_14114_18824 n3_14114_19007 1.161905e-01
R42274 n3_14114_19007 n3_14114_19040 2.095238e-02
R42275 n3_14114_19040 n3_14114_19223 1.161905e-01
R42276 n3_14114_19223 n3_14114_19256 2.095238e-02
R42277 n3_14114_19256 n3_14114_19404 9.396825e-02
R42278 n3_14114_19404 n3_14114_19439 2.222222e-02
R42279 n3_14114_19439 n3_14114_19472 2.095238e-02
R42280 n3_14114_19472 n3_14114_19655 1.161905e-01
R42281 n3_14114_19655 n3_14114_19688 2.095238e-02
R42282 n3_14114_19688 n3_14114_19871 1.161905e-01
R42283 n3_14114_19871 n3_14114_19904 2.095238e-02
R42284 n3_14114_19904 n3_14114_20087 1.161905e-01
R42285 n3_14114_20087 n3_14114_20120 2.095238e-02
R42286 n3_14114_20120 n3_14114_20303 1.161905e-01
R42287 n3_14114_20303 n3_14114_20336 2.095238e-02
R42288 n3_14114_20336 n3_14114_20519 1.161905e-01
R42289 n3_14114_20519 n3_14114_20552 2.095238e-02
R42290 n3_14114_20552 n3_14114_20687 8.571429e-02
R42291 n3_14114_20687 n3_14114_20735 3.047619e-02
R42292 n3_14114_20735 n3_14114_20768 2.095238e-02
R42293 n3_14114_20768 n3_14114_20951 1.161905e-01
R42294 n3_14114_20951 n3_14114_20984 2.095238e-02
R42295 n3_15900_215 n3_15900_248 2.095238e-02
R42296 n3_15900_248 n3_15900_383 8.571429e-02
R42297 n3_15900_383 n3_15900_431 3.047619e-02
R42298 n3_15900_431 n3_15900_464 2.095238e-02
R42299 n3_15900_464 n3_15900_647 1.161905e-01
R42300 n3_15900_647 n3_15900_680 2.095238e-02
R42301 n3_15900_680 n3_15900_863 1.161905e-01
R42302 n3_15900_863 n3_15900_896 2.095238e-02
R42303 n3_15900_896 n3_15900_1079 1.161905e-01
R42304 n3_15900_1079 n3_15900_1112 2.095238e-02
R42305 n3_15900_1112 n3_15900_1295 1.161905e-01
R42306 n3_15900_1295 n3_15900_1328 2.095238e-02
R42307 n3_15900_1328 n3_15900_1511 1.161905e-01
R42308 n3_15900_1511 n3_15900_1544 2.095238e-02
R42309 n3_15900_1544 n3_15900_1727 1.161905e-01
R42310 n3_15900_1727 n3_15900_1760 2.095238e-02
R42311 n3_15900_1760 n3_15900_1894 8.507937e-02
R42312 n3_15900_1894 n3_15900_1943 3.111111e-02
R42313 n3_15900_1943 n3_15900_1976 2.095238e-02
R42314 n3_15900_1976 n3_15900_2159 1.161905e-01
R42315 n3_15900_2159 n3_15900_2192 2.095238e-02
R42316 n3_15900_2192 n3_15900_2375 1.161905e-01
R42317 n3_15900_2375 n3_15900_2408 2.095238e-02
R42318 n3_15900_2408 n3_15900_2445 2.349206e-02
R42319 n3_15900_2445 n3_15900_2542 6.158730e-02
R42320 n3_15900_2542 n3_15900_2543 6.349206e-04
R42321 n3_15900_2543 n3_15900_2591 3.047619e-02
R42322 n3_15900_2591 n3_15900_2624 2.095238e-02
R42323 n3_15900_18527 n3_15900_18575 3.047619e-02
R42324 n3_15900_18575 n3_15900_18608 2.095238e-02
R42325 n3_15900_18608 n3_15900_18764 9.904762e-02
R42326 n3_15900_18764 n3_15900_18791 1.714286e-02
R42327 n3_15900_18791 n3_15900_18824 2.095238e-02
R42328 n3_15900_18824 n3_15900_19007 1.161905e-01
R42329 n3_15900_19007 n3_15900_19040 2.095238e-02
R42330 n3_15900_19040 n3_15900_19223 1.161905e-01
R42331 n3_15900_19223 n3_15900_19256 2.095238e-02
R42332 n3_15900_19256 n3_15900_19412 9.904762e-02
R42333 n3_15900_19412 n3_15900_19439 1.714286e-02
R42334 n3_15900_19439 n3_15900_19472 2.095238e-02
R42335 n3_15900_19472 n3_15900_19655 1.161905e-01
R42336 n3_15900_19655 n3_15900_19688 2.095238e-02
R42337 n3_15900_19688 n3_15900_19871 1.161905e-01
R42338 n3_15900_19871 n3_15900_19904 2.095238e-02
R42339 n3_15900_19904 n3_15900_20087 1.161905e-01
R42340 n3_15900_20087 n3_15900_20120 2.095238e-02
R42341 n3_15900_20120 n3_15900_20303 1.161905e-01
R42342 n3_15900_20303 n3_15900_20336 2.095238e-02
R42343 n3_15900_20336 n3_15900_20519 1.161905e-01
R42344 n3_15900_20519 n3_15900_20552 2.095238e-02
R42345 n3_15900_20552 n3_15900_20687 8.571429e-02
R42346 n3_15900_20687 n3_15900_20735 3.047619e-02
R42347 n3_15900_20735 n3_15900_20768 2.095238e-02
R42348 n3_15900_20768 n3_15900_20951 1.161905e-01
R42349 n3_15900_20951 n3_15900_20984 2.095238e-02
R42350 n3_16083_424 n3_16130_424 2.984127e-02
R42351 n3_16130_424 n3_16271_424 8.952381e-02
R42352 n3_16083_520 n3_16130_520 2.984127e-02
R42353 n3_16130_520 n3_16271_520 8.952381e-02
R42354 n3_16083_2674 n3_16130_2674 2.984127e-02
R42355 n3_16130_2674 n3_16271_2674 8.952381e-02
R42356 n3_16083_2770 n3_16130_2770 2.984127e-02
R42357 n3_16130_2770 n3_16271_2770 8.952381e-02
R42358 n3_16083_4924 n3_16130_4924 2.984127e-02
R42359 n3_16130_4924 n3_16271_4924 8.952381e-02
R42360 n3_16083_5020 n3_16130_5020 2.984127e-02
R42361 n3_16130_5020 n3_16271_5020 8.952381e-02
R42362 n3_16083_7174 n3_16130_7174 2.984127e-02
R42363 n3_16130_7174 n3_16271_7174 8.952381e-02
R42364 n3_16083_7270 n3_16130_7270 2.984127e-02
R42365 n3_16130_7270 n3_16271_7270 8.952381e-02
R42366 n3_16083_9424 n3_16130_9424 2.984127e-02
R42367 n3_16130_9424 n3_16271_9424 8.952381e-02
R42368 n3_16083_9520 n3_16130_9520 2.984127e-02
R42369 n3_16130_9520 n3_16271_9520 8.952381e-02
R42370 n3_16083_11674 n3_16130_11674 2.984127e-02
R42371 n3_16130_11674 n3_16271_11674 8.952381e-02
R42372 n3_16083_11770 n3_16130_11770 2.984127e-02
R42373 n3_16130_11770 n3_16271_11770 8.952381e-02
R42374 n3_16083_13924 n3_16130_13924 2.984127e-02
R42375 n3_16130_13924 n3_16271_13924 8.952381e-02
R42376 n3_16083_14020 n3_16130_14020 2.984127e-02
R42377 n3_16130_14020 n3_16271_14020 8.952381e-02
R42378 n3_16083_16174 n3_16130_16174 2.984127e-02
R42379 n3_16130_16174 n3_16271_16174 8.952381e-02
R42380 n3_16083_16270 n3_16130_16270 2.984127e-02
R42381 n3_16130_16270 n3_16271_16270 8.952381e-02
R42382 n3_16083_18424 n3_16130_18424 2.984127e-02
R42383 n3_16130_18424 n3_16271_18424 8.952381e-02
R42384 n3_16083_18520 n3_16130_18520 2.984127e-02
R42385 n3_16130_18520 n3_16271_18520 8.952381e-02
R42386 n3_16083_20674 n3_16130_20674 2.984127e-02
R42387 n3_16130_20674 n3_16271_20674 8.952381e-02
R42388 n3_16083_20770 n3_16130_20770 2.984127e-02
R42389 n3_16130_20770 n3_16271_20770 8.952381e-02
R42390 n3_16083_215 n3_16083_248 2.095238e-02
R42391 n3_16083_248 n3_16083_383 8.571429e-02
R42392 n3_16083_383 n3_16083_424 2.603175e-02
R42393 n3_16083_424 n3_16083_431 4.444444e-03
R42394 n3_16083_431 n3_16083_464 2.095238e-02
R42395 n3_16083_464 n3_16083_520 3.555556e-02
R42396 n3_16083_520 n3_16083_647 8.063492e-02
R42397 n3_16083_647 n3_16083_680 2.095238e-02
R42398 n3_16083_680 n3_16083_863 1.161905e-01
R42399 n3_16083_863 n3_16083_896 2.095238e-02
R42400 n3_16083_896 n3_16083_1079 1.161905e-01
R42401 n3_16083_1079 n3_16083_1112 2.095238e-02
R42402 n3_16083_1112 n3_16083_1295 1.161905e-01
R42403 n3_16083_1295 n3_16083_1328 2.095238e-02
R42404 n3_16083_1727 n3_16083_1760 2.095238e-02
R42405 n3_16083_1760 n3_16083_1894 8.507937e-02
R42406 n3_16083_1894 n3_16083_1943 3.111111e-02
R42407 n3_16083_1943 n3_16083_1976 2.095238e-02
R42408 n3_16083_1976 n3_16083_2159 1.161905e-01
R42409 n3_16083_2159 n3_16083_2192 2.095238e-02
R42410 n3_16083_2192 n3_16083_2375 1.161905e-01
R42411 n3_16083_2375 n3_16083_2408 2.095238e-02
R42412 n3_16083_2408 n3_16083_2445 2.349206e-02
R42413 n3_16083_2445 n3_16083_2542 6.158730e-02
R42414 n3_16083_2542 n3_16083_2543 6.349206e-04
R42415 n3_16083_2543 n3_16083_2591 3.047619e-02
R42416 n3_16083_2591 n3_16083_2624 2.095238e-02
R42417 n3_16083_2624 n3_16083_2674 3.174603e-02
R42418 n3_16083_2674 n3_16083_2770 6.095238e-02
R42419 n3_16083_2770 n3_16083_2807 2.349206e-02
R42420 n3_16083_2807 n3_16083_2840 2.095238e-02
R42421 n3_16083_2840 n3_16083_2877 2.349206e-02
R42422 n3_16083_2877 n3_16083_2974 6.158730e-02
R42423 n3_16083_2974 n3_16083_3023 3.111111e-02
R42424 n3_16083_3023 n3_16083_3056 2.095238e-02
R42425 n3_16083_3056 n3_16083_3239 1.161905e-01
R42426 n3_16083_3239 n3_16083_3272 2.095238e-02
R42427 n3_16083_3272 n3_16083_3406 8.507937e-02
R42428 n3_16083_3406 n3_16083_3455 3.111111e-02
R42429 n3_16083_3455 n3_16083_3488 2.095238e-02
R42430 n3_16083_3488 n3_16083_3671 1.161905e-01
R42431 n3_16083_3671 n3_16083_3704 2.095238e-02
R42432 n3_16083_4103 n3_16083_4136 2.095238e-02
R42433 n3_16083_4136 n3_16083_4319 1.161905e-01
R42434 n3_16083_4319 n3_16083_4352 2.095238e-02
R42435 n3_16083_4352 n3_16083_4486 8.507937e-02
R42436 n3_16083_4486 n3_16083_4535 3.111111e-02
R42437 n3_16083_4535 n3_16083_4568 2.095238e-02
R42438 n3_16083_4568 n3_16083_4702 8.507937e-02
R42439 n3_16083_4702 n3_16083_4751 3.111111e-02
R42440 n3_16083_4751 n3_16083_4784 2.095238e-02
R42441 n3_16083_4784 n3_16083_4919 8.571429e-02
R42442 n3_16083_4919 n3_16083_4924 3.174603e-03
R42443 n3_16083_4924 n3_16083_4967 2.730159e-02
R42444 n3_16083_4967 n3_16083_5000 2.095238e-02
R42445 n3_16083_5000 n3_16083_5020 1.269841e-02
R42446 n3_16083_5020 n3_16083_5134 7.238095e-02
R42447 n3_16083_5134 n3_16083_5183 3.111111e-02
R42448 n3_16083_5183 n3_16083_5216 2.095238e-02
R42449 n3_16083_5216 n3_16083_5253 2.349206e-02
R42450 n3_16083_5253 n3_16083_5350 6.158730e-02
R42451 n3_16083_5350 n3_16083_5399 3.111111e-02
R42452 n3_16083_5399 n3_16083_5432 2.095238e-02
R42453 n3_16083_5432 n3_16083_5566 8.507937e-02
R42454 n3_16083_5566 n3_16083_5615 3.111111e-02
R42455 n3_16083_5615 n3_16083_5648 2.095238e-02
R42456 n3_16083_5648 n3_16083_5831 1.161905e-01
R42457 n3_16083_5831 n3_16083_5864 2.095238e-02
R42458 n3_16083_6263 n3_16083_6296 2.095238e-02
R42459 n3_16083_6296 n3_16083_6333 2.349206e-02
R42460 n3_16083_6333 n3_16083_6430 6.158730e-02
R42461 n3_16083_6430 n3_16083_6479 3.111111e-02
R42462 n3_16083_6479 n3_16083_6512 2.095238e-02
R42463 n3_16083_6512 n3_16083_6695 1.161905e-01
R42464 n3_16083_6695 n3_16083_6728 2.095238e-02
R42465 n3_16083_6728 n3_16083_6911 1.161905e-01
R42466 n3_16083_6911 n3_16083_6944 2.095238e-02
R42467 n3_16083_6944 n3_16083_7127 1.161905e-01
R42468 n3_16083_7127 n3_16083_7160 2.095238e-02
R42469 n3_16083_7160 n3_16083_7174 8.888889e-03
R42470 n3_16083_7174 n3_16083_7270 6.095238e-02
R42471 n3_16083_7270 n3_16083_7343 4.634921e-02
R42472 n3_16083_7343 n3_16083_7376 2.095238e-02
R42473 n3_16083_7376 n3_16083_7559 1.161905e-01
R42474 n3_16083_7559 n3_16083_7592 2.095238e-02
R42475 n3_16083_7592 n3_16083_7775 1.161905e-01
R42476 n3_16083_7775 n3_16083_7808 2.095238e-02
R42477 n3_16083_7808 n3_16083_7845 2.349206e-02
R42478 n3_16083_7845 n3_16083_7942 6.158730e-02
R42479 n3_16083_7942 n3_16083_7991 3.111111e-02
R42480 n3_16083_7991 n3_16083_8024 2.095238e-02
R42481 n3_16083_8024 n3_16083_8207 1.161905e-01
R42482 n3_16083_8207 n3_16083_8240 2.095238e-02
R42483 n3_16083_8456 n3_16083_8639 1.161905e-01
R42484 n3_16083_8639 n3_16083_8672 2.095238e-02
R42485 n3_16083_8672 n3_16083_8855 1.161905e-01
R42486 n3_16083_8855 n3_16083_8888 2.095238e-02
R42487 n3_16083_8888 n3_16083_8925 2.349206e-02
R42488 n3_16083_8925 n3_16083_9022 6.158730e-02
R42489 n3_16083_9022 n3_16083_9071 3.111111e-02
R42490 n3_16083_9071 n3_16083_9104 2.095238e-02
R42491 n3_16083_9104 n3_16083_9287 1.161905e-01
R42492 n3_16083_9287 n3_16083_9320 2.095238e-02
R42493 n3_16083_9320 n3_16083_9424 6.603175e-02
R42494 n3_16083_9424 n3_16083_9503 5.015873e-02
R42495 n3_16083_9503 n3_16083_9520 1.079365e-02
R42496 n3_16083_9520 n3_16083_9536 1.015873e-02
R42497 n3_16083_9536 n3_16083_9719 1.161905e-01
R42498 n3_16083_9719 n3_16083_9752 2.095238e-02
R42499 n3_16083_9752 n3_16083_9935 1.161905e-01
R42500 n3_16083_9935 n3_16083_9968 2.095238e-02
R42501 n3_16083_9968 n3_16083_10005 2.349206e-02
R42502 n3_16083_10005 n3_16083_10102 6.158730e-02
R42503 n3_16083_10102 n3_16083_10151 3.111111e-02
R42504 n3_16083_10151 n3_16083_10184 2.095238e-02
R42505 n3_16083_10184 n3_16083_10367 1.161905e-01
R42506 n3_16083_10367 n3_16083_10400 2.095238e-02
R42507 n3_16083_10799 n3_16083_10832 2.095238e-02
R42508 n3_16083_10832 n3_16083_11015 1.161905e-01
R42509 n3_16083_11015 n3_16083_11048 2.095238e-02
R42510 n3_16083_11048 n3_16083_11196 9.396825e-02
R42511 n3_16083_11196 n3_16083_11204 5.079365e-03
R42512 n3_16083_11204 n3_16083_11231 1.714286e-02
R42513 n3_16083_11231 n3_16083_11264 2.095238e-02
R42514 n3_16083_11264 n3_16083_11447 1.161905e-01
R42515 n3_16083_11447 n3_16083_11480 2.095238e-02
R42516 n3_16083_11480 n3_16083_11663 1.161905e-01
R42517 n3_16083_11663 n3_16083_11674 6.984127e-03
R42518 n3_16083_11674 n3_16083_11696 1.396825e-02
R42519 n3_16083_11696 n3_16083_11770 4.698413e-02
R42520 n3_16083_11770 n3_16083_11879 6.920635e-02
R42521 n3_16083_11879 n3_16083_11912 2.095238e-02
R42522 n3_16083_11912 n3_16083_12095 1.161905e-01
R42523 n3_16083_12095 n3_16083_12128 2.095238e-02
R42524 n3_16083_12128 n3_16083_12276 9.396825e-02
R42525 n3_16083_12276 n3_16083_12284 5.079365e-03
R42526 n3_16083_12284 n3_16083_12311 1.714286e-02
R42527 n3_16083_12311 n3_16083_12344 2.095238e-02
R42528 n3_16083_12344 n3_16083_12527 1.161905e-01
R42529 n3_16083_12527 n3_16083_12560 2.095238e-02
R42530 n3_16083_12560 n3_16083_12743 1.161905e-01
R42531 n3_16083_12959 n3_16083_12992 2.095238e-02
R42532 n3_16083_12992 n3_16083_13175 1.161905e-01
R42533 n3_16083_13175 n3_16083_13208 2.095238e-02
R42534 n3_16083_13208 n3_16083_13391 1.161905e-01
R42535 n3_16083_13391 n3_16083_13424 2.095238e-02
R42536 n3_16083_13424 n3_16083_13607 1.161905e-01
R42537 n3_16083_13607 n3_16083_13640 2.095238e-02
R42538 n3_16083_13640 n3_16083_13788 9.396825e-02
R42539 n3_16083_13788 n3_16083_13823 2.222222e-02
R42540 n3_16083_13823 n3_16083_13856 2.095238e-02
R42541 n3_16083_13856 n3_16083_13924 4.317460e-02
R42542 n3_16083_13924 n3_16083_14020 6.095238e-02
R42543 n3_16083_14020 n3_16083_14039 1.206349e-02
R42544 n3_16083_14039 n3_16083_14072 2.095238e-02
R42545 n3_16083_14072 n3_16083_14255 1.161905e-01
R42546 n3_16083_14255 n3_16083_14288 2.095238e-02
R42547 n3_16083_14288 n3_16083_14471 1.161905e-01
R42548 n3_16083_14471 n3_16083_14504 2.095238e-02
R42549 n3_16083_14504 n3_16083_14652 9.396825e-02
R42550 n3_16083_14652 n3_16083_14687 2.222222e-02
R42551 n3_16083_14687 n3_16083_14720 2.095238e-02
R42552 n3_16083_14720 n3_16083_14903 1.161905e-01
R42553 n3_16083_14903 n3_16083_14936 2.095238e-02
R42554 n3_16083_15300 n3_16083_15335 2.222222e-02
R42555 n3_16083_15335 n3_16083_15368 2.095238e-02
R42556 n3_16083_15368 n3_16083_15551 1.161905e-01
R42557 n3_16083_15551 n3_16083_15584 2.095238e-02
R42558 n3_16083_15584 n3_16083_15740 9.904762e-02
R42559 n3_16083_15740 n3_16083_15767 1.714286e-02
R42560 n3_16083_15767 n3_16083_15800 2.095238e-02
R42561 n3_16083_15800 n3_16083_15983 1.161905e-01
R42562 n3_16083_15983 n3_16083_16016 2.095238e-02
R42563 n3_16083_16016 n3_16083_16174 1.003175e-01
R42564 n3_16083_16174 n3_16083_16199 1.587302e-02
R42565 n3_16083_16199 n3_16083_16232 2.095238e-02
R42566 n3_16083_16232 n3_16083_16270 2.412698e-02
R42567 n3_16083_16270 n3_16083_16415 9.206349e-02
R42568 n3_16083_16415 n3_16083_16448 2.095238e-02
R42569 n3_16083_16448 n3_16083_16604 9.904762e-02
R42570 n3_16083_16604 n3_16083_16631 1.714286e-02
R42571 n3_16083_16631 n3_16083_16664 2.095238e-02
R42572 n3_16083_16664 n3_16083_16798 8.507937e-02
R42573 n3_16083_16798 n3_16083_16820 1.396825e-02
R42574 n3_16083_16820 n3_16083_16847 1.714286e-02
R42575 n3_16083_16847 n3_16083_16880 2.095238e-02
R42576 n3_16083_16880 n3_16083_17063 1.161905e-01
R42577 n3_16083_17063 n3_16083_17096 2.095238e-02
R42578 n3_16083_17495 n3_16083_17528 2.095238e-02
R42579 n3_16083_17528 n3_16083_17676 9.396825e-02
R42580 n3_16083_17676 n3_16083_17684 5.079365e-03
R42581 n3_16083_17684 n3_16083_17711 1.714286e-02
R42582 n3_16083_17711 n3_16083_17744 2.095238e-02
R42583 n3_16083_17744 n3_16083_17927 1.161905e-01
R42584 n3_16083_17927 n3_16083_17960 2.095238e-02
R42585 n3_16083_17960 n3_16083_18143 1.161905e-01
R42586 n3_16083_18143 n3_16083_18176 2.095238e-02
R42587 n3_16083_18176 n3_16083_18332 9.904762e-02
R42588 n3_16083_18332 n3_16083_18359 1.714286e-02
R42589 n3_16083_18359 n3_16083_18392 2.095238e-02
R42590 n3_16083_18392 n3_16083_18424 2.031746e-02
R42591 n3_16083_18424 n3_16083_18520 6.095238e-02
R42592 n3_16083_18520 n3_16083_18527 4.444444e-03
R42593 n3_16083_18527 n3_16083_18575 3.047619e-02
R42594 n3_16083_18575 n3_16083_18608 2.095238e-02
R42595 n3_16083_18608 n3_16083_18764 9.904762e-02
R42596 n3_16083_18764 n3_16083_18791 1.714286e-02
R42597 n3_16083_18791 n3_16083_18824 2.095238e-02
R42598 n3_16083_18824 n3_16083_19007 1.161905e-01
R42599 n3_16083_19007 n3_16083_19040 2.095238e-02
R42600 n3_16083_19040 n3_16083_19196 9.904762e-02
R42601 n3_16083_19196 n3_16083_19223 1.714286e-02
R42602 n3_16083_19223 n3_16083_19256 2.095238e-02
R42603 n3_16083_19256 n3_16083_19412 9.904762e-02
R42604 n3_16083_19412 n3_16083_19439 1.714286e-02
R42605 n3_16083_19439 n3_16083_19472 2.095238e-02
R42606 n3_16083_19871 n3_16083_19904 2.095238e-02
R42607 n3_16083_19904 n3_16083_20087 1.161905e-01
R42608 n3_16083_20087 n3_16083_20120 2.095238e-02
R42609 n3_16083_20120 n3_16083_20303 1.161905e-01
R42610 n3_16083_20303 n3_16083_20336 2.095238e-02
R42611 n3_16083_20336 n3_16083_20519 1.161905e-01
R42612 n3_16083_20519 n3_16083_20552 2.095238e-02
R42613 n3_16083_20552 n3_16083_20674 7.746032e-02
R42614 n3_16083_20674 n3_16083_20687 8.253968e-03
R42615 n3_16083_20687 n3_16083_20735 3.047619e-02
R42616 n3_16083_20735 n3_16083_20768 2.095238e-02
R42617 n3_16083_20768 n3_16083_20770 1.269841e-03
R42618 n3_16083_20770 n3_16083_20951 1.149206e-01
R42619 n3_16083_20951 n3_16083_20984 2.095238e-02
R42620 n3_16271_215 n3_16271_248 2.095238e-02
R42621 n3_16271_248 n3_16271_383 8.571429e-02
R42622 n3_16271_383 n3_16271_424 2.603175e-02
R42623 n3_16271_424 n3_16271_431 4.444444e-03
R42624 n3_16271_520 n3_16271_647 8.063492e-02
R42625 n3_16271_647 n3_16271_680 2.095238e-02
R42626 n3_16271_680 n3_16271_863 1.161905e-01
R42627 n3_16271_863 n3_16271_896 2.095238e-02
R42628 n3_16271_896 n3_16271_1079 1.161905e-01
R42629 n3_16271_1079 n3_16271_1112 2.095238e-02
R42630 n3_16271_1112 n3_16271_1295 1.161905e-01
R42631 n3_16271_1295 n3_16271_1328 2.095238e-02
R42632 n3_16271_1328 n3_16271_1511 1.161905e-01
R42633 n3_16271_1511 n3_16271_1544 2.095238e-02
R42634 n3_16271_1544 n3_16271_1727 1.161905e-01
R42635 n3_16271_1727 n3_16271_1760 2.095238e-02
R42636 n3_16271_1760 n3_16271_1894 8.507937e-02
R42637 n3_16271_1894 n3_16271_1943 3.111111e-02
R42638 n3_16271_1943 n3_16271_1976 2.095238e-02
R42639 n3_16271_1976 n3_16271_2159 1.161905e-01
R42640 n3_16271_2159 n3_16271_2192 2.095238e-02
R42641 n3_16271_2192 n3_16271_2375 1.161905e-01
R42642 n3_16271_2375 n3_16271_2408 2.095238e-02
R42643 n3_16271_2408 n3_16271_2445 2.349206e-02
R42644 n3_16271_2445 n3_16271_2542 6.158730e-02
R42645 n3_16271_2542 n3_16271_2543 6.349206e-04
R42646 n3_16271_2543 n3_16271_2591 3.047619e-02
R42647 n3_16271_2591 n3_16271_2624 2.095238e-02
R42648 n3_16271_2624 n3_16271_2674 3.174603e-02
R42649 n3_16271_2770 n3_16271_2807 2.349206e-02
R42650 n3_16271_2807 n3_16271_2840 2.095238e-02
R42651 n3_16271_2840 n3_16271_2877 2.349206e-02
R42652 n3_16271_2877 n3_16271_2974 6.158730e-02
R42653 n3_16271_2974 n3_16271_3023 3.111111e-02
R42654 n3_16271_3023 n3_16271_3056 2.095238e-02
R42655 n3_16271_3056 n3_16271_3239 1.161905e-01
R42656 n3_16271_3239 n3_16271_3272 2.095238e-02
R42657 n3_16271_3272 n3_16271_3406 8.507937e-02
R42658 n3_16271_3406 n3_16271_3455 3.111111e-02
R42659 n3_16271_3455 n3_16271_3488 2.095238e-02
R42660 n3_16271_3488 n3_16271_3671 1.161905e-01
R42661 n3_16271_3671 n3_16271_3704 2.095238e-02
R42662 n3_16271_3704 n3_16271_3887 1.161905e-01
R42663 n3_16271_3887 n3_16271_3920 2.095238e-02
R42664 n3_16271_3920 n3_16271_4103 1.161905e-01
R42665 n3_16271_4103 n3_16271_4136 2.095238e-02
R42666 n3_16271_4136 n3_16271_4319 1.161905e-01
R42667 n3_16271_4319 n3_16271_4352 2.095238e-02
R42668 n3_16271_4352 n3_16271_4486 8.507937e-02
R42669 n3_16271_4486 n3_16271_4535 3.111111e-02
R42670 n3_16271_4535 n3_16271_4568 2.095238e-02
R42671 n3_16271_4568 n3_16271_4702 8.507937e-02
R42672 n3_16271_4702 n3_16271_4751 3.111111e-02
R42673 n3_16271_4751 n3_16271_4784 2.095238e-02
R42674 n3_16271_4784 n3_16271_4919 8.571429e-02
R42675 n3_16271_4919 n3_16271_4924 3.174603e-03
R42676 n3_16271_5000 n3_16271_5020 1.269841e-02
R42677 n3_16271_5020 n3_16271_5134 7.238095e-02
R42678 n3_16271_5134 n3_16271_5183 3.111111e-02
R42679 n3_16271_5183 n3_16271_5216 2.095238e-02
R42680 n3_16271_5216 n3_16271_5253 2.349206e-02
R42681 n3_16271_5253 n3_16271_5350 6.158730e-02
R42682 n3_16271_5350 n3_16271_5399 3.111111e-02
R42683 n3_16271_5399 n3_16271_5432 2.095238e-02
R42684 n3_16271_5432 n3_16271_5566 8.507937e-02
R42685 n3_16271_5566 n3_16271_5615 3.111111e-02
R42686 n3_16271_5615 n3_16271_5648 2.095238e-02
R42687 n3_16271_5648 n3_16271_5831 1.161905e-01
R42688 n3_16271_5831 n3_16271_5864 2.095238e-02
R42689 n3_16271_5864 n3_16271_6047 1.161905e-01
R42690 n3_16271_6047 n3_16271_6080 2.095238e-02
R42691 n3_16271_6080 n3_16271_6263 1.161905e-01
R42692 n3_16271_6263 n3_16271_6296 2.095238e-02
R42693 n3_16271_6296 n3_16271_6333 2.349206e-02
R42694 n3_16271_6333 n3_16271_6430 6.158730e-02
R42695 n3_16271_6430 n3_16271_6479 3.111111e-02
R42696 n3_16271_6479 n3_16271_6512 2.095238e-02
R42697 n3_16271_6512 n3_16271_6695 1.161905e-01
R42698 n3_16271_6695 n3_16271_6728 2.095238e-02
R42699 n3_16271_6728 n3_16271_6911 1.161905e-01
R42700 n3_16271_6911 n3_16271_6944 2.095238e-02
R42701 n3_16271_6944 n3_16271_7127 1.161905e-01
R42702 n3_16271_7127 n3_16271_7160 2.095238e-02
R42703 n3_16271_7160 n3_16271_7174 8.888889e-03
R42704 n3_16271_7270 n3_16271_7343 4.634921e-02
R42705 n3_16271_7343 n3_16271_7376 2.095238e-02
R42706 n3_16271_7376 n3_16271_7559 1.161905e-01
R42707 n3_16271_7559 n3_16271_7592 2.095238e-02
R42708 n3_16271_7592 n3_16271_7775 1.161905e-01
R42709 n3_16271_7775 n3_16271_7808 2.095238e-02
R42710 n3_16271_7808 n3_16271_7845 2.349206e-02
R42711 n3_16271_7845 n3_16271_7942 6.158730e-02
R42712 n3_16271_7942 n3_16271_7991 3.111111e-02
R42713 n3_16271_7991 n3_16271_8024 2.095238e-02
R42714 n3_16271_8024 n3_16271_8207 1.161905e-01
R42715 n3_16271_8207 n3_16271_8240 2.095238e-02
R42716 n3_16271_8240 n3_16271_8423 1.161905e-01
R42717 n3_16271_8423 n3_16271_8456 2.095238e-02
R42718 n3_16271_8456 n3_16271_8639 1.161905e-01
R42719 n3_16271_8639 n3_16271_8672 2.095238e-02
R42720 n3_16271_8672 n3_16271_8855 1.161905e-01
R42721 n3_16271_8855 n3_16271_8888 2.095238e-02
R42722 n3_16271_8888 n3_16271_8925 2.349206e-02
R42723 n3_16271_8925 n3_16271_9022 6.158730e-02
R42724 n3_16271_9022 n3_16271_9071 3.111111e-02
R42725 n3_16271_9071 n3_16271_9104 2.095238e-02
R42726 n3_16271_9104 n3_16271_9287 1.161905e-01
R42727 n3_16271_9287 n3_16271_9320 2.095238e-02
R42728 n3_16271_9320 n3_16271_9424 6.603175e-02
R42729 n3_16271_9503 n3_16271_9520 1.079365e-02
R42730 n3_16271_9520 n3_16271_9536 1.015873e-02
R42731 n3_16271_9536 n3_16271_9719 1.161905e-01
R42732 n3_16271_9719 n3_16271_9752 2.095238e-02
R42733 n3_16271_9752 n3_16271_9935 1.161905e-01
R42734 n3_16271_9935 n3_16271_9968 2.095238e-02
R42735 n3_16271_9968 n3_16271_10005 2.349206e-02
R42736 n3_16271_10005 n3_16271_10102 6.158730e-02
R42737 n3_16271_10102 n3_16271_10151 3.111111e-02
R42738 n3_16271_10151 n3_16271_10184 2.095238e-02
R42739 n3_16271_10184 n3_16271_10367 1.161905e-01
R42740 n3_16271_10367 n3_16271_10400 2.095238e-02
R42741 n3_16271_10616 n3_16271_10799 1.161905e-01
R42742 n3_16271_10799 n3_16271_10832 2.095238e-02
R42743 n3_16271_10832 n3_16271_11015 1.161905e-01
R42744 n3_16271_11015 n3_16271_11048 2.095238e-02
R42745 n3_16271_11048 n3_16271_11196 9.396825e-02
R42746 n3_16271_11196 n3_16271_11204 5.079365e-03
R42747 n3_16271_11204 n3_16271_11231 1.714286e-02
R42748 n3_16271_11231 n3_16271_11264 2.095238e-02
R42749 n3_16271_11264 n3_16271_11447 1.161905e-01
R42750 n3_16271_11447 n3_16271_11480 2.095238e-02
R42751 n3_16271_11480 n3_16271_11663 1.161905e-01
R42752 n3_16271_11663 n3_16271_11674 6.984127e-03
R42753 n3_16271_11674 n3_16271_11696 1.396825e-02
R42754 n3_16271_11770 n3_16271_11879 6.920635e-02
R42755 n3_16271_11879 n3_16271_11912 2.095238e-02
R42756 n3_16271_11912 n3_16271_12095 1.161905e-01
R42757 n3_16271_12095 n3_16271_12128 2.095238e-02
R42758 n3_16271_12128 n3_16271_12276 9.396825e-02
R42759 n3_16271_12276 n3_16271_12284 5.079365e-03
R42760 n3_16271_12284 n3_16271_12311 1.714286e-02
R42761 n3_16271_12311 n3_16271_12344 2.095238e-02
R42762 n3_16271_12344 n3_16271_12527 1.161905e-01
R42763 n3_16271_12527 n3_16271_12560 2.095238e-02
R42764 n3_16271_12560 n3_16271_12743 1.161905e-01
R42765 n3_16271_12743 n3_16271_12776 2.095238e-02
R42766 n3_16271_12776 n3_16271_12959 1.161905e-01
R42767 n3_16271_12959 n3_16271_12992 2.095238e-02
R42768 n3_16271_12992 n3_16271_13175 1.161905e-01
R42769 n3_16271_13175 n3_16271_13208 2.095238e-02
R42770 n3_16271_13208 n3_16271_13391 1.161905e-01
R42771 n3_16271_13391 n3_16271_13424 2.095238e-02
R42772 n3_16271_13424 n3_16271_13607 1.161905e-01
R42773 n3_16271_13607 n3_16271_13640 2.095238e-02
R42774 n3_16271_13640 n3_16271_13788 9.396825e-02
R42775 n3_16271_13788 n3_16271_13823 2.222222e-02
R42776 n3_16271_13823 n3_16271_13856 2.095238e-02
R42777 n3_16271_13856 n3_16271_13924 4.317460e-02
R42778 n3_16271_14020 n3_16271_14039 1.206349e-02
R42779 n3_16271_14039 n3_16271_14072 2.095238e-02
R42780 n3_16271_14072 n3_16271_14255 1.161905e-01
R42781 n3_16271_14255 n3_16271_14288 2.095238e-02
R42782 n3_16271_14288 n3_16271_14471 1.161905e-01
R42783 n3_16271_14471 n3_16271_14504 2.095238e-02
R42784 n3_16271_14504 n3_16271_14652 9.396825e-02
R42785 n3_16271_14652 n3_16271_14687 2.222222e-02
R42786 n3_16271_14687 n3_16271_14720 2.095238e-02
R42787 n3_16271_14720 n3_16271_14903 1.161905e-01
R42788 n3_16271_14903 n3_16271_14936 2.095238e-02
R42789 n3_16271_14936 n3_16271_15084 9.396825e-02
R42790 n3_16271_15084 n3_16271_15119 2.222222e-02
R42791 n3_16271_15119 n3_16271_15152 2.095238e-02
R42792 n3_16271_15152 n3_16271_15300 9.396825e-02
R42793 n3_16271_15300 n3_16271_15335 2.222222e-02
R42794 n3_16271_15335 n3_16271_15368 2.095238e-02
R42795 n3_16271_15368 n3_16271_15551 1.161905e-01
R42796 n3_16271_15551 n3_16271_15584 2.095238e-02
R42797 n3_16271_15584 n3_16271_15740 9.904762e-02
R42798 n3_16271_15740 n3_16271_15767 1.714286e-02
R42799 n3_16271_15767 n3_16271_15800 2.095238e-02
R42800 n3_16271_15800 n3_16271_15983 1.161905e-01
R42801 n3_16271_15983 n3_16271_16016 2.095238e-02
R42802 n3_16271_16016 n3_16271_16174 1.003175e-01
R42803 n3_16271_16174 n3_16271_16199 1.587302e-02
R42804 n3_16271_16270 n3_16271_16415 9.206349e-02
R42805 n3_16271_16415 n3_16271_16448 2.095238e-02
R42806 n3_16271_16448 n3_16271_16604 9.904762e-02
R42807 n3_16271_16604 n3_16271_16631 1.714286e-02
R42808 n3_16271_16631 n3_16271_16664 2.095238e-02
R42809 n3_16271_16664 n3_16271_16798 8.507937e-02
R42810 n3_16271_16798 n3_16271_16820 1.396825e-02
R42811 n3_16271_16820 n3_16271_16847 1.714286e-02
R42812 n3_16271_16847 n3_16271_16880 2.095238e-02
R42813 n3_16271_16880 n3_16271_17063 1.161905e-01
R42814 n3_16271_17063 n3_16271_17096 2.095238e-02
R42815 n3_16271_17096 n3_16271_17252 9.904762e-02
R42816 n3_16271_17252 n3_16271_17279 1.714286e-02
R42817 n3_16271_17279 n3_16271_17312 2.095238e-02
R42818 n3_16271_17312 n3_16271_17495 1.161905e-01
R42819 n3_16271_17495 n3_16271_17528 2.095238e-02
R42820 n3_16271_17528 n3_16271_17676 9.396825e-02
R42821 n3_16271_17676 n3_16271_17684 5.079365e-03
R42822 n3_16271_17684 n3_16271_17711 1.714286e-02
R42823 n3_16271_17711 n3_16271_17744 2.095238e-02
R42824 n3_16271_17744 n3_16271_17927 1.161905e-01
R42825 n3_16271_17927 n3_16271_17960 2.095238e-02
R42826 n3_16271_17960 n3_16271_18143 1.161905e-01
R42827 n3_16271_18143 n3_16271_18176 2.095238e-02
R42828 n3_16271_18176 n3_16271_18332 9.904762e-02
R42829 n3_16271_18332 n3_16271_18359 1.714286e-02
R42830 n3_16271_18359 n3_16271_18392 2.095238e-02
R42831 n3_16271_18392 n3_16271_18424 2.031746e-02
R42832 n3_16271_18520 n3_16271_18527 4.444444e-03
R42833 n3_16271_18527 n3_16271_18575 3.047619e-02
R42834 n3_16271_18575 n3_16271_18608 2.095238e-02
R42835 n3_16271_18608 n3_16271_18764 9.904762e-02
R42836 n3_16271_18764 n3_16271_18791 1.714286e-02
R42837 n3_16271_18791 n3_16271_18824 2.095238e-02
R42838 n3_16271_18824 n3_16271_19007 1.161905e-01
R42839 n3_16271_19007 n3_16271_19040 2.095238e-02
R42840 n3_16271_19040 n3_16271_19196 9.904762e-02
R42841 n3_16271_19196 n3_16271_19223 1.714286e-02
R42842 n3_16271_19223 n3_16271_19256 2.095238e-02
R42843 n3_16271_19256 n3_16271_19412 9.904762e-02
R42844 n3_16271_19412 n3_16271_19439 1.714286e-02
R42845 n3_16271_19439 n3_16271_19472 2.095238e-02
R42846 n3_16271_19472 n3_16271_19655 1.161905e-01
R42847 n3_16271_19655 n3_16271_19688 2.095238e-02
R42848 n3_16271_19688 n3_16271_19871 1.161905e-01
R42849 n3_16271_19871 n3_16271_19904 2.095238e-02
R42850 n3_16271_19904 n3_16271_20087 1.161905e-01
R42851 n3_16271_20087 n3_16271_20120 2.095238e-02
R42852 n3_16271_20120 n3_16271_20303 1.161905e-01
R42853 n3_16271_20303 n3_16271_20336 2.095238e-02
R42854 n3_16271_20336 n3_16271_20519 1.161905e-01
R42855 n3_16271_20519 n3_16271_20552 2.095238e-02
R42856 n3_16271_20552 n3_16271_20674 7.746032e-02
R42857 n3_16271_20674 n3_16271_20687 8.253968e-03
R42858 n3_16271_20768 n3_16271_20770 1.269841e-03
R42859 n3_16271_20770 n3_16271_20951 1.149206e-01
R42860 n3_16271_20951 n3_16271_20984 2.095238e-02
R42861 n3_16364_215 n3_16364_248 2.095238e-02
R42862 n3_16364_248 n3_16364_383 8.571429e-02
R42863 n3_16364_383 n3_16364_431 3.047619e-02
R42864 n3_16364_431 n3_16364_464 2.095238e-02
R42865 n3_16364_464 n3_16364_647 1.161905e-01
R42866 n3_16364_647 n3_16364_680 2.095238e-02
R42867 n3_16364_680 n3_16364_863 1.161905e-01
R42868 n3_16364_863 n3_16364_896 2.095238e-02
R42869 n3_16364_896 n3_16364_1079 1.161905e-01
R42870 n3_16364_1079 n3_16364_1112 2.095238e-02
R42871 n3_16364_1112 n3_16364_1295 1.161905e-01
R42872 n3_16364_1295 n3_16364_1328 2.095238e-02
R42873 n3_16364_1328 n3_16364_1511 1.161905e-01
R42874 n3_16364_1511 n3_16364_1544 2.095238e-02
R42875 n3_16364_1544 n3_16364_1727 1.161905e-01
R42876 n3_16364_1727 n3_16364_1760 2.095238e-02
R42877 n3_16364_1760 n3_16364_1894 8.507937e-02
R42878 n3_16364_1894 n3_16364_1943 3.111111e-02
R42879 n3_16364_1943 n3_16364_1976 2.095238e-02
R42880 n3_16364_1976 n3_16364_2159 1.161905e-01
R42881 n3_16364_2159 n3_16364_2192 2.095238e-02
R42882 n3_16364_2192 n3_16364_2375 1.161905e-01
R42883 n3_16364_2375 n3_16364_2408 2.095238e-02
R42884 n3_16364_2408 n3_16364_2445 2.349206e-02
R42885 n3_16364_2445 n3_16364_2542 6.158730e-02
R42886 n3_16364_2542 n3_16364_2543 6.349206e-04
R42887 n3_16364_2543 n3_16364_2591 3.047619e-02
R42888 n3_16364_2591 n3_16364_2624 2.095238e-02
R42889 n3_16364_18527 n3_16364_18575 3.047619e-02
R42890 n3_16364_18575 n3_16364_18608 2.095238e-02
R42891 n3_16364_18608 n3_16364_18791 1.161905e-01
R42892 n3_16364_18791 n3_16364_18824 2.095238e-02
R42893 n3_16364_18824 n3_16364_19007 1.161905e-01
R42894 n3_16364_19007 n3_16364_19040 2.095238e-02
R42895 n3_16364_19040 n3_16364_19196 9.904762e-02
R42896 n3_16364_19196 n3_16364_19223 1.714286e-02
R42897 n3_16364_19223 n3_16364_19256 2.095238e-02
R42898 n3_16364_19256 n3_16364_19439 1.161905e-01
R42899 n3_16364_19439 n3_16364_19472 2.095238e-02
R42900 n3_16364_19472 n3_16364_19655 1.161905e-01
R42901 n3_16364_19655 n3_16364_19688 2.095238e-02
R42902 n3_16364_19688 n3_16364_19871 1.161905e-01
R42903 n3_16364_19871 n3_16364_19904 2.095238e-02
R42904 n3_16364_19904 n3_16364_20087 1.161905e-01
R42905 n3_16364_20087 n3_16364_20120 2.095238e-02
R42906 n3_16364_20120 n3_16364_20303 1.161905e-01
R42907 n3_16364_20303 n3_16364_20336 2.095238e-02
R42908 n3_16364_20336 n3_16364_20519 1.161905e-01
R42909 n3_16364_20519 n3_16364_20552 2.095238e-02
R42910 n3_16364_20552 n3_16364_20687 8.571429e-02
R42911 n3_16364_20687 n3_16364_20735 3.047619e-02
R42912 n3_16364_20735 n3_16364_20768 2.095238e-02
R42913 n3_16364_20768 n3_16364_20951 1.161905e-01
R42914 n3_16364_20951 n3_16364_20984 2.095238e-02
R42915 n3_18150_215 n3_18150_248 2.095238e-02
R42916 n3_18150_248 n3_18150_383 8.571429e-02
R42917 n3_18150_383 n3_18150_431 3.047619e-02
R42918 n3_18150_431 n3_18150_464 2.095238e-02
R42919 n3_18150_464 n3_18150_647 1.161905e-01
R42920 n3_18150_647 n3_18150_680 2.095238e-02
R42921 n3_18150_680 n3_18150_863 1.161905e-01
R42922 n3_18150_863 n3_18150_896 2.095238e-02
R42923 n3_18150_896 n3_18150_1079 1.161905e-01
R42924 n3_18150_1079 n3_18150_1112 2.095238e-02
R42925 n3_18150_1112 n3_18150_1295 1.161905e-01
R42926 n3_18150_1295 n3_18150_1328 2.095238e-02
R42927 n3_18150_1328 n3_18150_1511 1.161905e-01
R42928 n3_18150_1511 n3_18150_1544 2.095238e-02
R42929 n3_18150_1544 n3_18150_1727 1.161905e-01
R42930 n3_18150_1727 n3_18150_1760 2.095238e-02
R42931 n3_18150_1760 n3_18150_1894 8.507937e-02
R42932 n3_18150_1894 n3_18150_1943 3.111111e-02
R42933 n3_18150_1943 n3_18150_1976 2.095238e-02
R42934 n3_18150_1976 n3_18150_2159 1.161905e-01
R42935 n3_18150_2159 n3_18150_2192 2.095238e-02
R42936 n3_18150_2192 n3_18150_2375 1.161905e-01
R42937 n3_18150_2375 n3_18150_2408 2.095238e-02
R42938 n3_18150_2408 n3_18150_2542 8.507937e-02
R42939 n3_18150_2542 n3_18150_2543 6.349206e-04
R42940 n3_18150_2543 n3_18150_2591 3.047619e-02
R42941 n3_18150_2591 n3_18150_2624 2.095238e-02
R42942 n3_18150_18527 n3_18150_18575 3.047619e-02
R42943 n3_18150_18575 n3_18150_18608 2.095238e-02
R42944 n3_18150_18608 n3_18150_18791 1.161905e-01
R42945 n3_18150_18791 n3_18150_18824 2.095238e-02
R42946 n3_18150_18824 n3_18150_19007 1.161905e-01
R42947 n3_18150_19007 n3_18150_19040 2.095238e-02
R42948 n3_18150_19040 n3_18150_19223 1.161905e-01
R42949 n3_18150_19223 n3_18150_19256 2.095238e-02
R42950 n3_18150_19256 n3_18150_19439 1.161905e-01
R42951 n3_18150_19439 n3_18150_19472 2.095238e-02
R42952 n3_18150_19472 n3_18150_19655 1.161905e-01
R42953 n3_18150_19655 n3_18150_19688 2.095238e-02
R42954 n3_18150_19688 n3_18150_19871 1.161905e-01
R42955 n3_18150_19871 n3_18150_19904 2.095238e-02
R42956 n3_18150_19904 n3_18150_20087 1.161905e-01
R42957 n3_18150_20087 n3_18150_20120 2.095238e-02
R42958 n3_18150_20120 n3_18150_20303 1.161905e-01
R42959 n3_18150_20303 n3_18150_20336 2.095238e-02
R42960 n3_18150_20336 n3_18150_20519 1.161905e-01
R42961 n3_18150_20519 n3_18150_20552 2.095238e-02
R42962 n3_18150_20552 n3_18150_20687 8.571429e-02
R42963 n3_18150_20687 n3_18150_20735 3.047619e-02
R42964 n3_18150_20735 n3_18150_20768 2.095238e-02
R42965 n3_18150_20768 n3_18150_20951 1.161905e-01
R42966 n3_18150_20951 n3_18150_20984 2.095238e-02
R42967 n3_18333_424 n3_18380_424 2.984127e-02
R42968 n3_18380_424 n3_18521_424 8.952381e-02
R42969 n3_18333_520 n3_18380_520 2.984127e-02
R42970 n3_18380_520 n3_18521_520 8.952381e-02
R42971 n3_18333_2674 n3_18380_2674 2.984127e-02
R42972 n3_18380_2674 n3_18521_2674 8.952381e-02
R42973 n3_18333_2770 n3_18380_2770 2.984127e-02
R42974 n3_18380_2770 n3_18521_2770 8.952381e-02
R42975 n3_18333_4924 n3_18380_4924 2.984127e-02
R42976 n3_18380_4924 n3_18521_4924 8.952381e-02
R42977 n3_18333_5020 n3_18380_5020 2.984127e-02
R42978 n3_18380_5020 n3_18521_5020 8.952381e-02
R42979 n3_18333_7174 n3_18380_7174 2.984127e-02
R42980 n3_18380_7174 n3_18521_7174 8.952381e-02
R42981 n3_18333_7270 n3_18380_7270 2.984127e-02
R42982 n3_18380_7270 n3_18521_7270 8.952381e-02
R42983 n3_18333_9424 n3_18380_9424 2.984127e-02
R42984 n3_18380_9424 n3_18521_9424 8.952381e-02
R42985 n3_18333_9520 n3_18380_9520 2.984127e-02
R42986 n3_18380_9520 n3_18521_9520 8.952381e-02
R42987 n3_18333_11674 n3_18380_11674 2.984127e-02
R42988 n3_18380_11674 n3_18521_11674 8.952381e-02
R42989 n3_18333_11770 n3_18380_11770 2.984127e-02
R42990 n3_18380_11770 n3_18521_11770 8.952381e-02
R42991 n3_18333_13924 n3_18380_13924 2.984127e-02
R42992 n3_18380_13924 n3_18521_13924 8.952381e-02
R42993 n3_18333_14020 n3_18380_14020 2.984127e-02
R42994 n3_18380_14020 n3_18521_14020 8.952381e-02
R42995 n3_18333_16174 n3_18380_16174 2.984127e-02
R42996 n3_18380_16174 n3_18521_16174 8.952381e-02
R42997 n3_18333_16270 n3_18380_16270 2.984127e-02
R42998 n3_18380_16270 n3_18521_16270 8.952381e-02
R42999 n3_18333_18424 n3_18380_18424 2.984127e-02
R43000 n3_18380_18424 n3_18521_18424 8.952381e-02
R43001 n3_18333_18520 n3_18380_18520 2.984127e-02
R43002 n3_18380_18520 n3_18521_18520 8.952381e-02
R43003 n3_18333_20674 n3_18380_20674 2.984127e-02
R43004 n3_18380_20674 n3_18521_20674 8.952381e-02
R43005 n3_18333_20770 n3_18380_20770 2.984127e-02
R43006 n3_18380_20770 n3_18521_20770 8.952381e-02
R43007 n3_18333_215 n3_18333_248 2.095238e-02
R43008 n3_18333_248 n3_18333_383 8.571429e-02
R43009 n3_18333_383 n3_18333_424 2.603175e-02
R43010 n3_18333_424 n3_18333_431 4.444444e-03
R43011 n3_18333_431 n3_18333_464 2.095238e-02
R43012 n3_18333_464 n3_18333_520 3.555556e-02
R43013 n3_18333_520 n3_18333_647 8.063492e-02
R43014 n3_18333_647 n3_18333_680 2.095238e-02
R43015 n3_18333_680 n3_18333_863 1.161905e-01
R43016 n3_18333_863 n3_18333_896 2.095238e-02
R43017 n3_18333_896 n3_18333_1079 1.161905e-01
R43018 n3_18333_1079 n3_18333_1112 2.095238e-02
R43019 n3_18333_1112 n3_18333_1295 1.161905e-01
R43020 n3_18333_1295 n3_18333_1328 2.095238e-02
R43021 n3_18333_1727 n3_18333_1760 2.095238e-02
R43022 n3_18333_1760 n3_18333_1894 8.507937e-02
R43023 n3_18333_1894 n3_18333_1943 3.111111e-02
R43024 n3_18333_1943 n3_18333_1976 2.095238e-02
R43025 n3_18333_1976 n3_18333_2110 8.507937e-02
R43026 n3_18333_2110 n3_18333_2159 3.111111e-02
R43027 n3_18333_2159 n3_18333_2192 2.095238e-02
R43028 n3_18333_2192 n3_18333_2375 1.161905e-01
R43029 n3_18333_2375 n3_18333_2408 2.095238e-02
R43030 n3_18333_2408 n3_18333_2542 8.507937e-02
R43031 n3_18333_2542 n3_18333_2543 6.349206e-04
R43032 n3_18333_2543 n3_18333_2591 3.047619e-02
R43033 n3_18333_2591 n3_18333_2624 2.095238e-02
R43034 n3_18333_2624 n3_18333_2674 3.174603e-02
R43035 n3_18333_2674 n3_18333_2770 6.095238e-02
R43036 n3_18333_2770 n3_18333_2807 2.349206e-02
R43037 n3_18333_2807 n3_18333_2840 2.095238e-02
R43038 n3_18333_2840 n3_18333_3023 1.161905e-01
R43039 n3_18333_3023 n3_18333_3056 2.095238e-02
R43040 n3_18333_3056 n3_18333_3239 1.161905e-01
R43041 n3_18333_3239 n3_18333_3272 2.095238e-02
R43042 n3_18333_3272 n3_18333_3406 8.507937e-02
R43043 n3_18333_3406 n3_18333_3455 3.111111e-02
R43044 n3_18333_3455 n3_18333_3488 2.095238e-02
R43045 n3_18333_3488 n3_18333_3671 1.161905e-01
R43046 n3_18333_3671 n3_18333_3704 2.095238e-02
R43047 n3_18333_4103 n3_18333_4136 2.095238e-02
R43048 n3_18333_4136 n3_18333_4319 1.161905e-01
R43049 n3_18333_4319 n3_18333_4352 2.095238e-02
R43050 n3_18333_4352 n3_18333_4486 8.507937e-02
R43051 n3_18333_4486 n3_18333_4535 3.111111e-02
R43052 n3_18333_4535 n3_18333_4568 2.095238e-02
R43053 n3_18333_4568 n3_18333_4702 8.507937e-02
R43054 n3_18333_4702 n3_18333_4751 3.111111e-02
R43055 n3_18333_4751 n3_18333_4784 2.095238e-02
R43056 n3_18333_4784 n3_18333_4920 8.634921e-02
R43057 n3_18333_4920 n3_18333_4924 2.539683e-03
R43058 n3_18333_4924 n3_18333_4967 2.730159e-02
R43059 n3_18333_4967 n3_18333_5000 2.095238e-02
R43060 n3_18333_5000 n3_18333_5020 1.269841e-02
R43061 n3_18333_5020 n3_18333_5134 7.238095e-02
R43062 n3_18333_5134 n3_18333_5183 3.111111e-02
R43063 n3_18333_5183 n3_18333_5216 2.095238e-02
R43064 n3_18333_5216 n3_18333_5253 2.349206e-02
R43065 n3_18333_5253 n3_18333_5350 6.158730e-02
R43066 n3_18333_5350 n3_18333_5399 3.111111e-02
R43067 n3_18333_5399 n3_18333_5432 2.095238e-02
R43068 n3_18333_5432 n3_18333_5566 8.507937e-02
R43069 n3_18333_5566 n3_18333_5615 3.111111e-02
R43070 n3_18333_5615 n3_18333_5648 2.095238e-02
R43071 n3_18333_5648 n3_18333_5831 1.161905e-01
R43072 n3_18333_5831 n3_18333_5864 2.095238e-02
R43073 n3_18333_6263 n3_18333_6296 2.095238e-02
R43074 n3_18333_6296 n3_18333_6333 2.349206e-02
R43075 n3_18333_6333 n3_18333_6430 6.158730e-02
R43076 n3_18333_6430 n3_18333_6479 3.111111e-02
R43077 n3_18333_6479 n3_18333_6512 2.095238e-02
R43078 n3_18333_6512 n3_18333_6695 1.161905e-01
R43079 n3_18333_6695 n3_18333_6728 2.095238e-02
R43080 n3_18333_6728 n3_18333_6911 1.161905e-01
R43081 n3_18333_6911 n3_18333_6944 2.095238e-02
R43082 n3_18333_6944 n3_18333_7127 1.161905e-01
R43083 n3_18333_7127 n3_18333_7160 2.095238e-02
R43084 n3_18333_7160 n3_18333_7174 8.888889e-03
R43085 n3_18333_7174 n3_18333_7270 6.095238e-02
R43086 n3_18333_7270 n3_18333_7343 4.634921e-02
R43087 n3_18333_7343 n3_18333_7376 2.095238e-02
R43088 n3_18333_7376 n3_18333_7559 1.161905e-01
R43089 n3_18333_7559 n3_18333_7592 2.095238e-02
R43090 n3_18333_7592 n3_18333_7775 1.161905e-01
R43091 n3_18333_7775 n3_18333_7808 2.095238e-02
R43092 n3_18333_7808 n3_18333_7845 2.349206e-02
R43093 n3_18333_7845 n3_18333_7942 6.158730e-02
R43094 n3_18333_7942 n3_18333_7991 3.111111e-02
R43095 n3_18333_7991 n3_18333_8024 2.095238e-02
R43096 n3_18333_8024 n3_18333_8207 1.161905e-01
R43097 n3_18333_8207 n3_18333_8240 2.095238e-02
R43098 n3_18333_8456 n3_18333_8639 1.161905e-01
R43099 n3_18333_8639 n3_18333_8672 2.095238e-02
R43100 n3_18333_8672 n3_18333_8855 1.161905e-01
R43101 n3_18333_8855 n3_18333_8888 2.095238e-02
R43102 n3_18333_8888 n3_18333_8925 2.349206e-02
R43103 n3_18333_8925 n3_18333_9022 6.158730e-02
R43104 n3_18333_9022 n3_18333_9071 3.111111e-02
R43105 n3_18333_9071 n3_18333_9104 2.095238e-02
R43106 n3_18333_9104 n3_18333_9287 1.161905e-01
R43107 n3_18333_9287 n3_18333_9320 2.095238e-02
R43108 n3_18333_9320 n3_18333_9424 6.603175e-02
R43109 n3_18333_9424 n3_18333_9503 5.015873e-02
R43110 n3_18333_9503 n3_18333_9520 1.079365e-02
R43111 n3_18333_9520 n3_18333_9536 1.015873e-02
R43112 n3_18333_9536 n3_18333_9719 1.161905e-01
R43113 n3_18333_9719 n3_18333_9752 2.095238e-02
R43114 n3_18333_9752 n3_18333_9935 1.161905e-01
R43115 n3_18333_9935 n3_18333_9968 2.095238e-02
R43116 n3_18333_9968 n3_18333_10005 2.349206e-02
R43117 n3_18333_10005 n3_18333_10102 6.158730e-02
R43118 n3_18333_10102 n3_18333_10151 3.111111e-02
R43119 n3_18333_10151 n3_18333_10184 2.095238e-02
R43120 n3_18333_10184 n3_18333_10367 1.161905e-01
R43121 n3_18333_10367 n3_18333_10400 2.095238e-02
R43122 n3_18333_10799 n3_18333_10832 2.095238e-02
R43123 n3_18333_10832 n3_18333_11015 1.161905e-01
R43124 n3_18333_11015 n3_18333_11048 2.095238e-02
R43125 n3_18333_11048 n3_18333_11196 9.396825e-02
R43126 n3_18333_11196 n3_18333_11231 2.222222e-02
R43127 n3_18333_11231 n3_18333_11264 2.095238e-02
R43128 n3_18333_11264 n3_18333_11447 1.161905e-01
R43129 n3_18333_11447 n3_18333_11480 2.095238e-02
R43130 n3_18333_11480 n3_18333_11663 1.161905e-01
R43131 n3_18333_11663 n3_18333_11674 6.984127e-03
R43132 n3_18333_11674 n3_18333_11696 1.396825e-02
R43133 n3_18333_11696 n3_18333_11770 4.698413e-02
R43134 n3_18333_11770 n3_18333_11879 6.920635e-02
R43135 n3_18333_11879 n3_18333_11912 2.095238e-02
R43136 n3_18333_11912 n3_18333_12095 1.161905e-01
R43137 n3_18333_12095 n3_18333_12128 2.095238e-02
R43138 n3_18333_12128 n3_18333_12284 9.904762e-02
R43139 n3_18333_12284 n3_18333_12311 1.714286e-02
R43140 n3_18333_12311 n3_18333_12344 2.095238e-02
R43141 n3_18333_12344 n3_18333_12527 1.161905e-01
R43142 n3_18333_12527 n3_18333_12560 2.095238e-02
R43143 n3_18333_12560 n3_18333_12743 1.161905e-01
R43144 n3_18333_12959 n3_18333_12992 2.095238e-02
R43145 n3_18333_12992 n3_18333_13175 1.161905e-01
R43146 n3_18333_13175 n3_18333_13208 2.095238e-02
R43147 n3_18333_13208 n3_18333_13391 1.161905e-01
R43148 n3_18333_13391 n3_18333_13424 2.095238e-02
R43149 n3_18333_13424 n3_18333_13607 1.161905e-01
R43150 n3_18333_13607 n3_18333_13640 2.095238e-02
R43151 n3_18333_13640 n3_18333_13788 9.396825e-02
R43152 n3_18333_13788 n3_18333_13796 5.079365e-03
R43153 n3_18333_13796 n3_18333_13823 1.714286e-02
R43154 n3_18333_13823 n3_18333_13856 2.095238e-02
R43155 n3_18333_13856 n3_18333_13924 4.317460e-02
R43156 n3_18333_13924 n3_18333_14020 6.095238e-02
R43157 n3_18333_14020 n3_18333_14039 1.206349e-02
R43158 n3_18333_14039 n3_18333_14072 2.095238e-02
R43159 n3_18333_14072 n3_18333_14255 1.161905e-01
R43160 n3_18333_14255 n3_18333_14288 2.095238e-02
R43161 n3_18333_14288 n3_18333_14471 1.161905e-01
R43162 n3_18333_14471 n3_18333_14504 2.095238e-02
R43163 n3_18333_14504 n3_18333_14652 9.396825e-02
R43164 n3_18333_14652 n3_18333_14660 5.079365e-03
R43165 n3_18333_14660 n3_18333_14687 1.714286e-02
R43166 n3_18333_14687 n3_18333_14720 2.095238e-02
R43167 n3_18333_14720 n3_18333_14903 1.161905e-01
R43168 n3_18333_14903 n3_18333_14936 2.095238e-02
R43169 n3_18333_15308 n3_18333_15335 1.714286e-02
R43170 n3_18333_15335 n3_18333_15368 2.095238e-02
R43171 n3_18333_15368 n3_18333_15551 1.161905e-01
R43172 n3_18333_15551 n3_18333_15584 2.095238e-02
R43173 n3_18333_15584 n3_18333_15740 9.904762e-02
R43174 n3_18333_15740 n3_18333_15767 1.714286e-02
R43175 n3_18333_15767 n3_18333_15800 2.095238e-02
R43176 n3_18333_15800 n3_18333_15983 1.161905e-01
R43177 n3_18333_15983 n3_18333_16016 2.095238e-02
R43178 n3_18333_16016 n3_18333_16174 1.003175e-01
R43179 n3_18333_16174 n3_18333_16199 1.587302e-02
R43180 n3_18333_16199 n3_18333_16232 2.095238e-02
R43181 n3_18333_16232 n3_18333_16270 2.412698e-02
R43182 n3_18333_16270 n3_18333_16415 9.206349e-02
R43183 n3_18333_16415 n3_18333_16448 2.095238e-02
R43184 n3_18333_16448 n3_18333_16631 1.161905e-01
R43185 n3_18333_16631 n3_18333_16664 2.095238e-02
R43186 n3_18333_16664 n3_18333_16812 9.396825e-02
R43187 n3_18333_16812 n3_18333_16820 5.079365e-03
R43188 n3_18333_16820 n3_18333_16847 1.714286e-02
R43189 n3_18333_16847 n3_18333_16880 2.095238e-02
R43190 n3_18333_16880 n3_18333_17063 1.161905e-01
R43191 n3_18333_17063 n3_18333_17096 2.095238e-02
R43192 n3_18333_17096 n3_18333_17230 8.507937e-02
R43193 n3_18333_17495 n3_18333_17528 2.095238e-02
R43194 n3_18333_17528 n3_18333_17711 1.161905e-01
R43195 n3_18333_17711 n3_18333_17744 2.095238e-02
R43196 n3_18333_17744 n3_18333_17900 9.904762e-02
R43197 n3_18333_17900 n3_18333_17927 1.714286e-02
R43198 n3_18333_17927 n3_18333_17960 2.095238e-02
R43199 n3_18333_17960 n3_18333_18143 1.161905e-01
R43200 n3_18333_18143 n3_18333_18176 2.095238e-02
R43201 n3_18333_18176 n3_18333_18359 1.161905e-01
R43202 n3_18333_18359 n3_18333_18392 2.095238e-02
R43203 n3_18333_18392 n3_18333_18424 2.031746e-02
R43204 n3_18333_18424 n3_18333_18520 6.095238e-02
R43205 n3_18333_18520 n3_18333_18527 4.444444e-03
R43206 n3_18333_18527 n3_18333_18575 3.047619e-02
R43207 n3_18333_18575 n3_18333_18608 2.095238e-02
R43208 n3_18333_18608 n3_18333_18791 1.161905e-01
R43209 n3_18333_18791 n3_18333_18824 2.095238e-02
R43210 n3_18333_18824 n3_18333_19007 1.161905e-01
R43211 n3_18333_19007 n3_18333_19040 2.095238e-02
R43212 n3_18333_19040 n3_18333_19223 1.161905e-01
R43213 n3_18333_19223 n3_18333_19256 2.095238e-02
R43214 n3_18333_19256 n3_18333_19439 1.161905e-01
R43215 n3_18333_19439 n3_18333_19472 2.095238e-02
R43216 n3_18333_19871 n3_18333_19904 2.095238e-02
R43217 n3_18333_19904 n3_18333_20087 1.161905e-01
R43218 n3_18333_20087 n3_18333_20120 2.095238e-02
R43219 n3_18333_20120 n3_18333_20303 1.161905e-01
R43220 n3_18333_20303 n3_18333_20336 2.095238e-02
R43221 n3_18333_20336 n3_18333_20519 1.161905e-01
R43222 n3_18333_20519 n3_18333_20552 2.095238e-02
R43223 n3_18333_20552 n3_18333_20674 7.746032e-02
R43224 n3_18333_20674 n3_18333_20687 8.253968e-03
R43225 n3_18333_20687 n3_18333_20735 3.047619e-02
R43226 n3_18333_20735 n3_18333_20768 2.095238e-02
R43227 n3_18333_20768 n3_18333_20770 1.269841e-03
R43228 n3_18333_20770 n3_18333_20951 1.149206e-01
R43229 n3_18333_20951 n3_18333_20984 2.095238e-02
R43230 n3_18521_215 n3_18521_248 2.095238e-02
R43231 n3_18521_248 n3_18521_383 8.571429e-02
R43232 n3_18521_383 n3_18521_424 2.603175e-02
R43233 n3_18521_424 n3_18521_431 4.444444e-03
R43234 n3_18521_520 n3_18521_647 8.063492e-02
R43235 n3_18521_647 n3_18521_680 2.095238e-02
R43236 n3_18521_680 n3_18521_863 1.161905e-01
R43237 n3_18521_863 n3_18521_896 2.095238e-02
R43238 n3_18521_896 n3_18521_1079 1.161905e-01
R43239 n3_18521_1079 n3_18521_1112 2.095238e-02
R43240 n3_18521_1112 n3_18521_1295 1.161905e-01
R43241 n3_18521_1295 n3_18521_1328 2.095238e-02
R43242 n3_18521_1328 n3_18521_1511 1.161905e-01
R43243 n3_18521_1511 n3_18521_1544 2.095238e-02
R43244 n3_18521_1544 n3_18521_1727 1.161905e-01
R43245 n3_18521_1727 n3_18521_1760 2.095238e-02
R43246 n3_18521_1760 n3_18521_1894 8.507937e-02
R43247 n3_18521_1894 n3_18521_1943 3.111111e-02
R43248 n3_18521_1943 n3_18521_1976 2.095238e-02
R43249 n3_18521_1976 n3_18521_2110 8.507937e-02
R43250 n3_18521_2110 n3_18521_2159 3.111111e-02
R43251 n3_18521_2159 n3_18521_2192 2.095238e-02
R43252 n3_18521_2192 n3_18521_2375 1.161905e-01
R43253 n3_18521_2375 n3_18521_2408 2.095238e-02
R43254 n3_18521_2408 n3_18521_2542 8.507937e-02
R43255 n3_18521_2542 n3_18521_2543 6.349206e-04
R43256 n3_18521_2543 n3_18521_2591 3.047619e-02
R43257 n3_18521_2591 n3_18521_2624 2.095238e-02
R43258 n3_18521_2624 n3_18521_2674 3.174603e-02
R43259 n3_18521_2770 n3_18521_2807 2.349206e-02
R43260 n3_18521_2807 n3_18521_2840 2.095238e-02
R43261 n3_18521_2840 n3_18521_3023 1.161905e-01
R43262 n3_18521_3023 n3_18521_3056 2.095238e-02
R43263 n3_18521_3056 n3_18521_3239 1.161905e-01
R43264 n3_18521_3239 n3_18521_3272 2.095238e-02
R43265 n3_18521_3272 n3_18521_3406 8.507937e-02
R43266 n3_18521_3406 n3_18521_3455 3.111111e-02
R43267 n3_18521_3455 n3_18521_3488 2.095238e-02
R43268 n3_18521_3488 n3_18521_3671 1.161905e-01
R43269 n3_18521_3671 n3_18521_3704 2.095238e-02
R43270 n3_18521_3704 n3_18521_3887 1.161905e-01
R43271 n3_18521_3887 n3_18521_3920 2.095238e-02
R43272 n3_18521_3920 n3_18521_4103 1.161905e-01
R43273 n3_18521_4103 n3_18521_4136 2.095238e-02
R43274 n3_18521_4136 n3_18521_4319 1.161905e-01
R43275 n3_18521_4319 n3_18521_4352 2.095238e-02
R43276 n3_18521_4352 n3_18521_4486 8.507937e-02
R43277 n3_18521_4486 n3_18521_4535 3.111111e-02
R43278 n3_18521_4535 n3_18521_4568 2.095238e-02
R43279 n3_18521_4568 n3_18521_4702 8.507937e-02
R43280 n3_18521_4702 n3_18521_4751 3.111111e-02
R43281 n3_18521_4751 n3_18521_4784 2.095238e-02
R43282 n3_18521_4784 n3_18521_4920 8.634921e-02
R43283 n3_18521_4920 n3_18521_4924 2.539683e-03
R43284 n3_18521_5000 n3_18521_5020 1.269841e-02
R43285 n3_18521_5020 n3_18521_5134 7.238095e-02
R43286 n3_18521_5134 n3_18521_5183 3.111111e-02
R43287 n3_18521_5183 n3_18521_5216 2.095238e-02
R43288 n3_18521_5216 n3_18521_5253 2.349206e-02
R43289 n3_18521_5253 n3_18521_5350 6.158730e-02
R43290 n3_18521_5350 n3_18521_5399 3.111111e-02
R43291 n3_18521_5399 n3_18521_5432 2.095238e-02
R43292 n3_18521_5432 n3_18521_5566 8.507937e-02
R43293 n3_18521_5566 n3_18521_5615 3.111111e-02
R43294 n3_18521_5615 n3_18521_5648 2.095238e-02
R43295 n3_18521_5648 n3_18521_5831 1.161905e-01
R43296 n3_18521_5831 n3_18521_5864 2.095238e-02
R43297 n3_18521_5864 n3_18521_6047 1.161905e-01
R43298 n3_18521_6047 n3_18521_6080 2.095238e-02
R43299 n3_18521_6080 n3_18521_6263 1.161905e-01
R43300 n3_18521_6263 n3_18521_6296 2.095238e-02
R43301 n3_18521_6296 n3_18521_6333 2.349206e-02
R43302 n3_18521_6333 n3_18521_6430 6.158730e-02
R43303 n3_18521_6430 n3_18521_6479 3.111111e-02
R43304 n3_18521_6479 n3_18521_6512 2.095238e-02
R43305 n3_18521_6512 n3_18521_6695 1.161905e-01
R43306 n3_18521_6695 n3_18521_6728 2.095238e-02
R43307 n3_18521_6728 n3_18521_6911 1.161905e-01
R43308 n3_18521_6911 n3_18521_6944 2.095238e-02
R43309 n3_18521_6944 n3_18521_7127 1.161905e-01
R43310 n3_18521_7127 n3_18521_7160 2.095238e-02
R43311 n3_18521_7160 n3_18521_7174 8.888889e-03
R43312 n3_18521_7270 n3_18521_7343 4.634921e-02
R43313 n3_18521_7343 n3_18521_7376 2.095238e-02
R43314 n3_18521_7376 n3_18521_7559 1.161905e-01
R43315 n3_18521_7559 n3_18521_7592 2.095238e-02
R43316 n3_18521_7592 n3_18521_7775 1.161905e-01
R43317 n3_18521_7775 n3_18521_7808 2.095238e-02
R43318 n3_18521_7808 n3_18521_7845 2.349206e-02
R43319 n3_18521_7845 n3_18521_7942 6.158730e-02
R43320 n3_18521_7942 n3_18521_7991 3.111111e-02
R43321 n3_18521_7991 n3_18521_8024 2.095238e-02
R43322 n3_18521_8024 n3_18521_8207 1.161905e-01
R43323 n3_18521_8207 n3_18521_8240 2.095238e-02
R43324 n3_18521_8240 n3_18521_8423 1.161905e-01
R43325 n3_18521_8423 n3_18521_8456 2.095238e-02
R43326 n3_18521_8456 n3_18521_8639 1.161905e-01
R43327 n3_18521_8639 n3_18521_8672 2.095238e-02
R43328 n3_18521_8672 n3_18521_8855 1.161905e-01
R43329 n3_18521_8855 n3_18521_8888 2.095238e-02
R43330 n3_18521_8888 n3_18521_8925 2.349206e-02
R43331 n3_18521_8925 n3_18521_9022 6.158730e-02
R43332 n3_18521_9022 n3_18521_9071 3.111111e-02
R43333 n3_18521_9071 n3_18521_9104 2.095238e-02
R43334 n3_18521_9104 n3_18521_9287 1.161905e-01
R43335 n3_18521_9287 n3_18521_9320 2.095238e-02
R43336 n3_18521_9320 n3_18521_9424 6.603175e-02
R43337 n3_18521_9503 n3_18521_9520 1.079365e-02
R43338 n3_18521_9520 n3_18521_9536 1.015873e-02
R43339 n3_18521_9536 n3_18521_9719 1.161905e-01
R43340 n3_18521_9719 n3_18521_9752 2.095238e-02
R43341 n3_18521_9752 n3_18521_9935 1.161905e-01
R43342 n3_18521_9935 n3_18521_9968 2.095238e-02
R43343 n3_18521_9968 n3_18521_10005 2.349206e-02
R43344 n3_18521_10005 n3_18521_10102 6.158730e-02
R43345 n3_18521_10102 n3_18521_10151 3.111111e-02
R43346 n3_18521_10151 n3_18521_10184 2.095238e-02
R43347 n3_18521_10184 n3_18521_10367 1.161905e-01
R43348 n3_18521_10367 n3_18521_10400 2.095238e-02
R43349 n3_18521_10616 n3_18521_10799 1.161905e-01
R43350 n3_18521_10799 n3_18521_10832 2.095238e-02
R43351 n3_18521_10832 n3_18521_11015 1.161905e-01
R43352 n3_18521_11015 n3_18521_11048 2.095238e-02
R43353 n3_18521_11048 n3_18521_11196 9.396825e-02
R43354 n3_18521_11196 n3_18521_11231 2.222222e-02
R43355 n3_18521_11231 n3_18521_11264 2.095238e-02
R43356 n3_18521_11264 n3_18521_11447 1.161905e-01
R43357 n3_18521_11447 n3_18521_11480 2.095238e-02
R43358 n3_18521_11480 n3_18521_11663 1.161905e-01
R43359 n3_18521_11663 n3_18521_11674 6.984127e-03
R43360 n3_18521_11674 n3_18521_11696 1.396825e-02
R43361 n3_18521_11770 n3_18521_11879 6.920635e-02
R43362 n3_18521_11879 n3_18521_11912 2.095238e-02
R43363 n3_18521_11912 n3_18521_12095 1.161905e-01
R43364 n3_18521_12095 n3_18521_12128 2.095238e-02
R43365 n3_18521_12128 n3_18521_12284 9.904762e-02
R43366 n3_18521_12284 n3_18521_12311 1.714286e-02
R43367 n3_18521_12311 n3_18521_12344 2.095238e-02
R43368 n3_18521_12344 n3_18521_12527 1.161905e-01
R43369 n3_18521_12527 n3_18521_12560 2.095238e-02
R43370 n3_18521_12560 n3_18521_12743 1.161905e-01
R43371 n3_18521_12743 n3_18521_12776 2.095238e-02
R43372 n3_18521_12776 n3_18521_12959 1.161905e-01
R43373 n3_18521_12959 n3_18521_12992 2.095238e-02
R43374 n3_18521_12992 n3_18521_13175 1.161905e-01
R43375 n3_18521_13175 n3_18521_13208 2.095238e-02
R43376 n3_18521_13208 n3_18521_13391 1.161905e-01
R43377 n3_18521_13391 n3_18521_13424 2.095238e-02
R43378 n3_18521_13424 n3_18521_13607 1.161905e-01
R43379 n3_18521_13607 n3_18521_13640 2.095238e-02
R43380 n3_18521_13640 n3_18521_13788 9.396825e-02
R43381 n3_18521_13788 n3_18521_13796 5.079365e-03
R43382 n3_18521_13796 n3_18521_13823 1.714286e-02
R43383 n3_18521_13823 n3_18521_13856 2.095238e-02
R43384 n3_18521_13856 n3_18521_13924 4.317460e-02
R43385 n3_18521_14020 n3_18521_14039 1.206349e-02
R43386 n3_18521_14039 n3_18521_14072 2.095238e-02
R43387 n3_18521_14072 n3_18521_14255 1.161905e-01
R43388 n3_18521_14255 n3_18521_14288 2.095238e-02
R43389 n3_18521_14288 n3_18521_14471 1.161905e-01
R43390 n3_18521_14471 n3_18521_14504 2.095238e-02
R43391 n3_18521_14504 n3_18521_14652 9.396825e-02
R43392 n3_18521_14652 n3_18521_14660 5.079365e-03
R43393 n3_18521_14660 n3_18521_14687 1.714286e-02
R43394 n3_18521_14687 n3_18521_14720 2.095238e-02
R43395 n3_18521_14720 n3_18521_14903 1.161905e-01
R43396 n3_18521_14903 n3_18521_14936 2.095238e-02
R43397 n3_18521_14936 n3_18521_15092 9.904762e-02
R43398 n3_18521_15092 n3_18521_15119 1.714286e-02
R43399 n3_18521_15119 n3_18521_15152 2.095238e-02
R43400 n3_18521_15152 n3_18521_15308 9.904762e-02
R43401 n3_18521_15308 n3_18521_15335 1.714286e-02
R43402 n3_18521_15335 n3_18521_15368 2.095238e-02
R43403 n3_18521_15368 n3_18521_15551 1.161905e-01
R43404 n3_18521_15551 n3_18521_15584 2.095238e-02
R43405 n3_18521_15584 n3_18521_15740 9.904762e-02
R43406 n3_18521_15740 n3_18521_15767 1.714286e-02
R43407 n3_18521_15767 n3_18521_15800 2.095238e-02
R43408 n3_18521_15800 n3_18521_15983 1.161905e-01
R43409 n3_18521_15983 n3_18521_16016 2.095238e-02
R43410 n3_18521_16016 n3_18521_16174 1.003175e-01
R43411 n3_18521_16174 n3_18521_16199 1.587302e-02
R43412 n3_18521_16270 n3_18521_16415 9.206349e-02
R43413 n3_18521_16415 n3_18521_16448 2.095238e-02
R43414 n3_18521_16448 n3_18521_16631 1.161905e-01
R43415 n3_18521_16631 n3_18521_16664 2.095238e-02
R43416 n3_18521_16664 n3_18521_16812 9.396825e-02
R43417 n3_18521_16812 n3_18521_16820 5.079365e-03
R43418 n3_18521_16820 n3_18521_16847 1.714286e-02
R43419 n3_18521_16847 n3_18521_16880 2.095238e-02
R43420 n3_18521_16880 n3_18521_17063 1.161905e-01
R43421 n3_18521_17063 n3_18521_17096 2.095238e-02
R43422 n3_18521_17096 n3_18521_17230 8.507937e-02
R43423 n3_18521_17230 n3_18521_17279 3.111111e-02
R43424 n3_18521_17279 n3_18521_17312 2.095238e-02
R43425 n3_18521_17312 n3_18521_17495 1.161905e-01
R43426 n3_18521_17495 n3_18521_17528 2.095238e-02
R43427 n3_18521_17528 n3_18521_17711 1.161905e-01
R43428 n3_18521_17711 n3_18521_17744 2.095238e-02
R43429 n3_18521_17744 n3_18521_17900 9.904762e-02
R43430 n3_18521_17900 n3_18521_17927 1.714286e-02
R43431 n3_18521_17927 n3_18521_17960 2.095238e-02
R43432 n3_18521_17960 n3_18521_18143 1.161905e-01
R43433 n3_18521_18143 n3_18521_18176 2.095238e-02
R43434 n3_18521_18176 n3_18521_18359 1.161905e-01
R43435 n3_18521_18359 n3_18521_18392 2.095238e-02
R43436 n3_18521_18392 n3_18521_18424 2.031746e-02
R43437 n3_18521_18520 n3_18521_18527 4.444444e-03
R43438 n3_18521_18527 n3_18521_18575 3.047619e-02
R43439 n3_18521_18575 n3_18521_18608 2.095238e-02
R43440 n3_18521_18608 n3_18521_18791 1.161905e-01
R43441 n3_18521_18791 n3_18521_18824 2.095238e-02
R43442 n3_18521_18824 n3_18521_19007 1.161905e-01
R43443 n3_18521_19007 n3_18521_19040 2.095238e-02
R43444 n3_18521_19040 n3_18521_19223 1.161905e-01
R43445 n3_18521_19223 n3_18521_19256 2.095238e-02
R43446 n3_18521_19256 n3_18521_19439 1.161905e-01
R43447 n3_18521_19439 n3_18521_19472 2.095238e-02
R43448 n3_18521_19472 n3_18521_19655 1.161905e-01
R43449 n3_18521_19655 n3_18521_19688 2.095238e-02
R43450 n3_18521_19688 n3_18521_19871 1.161905e-01
R43451 n3_18521_19871 n3_18521_19904 2.095238e-02
R43452 n3_18521_19904 n3_18521_20087 1.161905e-01
R43453 n3_18521_20087 n3_18521_20120 2.095238e-02
R43454 n3_18521_20120 n3_18521_20303 1.161905e-01
R43455 n3_18521_20303 n3_18521_20336 2.095238e-02
R43456 n3_18521_20336 n3_18521_20519 1.161905e-01
R43457 n3_18521_20519 n3_18521_20552 2.095238e-02
R43458 n3_18521_20552 n3_18521_20674 7.746032e-02
R43459 n3_18521_20674 n3_18521_20687 8.253968e-03
R43460 n3_18521_20768 n3_18521_20770 1.269841e-03
R43461 n3_18521_20770 n3_18521_20951 1.149206e-01
R43462 n3_18521_20951 n3_18521_20984 2.095238e-02
R43463 n3_18614_215 n3_18614_248 2.095238e-02
R43464 n3_18614_248 n3_18614_383 8.571429e-02
R43465 n3_18614_383 n3_18614_431 3.047619e-02
R43466 n3_18614_431 n3_18614_464 2.095238e-02
R43467 n3_18614_464 n3_18614_647 1.161905e-01
R43468 n3_18614_647 n3_18614_680 2.095238e-02
R43469 n3_18614_680 n3_18614_863 1.161905e-01
R43470 n3_18614_863 n3_18614_896 2.095238e-02
R43471 n3_18614_896 n3_18614_1079 1.161905e-01
R43472 n3_18614_1079 n3_18614_1112 2.095238e-02
R43473 n3_18614_1112 n3_18614_1295 1.161905e-01
R43474 n3_18614_1295 n3_18614_1328 2.095238e-02
R43475 n3_18614_1328 n3_18614_1511 1.161905e-01
R43476 n3_18614_1511 n3_18614_1544 2.095238e-02
R43477 n3_18614_1544 n3_18614_1727 1.161905e-01
R43478 n3_18614_1727 n3_18614_1760 2.095238e-02
R43479 n3_18614_1760 n3_18614_1943 1.161905e-01
R43480 n3_18614_1943 n3_18614_1976 2.095238e-02
R43481 n3_18614_1976 n3_18614_2110 8.507937e-02
R43482 n3_18614_2110 n3_18614_2159 3.111111e-02
R43483 n3_18614_2159 n3_18614_2192 2.095238e-02
R43484 n3_18614_2192 n3_18614_2375 1.161905e-01
R43485 n3_18614_2375 n3_18614_2408 2.095238e-02
R43486 n3_18614_2408 n3_18614_2543 8.571429e-02
R43487 n3_18614_2543 n3_18614_2591 3.047619e-02
R43488 n3_18614_2591 n3_18614_2624 2.095238e-02
R43489 n3_18614_18527 n3_18614_18575 3.047619e-02
R43490 n3_18614_18575 n3_18614_18608 2.095238e-02
R43491 n3_18614_18608 n3_18614_18791 1.161905e-01
R43492 n3_18614_18791 n3_18614_18824 2.095238e-02
R43493 n3_18614_18824 n3_18614_19007 1.161905e-01
R43494 n3_18614_19007 n3_18614_19040 2.095238e-02
R43495 n3_18614_19040 n3_18614_19223 1.161905e-01
R43496 n3_18614_19223 n3_18614_19256 2.095238e-02
R43497 n3_18614_19256 n3_18614_19439 1.161905e-01
R43498 n3_18614_19439 n3_18614_19472 2.095238e-02
R43499 n3_18614_19472 n3_18614_19655 1.161905e-01
R43500 n3_18614_19655 n3_18614_19688 2.095238e-02
R43501 n3_18614_19688 n3_18614_19871 1.161905e-01
R43502 n3_18614_19871 n3_18614_19904 2.095238e-02
R43503 n3_18614_19904 n3_18614_20087 1.161905e-01
R43504 n3_18614_20087 n3_18614_20120 2.095238e-02
R43505 n3_18614_20120 n3_18614_20303 1.161905e-01
R43506 n3_18614_20303 n3_18614_20336 2.095238e-02
R43507 n3_18614_20336 n3_18614_20519 1.161905e-01
R43508 n3_18614_20519 n3_18614_20552 2.095238e-02
R43509 n3_18614_20552 n3_18614_20687 8.571429e-02
R43510 n3_18614_20687 n3_18614_20735 3.047619e-02
R43511 n3_18614_20735 n3_18614_20768 2.095238e-02
R43512 n3_18614_20768 n3_18614_20951 1.161905e-01
R43513 n3_18614_20951 n3_18614_20984 2.095238e-02
R43514 n3_20583_424 n3_20630_424 2.984127e-02
R43515 n3_20583_520 n3_20630_520 2.984127e-02
R43516 n3_20630_520 n3_20771_520 8.952381e-02
R43517 n3_20583_2674 n3_20630_2674 2.984127e-02
R43518 n3_20630_2674 n3_20771_2674 8.952381e-02
R43519 n3_20583_2770 n3_20630_2770 2.984127e-02
R43520 n3_20630_2770 n3_20771_2770 8.952381e-02
R43521 n3_20583_4924 n3_20630_4924 2.984127e-02
R43522 n3_20630_4924 n3_20771_4924 8.952381e-02
R43523 n3_20583_5020 n3_20630_5020 2.984127e-02
R43524 n3_20630_5020 n3_20771_5020 8.952381e-02
R43525 n3_20583_7174 n3_20630_7174 2.984127e-02
R43526 n3_20630_7174 n3_20771_7174 8.952381e-02
R43527 n3_20583_7270 n3_20630_7270 2.984127e-02
R43528 n3_20630_7270 n3_20771_7270 8.952381e-02
R43529 n3_20583_9424 n3_20630_9424 2.984127e-02
R43530 n3_20630_9424 n3_20771_9424 8.952381e-02
R43531 n3_20583_9520 n3_20630_9520 2.984127e-02
R43532 n3_20630_9520 n3_20771_9520 8.952381e-02
R43533 n3_20583_11674 n3_20630_11674 2.984127e-02
R43534 n3_20630_11674 n3_20771_11674 8.952381e-02
R43535 n3_20583_11770 n3_20630_11770 2.984127e-02
R43536 n3_20630_11770 n3_20771_11770 8.952381e-02
R43537 n3_20583_13924 n3_20630_13924 2.984127e-02
R43538 n3_20630_13924 n3_20771_13924 8.952381e-02
R43539 n3_20583_14020 n3_20630_14020 2.984127e-02
R43540 n3_20630_14020 n3_20771_14020 8.952381e-02
R43541 n3_20583_16174 n3_20630_16174 2.984127e-02
R43542 n3_20630_16174 n3_20771_16174 8.952381e-02
R43543 n3_20583_16270 n3_20630_16270 2.984127e-02
R43544 n3_20630_16270 n3_20771_16270 8.952381e-02
R43545 n3_20583_18424 n3_20630_18424 2.984127e-02
R43546 n3_20630_18424 n3_20771_18424 8.952381e-02
R43547 n3_20583_18520 n3_20630_18520 2.984127e-02
R43548 n3_20630_18520 n3_20771_18520 8.952381e-02
R43549 n3_20583_20674 n3_20630_20674 2.984127e-02
R43550 n3_20630_20674 n3_20771_20674 8.952381e-02
R43551 n3_20583_20770 n3_20630_20770 2.984127e-02
R43552 n3_20583_215 n3_20583_248 2.095238e-02
R43553 n3_20583_248 n3_20583_383 8.571429e-02
R43554 n3_20583_383 n3_20583_424 2.603175e-02
R43555 n3_20583_424 n3_20583_431 4.444444e-03
R43556 n3_20583_431 n3_20583_464 2.095238e-02
R43557 n3_20583_464 n3_20583_520 3.555556e-02
R43558 n3_20583_520 n3_20583_647 8.063492e-02
R43559 n3_20583_647 n3_20583_680 2.095238e-02
R43560 n3_20583_680 n3_20583_863 1.161905e-01
R43561 n3_20583_863 n3_20583_896 2.095238e-02
R43562 n3_20583_896 n3_20583_1079 1.161905e-01
R43563 n3_20583_1079 n3_20583_1112 2.095238e-02
R43564 n3_20583_1112 n3_20583_1295 1.161905e-01
R43565 n3_20583_1295 n3_20583_1328 2.095238e-02
R43566 n3_20583_1727 n3_20583_1760 2.095238e-02
R43567 n3_20583_1760 n3_20583_1943 1.161905e-01
R43568 n3_20583_1943 n3_20583_1976 2.095238e-02
R43569 n3_20583_1976 n3_20583_2159 1.161905e-01
R43570 n3_20583_2159 n3_20583_2192 2.095238e-02
R43571 n3_20583_2192 n3_20583_2375 1.161905e-01
R43572 n3_20583_2375 n3_20583_2408 2.095238e-02
R43573 n3_20583_2408 n3_20583_2543 8.571429e-02
R43574 n3_20583_2543 n3_20583_2591 3.047619e-02
R43575 n3_20583_2591 n3_20583_2624 2.095238e-02
R43576 n3_20583_2624 n3_20583_2674 3.174603e-02
R43577 n3_20583_2674 n3_20583_2770 6.095238e-02
R43578 n3_20583_2770 n3_20583_2807 2.349206e-02
R43579 n3_20583_2807 n3_20583_2840 2.095238e-02
R43580 n3_20583_2840 n3_20583_3023 1.161905e-01
R43581 n3_20583_3023 n3_20583_3056 2.095238e-02
R43582 n3_20583_3056 n3_20583_3239 1.161905e-01
R43583 n3_20583_3239 n3_20583_3272 2.095238e-02
R43584 n3_20583_3272 n3_20583_3455 1.161905e-01
R43585 n3_20583_3455 n3_20583_3488 2.095238e-02
R43586 n3_20583_3488 n3_20583_3671 1.161905e-01
R43587 n3_20583_3671 n3_20583_3704 2.095238e-02
R43588 n3_20583_4103 n3_20583_4136 2.095238e-02
R43589 n3_20583_4136 n3_20583_4319 1.161905e-01
R43590 n3_20583_4319 n3_20583_4352 2.095238e-02
R43591 n3_20583_4352 n3_20583_4535 1.161905e-01
R43592 n3_20583_4535 n3_20583_4568 2.095238e-02
R43593 n3_20583_4568 n3_20583_4751 1.161905e-01
R43594 n3_20583_4751 n3_20583_4784 2.095238e-02
R43595 n3_20583_4784 n3_20583_4924 8.888889e-02
R43596 n3_20583_4924 n3_20583_4967 2.730159e-02
R43597 n3_20583_4967 n3_20583_5000 2.095238e-02
R43598 n3_20583_5000 n3_20583_5020 1.269841e-02
R43599 n3_20583_5020 n3_20583_5183 1.034921e-01
R43600 n3_20583_5183 n3_20583_5216 2.095238e-02
R43601 n3_20583_5216 n3_20583_5399 1.161905e-01
R43602 n3_20583_5399 n3_20583_5432 2.095238e-02
R43603 n3_20583_5432 n3_20583_5615 1.161905e-01
R43604 n3_20583_5615 n3_20583_5648 2.095238e-02
R43605 n3_20583_5648 n3_20583_5782 8.507937e-02
R43606 n3_20583_5782 n3_20583_5831 3.111111e-02
R43607 n3_20583_5831 n3_20583_5864 2.095238e-02
R43608 n3_20583_6263 n3_20583_6296 2.095238e-02
R43609 n3_20583_6296 n3_20583_6333 2.349206e-02
R43610 n3_20583_6333 n3_20583_6479 9.269841e-02
R43611 n3_20583_6479 n3_20583_6512 2.095238e-02
R43612 n3_20583_6512 n3_20583_6695 1.161905e-01
R43613 n3_20583_6695 n3_20583_6728 2.095238e-02
R43614 n3_20583_6728 n3_20583_6911 1.161905e-01
R43615 n3_20583_6911 n3_20583_6944 2.095238e-02
R43616 n3_20583_6944 n3_20583_7127 1.161905e-01
R43617 n3_20583_7127 n3_20583_7160 2.095238e-02
R43618 n3_20583_7160 n3_20583_7174 8.888889e-03
R43619 n3_20583_7174 n3_20583_7270 6.095238e-02
R43620 n3_20583_7270 n3_20583_7343 4.634921e-02
R43621 n3_20583_7343 n3_20583_7376 2.095238e-02
R43622 n3_20583_7376 n3_20583_7559 1.161905e-01
R43623 n3_20583_7559 n3_20583_7592 2.095238e-02
R43624 n3_20583_7592 n3_20583_7775 1.161905e-01
R43625 n3_20583_7775 n3_20583_7808 2.095238e-02
R43626 n3_20583_7808 n3_20583_7991 1.161905e-01
R43627 n3_20583_7991 n3_20583_8024 2.095238e-02
R43628 n3_20583_8024 n3_20583_8207 1.161905e-01
R43629 n3_20583_8207 n3_20583_8240 2.095238e-02
R43630 n3_20583_8456 n3_20583_8639 1.161905e-01
R43631 n3_20583_8639 n3_20583_8672 2.095238e-02
R43632 n3_20583_8672 n3_20583_8855 1.161905e-01
R43633 n3_20583_8855 n3_20583_8888 2.095238e-02
R43634 n3_20583_8888 n3_20583_9071 1.161905e-01
R43635 n3_20583_9071 n3_20583_9104 2.095238e-02
R43636 n3_20583_9104 n3_20583_9287 1.161905e-01
R43637 n3_20583_9287 n3_20583_9320 2.095238e-02
R43638 n3_20583_9320 n3_20583_9424 6.603175e-02
R43639 n3_20583_9424 n3_20583_9503 5.015873e-02
R43640 n3_20583_9503 n3_20583_9520 1.079365e-02
R43641 n3_20583_9520 n3_20583_9536 1.015873e-02
R43642 n3_20583_9536 n3_20583_9719 1.161905e-01
R43643 n3_20583_9719 n3_20583_9752 2.095238e-02
R43644 n3_20583_9752 n3_20583_9935 1.161905e-01
R43645 n3_20583_9935 n3_20583_9968 2.095238e-02
R43646 n3_20583_9968 n3_20583_10151 1.161905e-01
R43647 n3_20583_10151 n3_20583_10184 2.095238e-02
R43648 n3_20583_10184 n3_20583_10367 1.161905e-01
R43649 n3_20583_10367 n3_20583_10400 2.095238e-02
R43650 n3_20583_10799 n3_20583_10832 2.095238e-02
R43651 n3_20583_10832 n3_20583_11015 1.161905e-01
R43652 n3_20583_11015 n3_20583_11048 2.095238e-02
R43653 n3_20583_11048 n3_20583_11231 1.161905e-01
R43654 n3_20583_11231 n3_20583_11264 2.095238e-02
R43655 n3_20583_11264 n3_20583_11447 1.161905e-01
R43656 n3_20583_11447 n3_20583_11480 2.095238e-02
R43657 n3_20583_11480 n3_20583_11663 1.161905e-01
R43658 n3_20583_11663 n3_20583_11674 6.984127e-03
R43659 n3_20583_11674 n3_20583_11696 1.396825e-02
R43660 n3_20583_11696 n3_20583_11770 4.698413e-02
R43661 n3_20583_11770 n3_20583_11879 6.920635e-02
R43662 n3_20583_11879 n3_20583_11912 2.095238e-02
R43663 n3_20583_11912 n3_20583_12095 1.161905e-01
R43664 n3_20583_12095 n3_20583_12128 2.095238e-02
R43665 n3_20583_12128 n3_20583_12311 1.161905e-01
R43666 n3_20583_12311 n3_20583_12344 2.095238e-02
R43667 n3_20583_12344 n3_20583_12527 1.161905e-01
R43668 n3_20583_12527 n3_20583_12560 2.095238e-02
R43669 n3_20583_12560 n3_20583_12743 1.161905e-01
R43670 n3_20583_12959 n3_20583_12992 2.095238e-02
R43671 n3_20583_12992 n3_20583_13175 1.161905e-01
R43672 n3_20583_13175 n3_20583_13208 2.095238e-02
R43673 n3_20583_13208 n3_20583_13391 1.161905e-01
R43674 n3_20583_13391 n3_20583_13424 2.095238e-02
R43675 n3_20583_13424 n3_20583_13607 1.161905e-01
R43676 n3_20583_13607 n3_20583_13640 2.095238e-02
R43677 n3_20583_13640 n3_20583_13823 1.161905e-01
R43678 n3_20583_13823 n3_20583_13856 2.095238e-02
R43679 n3_20583_13856 n3_20583_13924 4.317460e-02
R43680 n3_20583_13924 n3_20583_14020 6.095238e-02
R43681 n3_20583_14020 n3_20583_14039 1.206349e-02
R43682 n3_20583_14039 n3_20583_14072 2.095238e-02
R43683 n3_20583_14072 n3_20583_14255 1.161905e-01
R43684 n3_20583_14255 n3_20583_14288 2.095238e-02
R43685 n3_20583_14288 n3_20583_14471 1.161905e-01
R43686 n3_20583_14471 n3_20583_14504 2.095238e-02
R43687 n3_20583_14504 n3_20583_14687 1.161905e-01
R43688 n3_20583_14687 n3_20583_14720 2.095238e-02
R43689 n3_20583_14720 n3_20583_14903 1.161905e-01
R43690 n3_20583_14903 n3_20583_14936 2.095238e-02
R43691 n3_20583_15308 n3_20583_15335 1.714286e-02
R43692 n3_20583_15335 n3_20583_15368 2.095238e-02
R43693 n3_20583_15368 n3_20583_15551 1.161905e-01
R43694 n3_20583_15551 n3_20583_15584 2.095238e-02
R43695 n3_20583_15584 n3_20583_15767 1.161905e-01
R43696 n3_20583_15767 n3_20583_15800 2.095238e-02
R43697 n3_20583_15800 n3_20583_15983 1.161905e-01
R43698 n3_20583_15983 n3_20583_16016 2.095238e-02
R43699 n3_20583_16016 n3_20583_16174 1.003175e-01
R43700 n3_20583_16174 n3_20583_16199 1.587302e-02
R43701 n3_20583_16199 n3_20583_16232 2.095238e-02
R43702 n3_20583_16232 n3_20583_16270 2.412698e-02
R43703 n3_20583_16270 n3_20583_16415 9.206349e-02
R43704 n3_20583_16415 n3_20583_16448 2.095238e-02
R43705 n3_20583_16448 n3_20583_16631 1.161905e-01
R43706 n3_20583_16631 n3_20583_16664 2.095238e-02
R43707 n3_20583_16664 n3_20583_16798 8.507937e-02
R43708 n3_20583_16798 n3_20583_16847 3.111111e-02
R43709 n3_20583_16847 n3_20583_16880 2.095238e-02
R43710 n3_20583_16880 n3_20583_17063 1.161905e-01
R43711 n3_20583_17063 n3_20583_17096 2.095238e-02
R43712 n3_20583_17495 n3_20583_17528 2.095238e-02
R43713 n3_20583_17528 n3_20583_17711 1.161905e-01
R43714 n3_20583_17711 n3_20583_17744 2.095238e-02
R43715 n3_20583_17744 n3_20583_17927 1.161905e-01
R43716 n3_20583_17927 n3_20583_17960 2.095238e-02
R43717 n3_20583_17960 n3_20583_18143 1.161905e-01
R43718 n3_20583_18143 n3_20583_18176 2.095238e-02
R43719 n3_20583_18176 n3_20583_18359 1.161905e-01
R43720 n3_20583_18359 n3_20583_18392 2.095238e-02
R43721 n3_20583_18392 n3_20583_18424 2.031746e-02
R43722 n3_20583_18424 n3_20583_18520 6.095238e-02
R43723 n3_20583_18520 n3_20583_18527 4.444444e-03
R43724 n3_20583_18527 n3_20583_18575 3.047619e-02
R43725 n3_20583_18575 n3_20583_18608 2.095238e-02
R43726 n3_20583_18608 n3_20583_18791 1.161905e-01
R43727 n3_20583_18791 n3_20583_18824 2.095238e-02
R43728 n3_20583_18824 n3_20583_19007 1.161905e-01
R43729 n3_20583_19007 n3_20583_19040 2.095238e-02
R43730 n3_20583_19040 n3_20583_19223 1.161905e-01
R43731 n3_20583_19223 n3_20583_19256 2.095238e-02
R43732 n3_20583_19256 n3_20583_19439 1.161905e-01
R43733 n3_20583_19439 n3_20583_19472 2.095238e-02
R43734 n3_20583_19871 n3_20583_19904 2.095238e-02
R43735 n3_20583_19904 n3_20583_20087 1.161905e-01
R43736 n3_20583_20087 n3_20583_20120 2.095238e-02
R43737 n3_20583_20120 n3_20583_20303 1.161905e-01
R43738 n3_20583_20303 n3_20583_20336 2.095238e-02
R43739 n3_20583_20336 n3_20583_20519 1.161905e-01
R43740 n3_20583_20519 n3_20583_20552 2.095238e-02
R43741 n3_20583_20552 n3_20583_20674 7.746032e-02
R43742 n3_20583_20674 n3_20583_20687 8.253968e-03
R43743 n3_20583_20687 n3_20583_20735 3.047619e-02
R43744 n3_20583_20735 n3_20583_20768 2.095238e-02
R43745 n3_20583_20768 n3_20583_20770 1.269841e-03
R43746 n3_20583_20770 n3_20583_20951 1.149206e-01
R43747 n3_20583_20951 n3_20583_20984 2.095238e-02
R43748 n3_20771_520 n3_20771_647 8.063492e-02
R43749 n3_20771_647 n3_20771_680 2.095238e-02
R43750 n3_20771_680 n3_20771_863 1.161905e-01
R43751 n3_20771_863 n3_20771_896 2.095238e-02
R43752 n3_20771_896 n3_20771_1079 1.161905e-01
R43753 n3_20771_1079 n3_20771_1112 2.095238e-02
R43754 n3_20771_1112 n3_20771_1295 1.161905e-01
R43755 n3_20771_1295 n3_20771_1328 2.095238e-02
R43756 n3_20771_1328 n3_20771_1511 1.161905e-01
R43757 n3_20771_1511 n3_20771_1544 2.095238e-02
R43758 n3_20771_1544 n3_20771_1727 1.161905e-01
R43759 n3_20771_1727 n3_20771_1760 2.095238e-02
R43760 n3_20771_1760 n3_20771_1943 1.161905e-01
R43761 n3_20771_1943 n3_20771_1976 2.095238e-02
R43762 n3_20771_1976 n3_20771_2159 1.161905e-01
R43763 n3_20771_2159 n3_20771_2192 2.095238e-02
R43764 n3_20771_2192 n3_20771_2375 1.161905e-01
R43765 n3_20771_2375 n3_20771_2408 2.095238e-02
R43766 n3_20771_2408 n3_20771_2543 8.571429e-02
R43767 n3_20771_2543 n3_20771_2591 3.047619e-02
R43768 n3_20771_2591 n3_20771_2624 2.095238e-02
R43769 n3_20771_2624 n3_20771_2674 3.174603e-02
R43770 n3_20771_2770 n3_20771_2807 2.349206e-02
R43771 n3_20771_2807 n3_20771_2840 2.095238e-02
R43772 n3_20771_2840 n3_20771_3023 1.161905e-01
R43773 n3_20771_3023 n3_20771_3056 2.095238e-02
R43774 n3_20771_3056 n3_20771_3239 1.161905e-01
R43775 n3_20771_3239 n3_20771_3272 2.095238e-02
R43776 n3_20771_3272 n3_20771_3455 1.161905e-01
R43777 n3_20771_3455 n3_20771_3488 2.095238e-02
R43778 n3_20771_3488 n3_20771_3671 1.161905e-01
R43779 n3_20771_3671 n3_20771_3704 2.095238e-02
R43780 n3_20771_3704 n3_20771_3887 1.161905e-01
R43781 n3_20771_3887 n3_20771_3920 2.095238e-02
R43782 n3_20771_3920 n3_20771_4103 1.161905e-01
R43783 n3_20771_4103 n3_20771_4136 2.095238e-02
R43784 n3_20771_4136 n3_20771_4319 1.161905e-01
R43785 n3_20771_4319 n3_20771_4352 2.095238e-02
R43786 n3_20771_4352 n3_20771_4535 1.161905e-01
R43787 n3_20771_4535 n3_20771_4568 2.095238e-02
R43788 n3_20771_4568 n3_20771_4751 1.161905e-01
R43789 n3_20771_4751 n3_20771_4784 2.095238e-02
R43790 n3_20771_4784 n3_20771_4924 8.888889e-02
R43791 n3_20771_5000 n3_20771_5020 1.269841e-02
R43792 n3_20771_5020 n3_20771_5183 1.034921e-01
R43793 n3_20771_5183 n3_20771_5216 2.095238e-02
R43794 n3_20771_5216 n3_20771_5399 1.161905e-01
R43795 n3_20771_5399 n3_20771_5432 2.095238e-02
R43796 n3_20771_5432 n3_20771_5615 1.161905e-01
R43797 n3_20771_5615 n3_20771_5648 2.095238e-02
R43798 n3_20771_5648 n3_20771_5782 8.507937e-02
R43799 n3_20771_5782 n3_20771_5831 3.111111e-02
R43800 n3_20771_5831 n3_20771_5864 2.095238e-02
R43801 n3_20771_5864 n3_20771_6047 1.161905e-01
R43802 n3_20771_6047 n3_20771_6080 2.095238e-02
R43803 n3_20771_6080 n3_20771_6263 1.161905e-01
R43804 n3_20771_6263 n3_20771_6296 2.095238e-02
R43805 n3_20771_6296 n3_20771_6479 1.161905e-01
R43806 n3_20771_6479 n3_20771_6512 2.095238e-02
R43807 n3_20771_6512 n3_20771_6695 1.161905e-01
R43808 n3_20771_6695 n3_20771_6728 2.095238e-02
R43809 n3_20771_6728 n3_20771_6911 1.161905e-01
R43810 n3_20771_6911 n3_20771_6944 2.095238e-02
R43811 n3_20771_6944 n3_20771_7127 1.161905e-01
R43812 n3_20771_7127 n3_20771_7160 2.095238e-02
R43813 n3_20771_7160 n3_20771_7174 8.888889e-03
R43814 n3_20771_7270 n3_20771_7343 4.634921e-02
R43815 n3_20771_7343 n3_20771_7376 2.095238e-02
R43816 n3_20771_7376 n3_20771_7559 1.161905e-01
R43817 n3_20771_7559 n3_20771_7592 2.095238e-02
R43818 n3_20771_7592 n3_20771_7775 1.161905e-01
R43819 n3_20771_7775 n3_20771_7808 2.095238e-02
R43820 n3_20771_7808 n3_20771_7991 1.161905e-01
R43821 n3_20771_7991 n3_20771_8024 2.095238e-02
R43822 n3_20771_8024 n3_20771_8207 1.161905e-01
R43823 n3_20771_8207 n3_20771_8240 2.095238e-02
R43824 n3_20771_8240 n3_20771_8423 1.161905e-01
R43825 n3_20771_8423 n3_20771_8456 2.095238e-02
R43826 n3_20771_8456 n3_20771_8639 1.161905e-01
R43827 n3_20771_8639 n3_20771_8672 2.095238e-02
R43828 n3_20771_8672 n3_20771_8855 1.161905e-01
R43829 n3_20771_8855 n3_20771_8888 2.095238e-02
R43830 n3_20771_8888 n3_20771_9071 1.161905e-01
R43831 n3_20771_9071 n3_20771_9104 2.095238e-02
R43832 n3_20771_9104 n3_20771_9287 1.161905e-01
R43833 n3_20771_9287 n3_20771_9320 2.095238e-02
R43834 n3_20771_9320 n3_20771_9424 6.603175e-02
R43835 n3_20771_9503 n3_20771_9520 1.079365e-02
R43836 n3_20771_9520 n3_20771_9536 1.015873e-02
R43837 n3_20771_9536 n3_20771_9719 1.161905e-01
R43838 n3_20771_9719 n3_20771_9752 2.095238e-02
R43839 n3_20771_9752 n3_20771_9935 1.161905e-01
R43840 n3_20771_9935 n3_20771_9968 2.095238e-02
R43841 n3_20771_9968 n3_20771_10151 1.161905e-01
R43842 n3_20771_10151 n3_20771_10184 2.095238e-02
R43843 n3_20771_10184 n3_20771_10367 1.161905e-01
R43844 n3_20771_10367 n3_20771_10400 2.095238e-02
R43845 n3_20771_10616 n3_20771_10799 1.161905e-01
R43846 n3_20771_10799 n3_20771_10832 2.095238e-02
R43847 n3_20771_10832 n3_20771_11015 1.161905e-01
R43848 n3_20771_11015 n3_20771_11048 2.095238e-02
R43849 n3_20771_11048 n3_20771_11231 1.161905e-01
R43850 n3_20771_11231 n3_20771_11264 2.095238e-02
R43851 n3_20771_11264 n3_20771_11447 1.161905e-01
R43852 n3_20771_11447 n3_20771_11480 2.095238e-02
R43853 n3_20771_11480 n3_20771_11663 1.161905e-01
R43854 n3_20771_11663 n3_20771_11674 6.984127e-03
R43855 n3_20771_11674 n3_20771_11696 1.396825e-02
R43856 n3_20771_11770 n3_20771_11879 6.920635e-02
R43857 n3_20771_11879 n3_20771_11912 2.095238e-02
R43858 n3_20771_11912 n3_20771_12095 1.161905e-01
R43859 n3_20771_12095 n3_20771_12128 2.095238e-02
R43860 n3_20771_12128 n3_20771_12311 1.161905e-01
R43861 n3_20771_12311 n3_20771_12344 2.095238e-02
R43862 n3_20771_12344 n3_20771_12527 1.161905e-01
R43863 n3_20771_12527 n3_20771_12560 2.095238e-02
R43864 n3_20771_12560 n3_20771_12743 1.161905e-01
R43865 n3_20771_12743 n3_20771_12776 2.095238e-02
R43866 n3_20771_12776 n3_20771_12959 1.161905e-01
R43867 n3_20771_12959 n3_20771_12992 2.095238e-02
R43868 n3_20771_12992 n3_20771_13175 1.161905e-01
R43869 n3_20771_13175 n3_20771_13208 2.095238e-02
R43870 n3_20771_13208 n3_20771_13391 1.161905e-01
R43871 n3_20771_13391 n3_20771_13424 2.095238e-02
R43872 n3_20771_13424 n3_20771_13607 1.161905e-01
R43873 n3_20771_13607 n3_20771_13640 2.095238e-02
R43874 n3_20771_13640 n3_20771_13823 1.161905e-01
R43875 n3_20771_13823 n3_20771_13856 2.095238e-02
R43876 n3_20771_13856 n3_20771_13924 4.317460e-02
R43877 n3_20771_14020 n3_20771_14039 1.206349e-02
R43878 n3_20771_14039 n3_20771_14072 2.095238e-02
R43879 n3_20771_14072 n3_20771_14255 1.161905e-01
R43880 n3_20771_14255 n3_20771_14288 2.095238e-02
R43881 n3_20771_14288 n3_20771_14471 1.161905e-01
R43882 n3_20771_14471 n3_20771_14504 2.095238e-02
R43883 n3_20771_14504 n3_20771_14687 1.161905e-01
R43884 n3_20771_14687 n3_20771_14720 2.095238e-02
R43885 n3_20771_14720 n3_20771_14903 1.161905e-01
R43886 n3_20771_14903 n3_20771_14936 2.095238e-02
R43887 n3_20771_14936 n3_20771_15092 9.904762e-02
R43888 n3_20771_15092 n3_20771_15119 1.714286e-02
R43889 n3_20771_15119 n3_20771_15152 2.095238e-02
R43890 n3_20771_15152 n3_20771_15308 9.904762e-02
R43891 n3_20771_15308 n3_20771_15335 1.714286e-02
R43892 n3_20771_15335 n3_20771_15368 2.095238e-02
R43893 n3_20771_15368 n3_20771_15551 1.161905e-01
R43894 n3_20771_15551 n3_20771_15584 2.095238e-02
R43895 n3_20771_15584 n3_20771_15767 1.161905e-01
R43896 n3_20771_15767 n3_20771_15800 2.095238e-02
R43897 n3_20771_15800 n3_20771_15983 1.161905e-01
R43898 n3_20771_15983 n3_20771_16016 2.095238e-02
R43899 n3_20771_16016 n3_20771_16174 1.003175e-01
R43900 n3_20771_16174 n3_20771_16199 1.587302e-02
R43901 n3_20771_16270 n3_20771_16415 9.206349e-02
R43902 n3_20771_16415 n3_20771_16448 2.095238e-02
R43903 n3_20771_16448 n3_20771_16631 1.161905e-01
R43904 n3_20771_16631 n3_20771_16664 2.095238e-02
R43905 n3_20771_16664 n3_20771_16798 8.507937e-02
R43906 n3_20771_16798 n3_20771_16847 3.111111e-02
R43907 n3_20771_16847 n3_20771_16880 2.095238e-02
R43908 n3_20771_16880 n3_20771_17063 1.161905e-01
R43909 n3_20771_17063 n3_20771_17096 2.095238e-02
R43910 n3_20771_17096 n3_20771_17279 1.161905e-01
R43911 n3_20771_17279 n3_20771_17312 2.095238e-02
R43912 n3_20771_17312 n3_20771_17495 1.161905e-01
R43913 n3_20771_17495 n3_20771_17528 2.095238e-02
R43914 n3_20771_17528 n3_20771_17711 1.161905e-01
R43915 n3_20771_17711 n3_20771_17744 2.095238e-02
R43916 n3_20771_17744 n3_20771_17927 1.161905e-01
R43917 n3_20771_17927 n3_20771_17960 2.095238e-02
R43918 n3_20771_17960 n3_20771_18143 1.161905e-01
R43919 n3_20771_18143 n3_20771_18176 2.095238e-02
R43920 n3_20771_18176 n3_20771_18359 1.161905e-01
R43921 n3_20771_18359 n3_20771_18392 2.095238e-02
R43922 n3_20771_18392 n3_20771_18424 2.031746e-02
R43923 n3_20771_18520 n3_20771_18527 4.444444e-03
R43924 n3_20771_18527 n3_20771_18575 3.047619e-02
R43925 n3_20771_18575 n3_20771_18608 2.095238e-02
R43926 n3_20771_18608 n3_20771_18791 1.161905e-01
R43927 n3_20771_18791 n3_20771_18824 2.095238e-02
R43928 n3_20771_18824 n3_20771_19007 1.161905e-01
R43929 n3_20771_19007 n3_20771_19040 2.095238e-02
R43930 n3_20771_19040 n3_20771_19223 1.161905e-01
R43931 n3_20771_19223 n3_20771_19256 2.095238e-02
R43932 n3_20771_19256 n3_20771_19439 1.161905e-01
R43933 n3_20771_19439 n3_20771_19472 2.095238e-02
R43934 n3_20771_19472 n3_20771_19655 1.161905e-01
R43935 n3_20771_19655 n3_20771_19688 2.095238e-02
R43936 n3_20771_19688 n3_20771_19871 1.161905e-01
R43937 n3_20771_19871 n3_20771_19904 2.095238e-02
R43938 n3_20771_19904 n3_20771_20087 1.161905e-01
R43939 n3_20771_20087 n3_20771_20120 2.095238e-02
R43940 n3_20771_20120 n3_20771_20303 1.161905e-01
R43941 n3_20771_20303 n3_20771_20336 2.095238e-02
R43942 n3_20771_20336 n3_20771_20519 1.161905e-01
R43943 n3_20771_20519 n3_20771_20552 2.095238e-02
R43944 n3_20771_20552 n3_20771_20674 7.746032e-02
R43945 n3_20771_20674 n3_20771_20687 8.253968e-03
R43946 n3_9380_20674 n3_9380_20687 2.600000e-02
R43947 n3_9380_20687 n3_9380_20721 6.800000e-02
R43948 n3_9380_20721 n3_9380_20735 2.800000e-02
R43949 n3_9380_20735 n3_9380_20768 6.600000e-02
R43950 n3_9380_20768 n3_9380_20770 4.000000e-03
R43951 n3_9380_18392 n3_9380_18424 6.400000e-02
R43952 n3_9380_18424 n3_9380_18471 9.400000e-02
R43953 n3_9380_18471 n3_9380_18520 9.800000e-02
R43954 n3_9380_18520 n3_9380_18527 1.400000e-02
R43955 n3_9380_18527 n3_9380_18548 4.200000e-02
R43956 n3_9380_16172 n3_9380_16174 4.000000e-03
R43957 n3_9380_16174 n3_9380_16199 5.000000e-02
R43958 n3_9380_16199 n3_9380_16221 4.400000e-02
R43959 n3_9380_16221 n3_9380_16232 2.200000e-02
R43960 n3_9380_16232 n3_9380_16270 7.600000e-02
R43961 n3_9380_13924 n3_9380_13971 9.400000e-02
R43962 n3_9380_13971 n3_9380_13990 3.800000e-02
R43963 n3_9380_13990 n3_9380_14012 4.400000e-02
R43964 n3_9380_14012 n3_9380_14020 1.600000e-02
R43965 n3_9380_14020 n3_9380_14039 3.800000e-02
R43966 n3_7130_20674 n3_7130_20687 2.600000e-02
R43967 n3_7130_20687 n3_7130_20721 6.800000e-02
R43968 n3_7130_20721 n3_7130_20735 2.800000e-02
R43969 n3_7130_20735 n3_7130_20768 6.600000e-02
R43970 n3_7130_20768 n3_7130_20770 4.000000e-03
R43971 n3_7130_18392 n3_7130_18424 6.400000e-02
R43972 n3_7130_18424 n3_7130_18471 9.400000e-02
R43973 n3_7130_18471 n3_7130_18520 9.800000e-02
R43974 n3_7130_18520 n3_7130_18526 1.200000e-02
R43975 n3_7130_18526 n3_7130_18527 2.000000e-03
R43976 n3_7130_18527 n3_7130_18548 4.200000e-02
R43977 n3_7130_16172 n3_7130_16174 4.000000e-03
R43978 n3_7130_16174 n3_7130_16199 5.000000e-02
R43979 n3_7130_16199 n3_7130_16221 4.400000e-02
R43980 n3_7130_16221 n3_7130_16232 2.200000e-02
R43981 n3_7130_16232 n3_7130_16270 7.600000e-02
R43982 n3_4880_20674 n3_4880_20687 2.600000e-02
R43983 n3_4880_20687 n3_4880_20721 6.800000e-02
R43984 n3_4880_20721 n3_4880_20735 2.800000e-02
R43985 n3_4880_20735 n3_4880_20768 6.600000e-02
R43986 n3_4880_20768 n3_4880_20770 4.000000e-03
R43987 n3_4880_18392 n3_4880_18424 6.400000e-02
R43988 n3_4880_18424 n3_4880_18471 9.400000e-02
R43989 n3_4880_18471 n3_4880_18520 9.800000e-02
R43990 n3_4880_18520 n3_4880_18527 1.400000e-02
R43991 n3_4880_18527 n3_4880_18548 4.200000e-02
R43992 n3_2630_20674 n3_2630_20687 2.600000e-02
R43993 n3_2630_20687 n3_2630_20721 6.800000e-02
R43994 n3_2630_20721 n3_2630_20735 2.800000e-02
R43995 n3_2630_20735 n3_2630_20768 6.600000e-02
R43996 n3_2630_20768 n3_2630_20770 4.000000e-03
R43997 n3_380_20674 n3_380_20687 2.600000e-02
R43998 n3_380_20687 n3_380_20721 6.800000e-02
R43999 n3_380_20721 n3_380_20735 2.800000e-02
R44000 n3_380_20735 n3_380_20768 6.600000e-02
R44001 n3_380_20768 n3_380_20770 4.000000e-03
R44002 n3_380_18392 n3_380_18424 6.400000e-02
R44003 n3_380_18424 n3_380_18471 9.400000e-02
R44004 n3_380_18471 n3_380_18520 9.800000e-02
R44005 n3_380_18520 n3_380_18527 1.400000e-02
R44006 n3_2630_18392 n3_2630_18424 6.400000e-02
R44007 n3_2630_18424 n3_2630_18471 9.400000e-02
R44008 n3_2630_18471 n3_2630_18520 9.800000e-02
R44009 n3_2630_18520 n3_2630_18527 1.400000e-02
R44010 n3_380_16174 n3_380_16199 5.000000e-02
R44011 n3_380_16199 n3_380_16221 4.400000e-02
R44012 n3_380_16221 n3_380_16232 2.200000e-02
R44013 n3_380_16232 n3_380_16270 7.600000e-02
R44014 n3_2630_16174 n3_2630_16199 5.000000e-02
R44015 n3_2630_16199 n3_2630_16221 4.400000e-02
R44016 n3_2630_16221 n3_2630_16232 2.200000e-02
R44017 n3_2630_16232 n3_2630_16270 7.600000e-02
R44018 n3_4880_16172 n3_4880_16174 4.000000e-03
R44019 n3_4880_16174 n3_4880_16199 5.000000e-02
R44020 n3_4880_16199 n3_4880_16221 4.400000e-02
R44021 n3_4880_16221 n3_4880_16232 2.200000e-02
R44022 n3_4880_16232 n3_4880_16270 7.600000e-02
R44023 n3_380_13924 n3_380_13971 9.400000e-02
R44024 n3_380_13971 n3_380_14020 9.800000e-02
R44025 n3_380_14020 n3_380_14039 3.800000e-02
R44026 n3_2630_13924 n3_2630_13971 9.400000e-02
R44027 n3_2630_13971 n3_2630_13990 3.800000e-02
R44028 n3_2630_13990 n3_2630_14020 6.000000e-02
R44029 n3_2630_14020 n3_2630_14039 3.800000e-02
R44030 n3_4880_13924 n3_4880_13971 9.400000e-02
R44031 n3_4880_13971 n3_4880_13990 3.800000e-02
R44032 n3_4880_13990 n3_4880_14020 6.000000e-02
R44033 n3_4880_14020 n3_4880_14039 3.800000e-02
R44034 n3_7130_13924 n3_7130_13971 9.400000e-02
R44035 n3_7130_13971 n3_7130_14020 9.800000e-02
R44036 n3_7130_14020 n3_7130_14039 3.800000e-02
R44037 n3_380_11663 n3_380_11674 2.200000e-02
R44038 n3_380_11674 n3_380_11696 4.400000e-02
R44039 n3_380_11696 n3_380_11721 5.000000e-02
R44040 n3_380_11721 n3_380_11770 9.800000e-02
R44041 n3_2630_11663 n3_2630_11674 2.200000e-02
R44042 n3_2630_11674 n3_2630_11696 4.400000e-02
R44043 n3_2630_11696 n3_2630_11721 5.000000e-02
R44044 n3_2630_11721 n3_2630_11770 9.800000e-02
R44045 n3_4880_11663 n3_4880_11674 2.200000e-02
R44046 n3_4880_11674 n3_4880_11696 4.400000e-02
R44047 n3_4880_11696 n3_4880_11721 5.000000e-02
R44048 n3_4880_11721 n3_4880_11770 9.800000e-02
R44049 n3_7130_11663 n3_7130_11674 2.200000e-02
R44050 n3_7130_11674 n3_7130_11696 4.400000e-02
R44051 n3_7130_11696 n3_7130_11721 5.000000e-02
R44052 n3_7130_11721 n3_7130_11770 9.800000e-02
R44053 n3_9380_11663 n3_9380_11674 2.200000e-02
R44054 n3_9380_11674 n3_9380_11696 4.400000e-02
R44055 n3_9380_11696 n3_9380_11721 5.000000e-02
R44056 n3_9380_11721 n3_9380_11770 9.800000e-02
R44057 n3_380_424 n3_380_431 1.400000e-02
R44058 n3_380_431 n3_380_464 6.600000e-02
R44059 n3_380_464 n3_380_471 1.400000e-02
R44060 n3_380_471 n3_380_520 9.800000e-02
R44061 n3_2630_424 n3_2630_431 1.400000e-02
R44062 n3_2630_431 n3_2630_464 6.600000e-02
R44063 n3_2630_464 n3_2630_471 1.400000e-02
R44064 n3_2630_471 n3_2630_520 9.800000e-02
R44065 n3_2630_2674 n3_2630_2721 9.400000e-02
R44066 n3_2630_2721 n3_2630_2770 9.800000e-02
R44067 n3_4880_424 n3_4880_431 1.400000e-02
R44068 n3_4880_431 n3_4880_464 6.600000e-02
R44069 n3_4880_464 n3_4880_471 1.400000e-02
R44070 n3_4880_471 n3_4880_513 8.400000e-02
R44071 n3_4880_513 n3_4880_520 1.400000e-02
R44072 n3_4880_2674 n3_4880_2721 9.400000e-02
R44073 n3_4880_2721 n3_4880_2770 9.800000e-02
R44074 n3_4880_4924 n3_4880_4967 8.600000e-02
R44075 n3_4880_4967 n3_4880_4971 8.000000e-03
R44076 n3_4880_4971 n3_4880_5000 5.800000e-02
R44077 n3_4880_5000 n3_4880_5020 4.000000e-02
R44078 n3_7130_424 n3_7130_431 1.400000e-02
R44079 n3_7130_431 n3_7130_464 6.600000e-02
R44080 n3_7130_464 n3_7130_471 1.400000e-02
R44081 n3_7130_471 n3_7130_520 9.800000e-02
R44082 n3_7130_2674 n3_7130_2721 9.400000e-02
R44083 n3_7130_2721 n3_7130_2770 9.800000e-02
R44084 n3_7130_4924 n3_7130_4967 8.600000e-02
R44085 n3_7130_4967 n3_7130_4971 8.000000e-03
R44086 n3_7130_4971 n3_7130_5000 5.800000e-02
R44087 n3_7130_5000 n3_7130_5020 4.000000e-02
R44088 n3_7130_7160 n3_7130_7174 2.800000e-02
R44089 n3_7130_7174 n3_7130_7221 9.400000e-02
R44090 n3_7130_7221 n3_7130_7270 9.800000e-02
R44091 n3_9380_424 n3_9380_431 1.400000e-02
R44092 n3_9380_431 n3_9380_464 6.600000e-02
R44093 n3_9380_464 n3_9380_471 1.400000e-02
R44094 n3_9380_471 n3_9380_520 9.800000e-02
R44095 n3_9380_2674 n3_9380_2721 9.400000e-02
R44096 n3_9380_2721 n3_9380_2770 9.800000e-02
R44097 n3_9380_4924 n3_9380_4967 8.600000e-02
R44098 n3_9380_4967 n3_9380_4971 8.000000e-03
R44099 n3_9380_4971 n3_9380_5000 5.800000e-02
R44100 n3_9380_5000 n3_9380_5020 4.000000e-02
R44101 n3_9380_7160 n3_9380_7174 2.800000e-02
R44102 n3_9380_7174 n3_9380_7221 9.400000e-02
R44103 n3_9380_7221 n3_9380_7270 9.800000e-02
R44104 n3_9380_9424 n3_9380_9471 9.400000e-02
R44105 n3_9380_9471 n3_9380_9503 6.400000e-02
R44106 n3_9380_9503 n3_9380_9520 3.400000e-02
R44107 n3_9380_9520 n3_9380_9536 3.200000e-02
R44108 n3_380_9424 n3_380_9471 9.400000e-02
R44109 n3_380_9471 n3_380_9503 6.400000e-02
R44110 n3_380_9503 n3_380_9520 3.400000e-02
R44111 n3_380_9520 n3_380_9536 3.200000e-02
R44112 n3_2630_9424 n3_2630_9471 9.400000e-02
R44113 n3_2630_9471 n3_2630_9503 6.400000e-02
R44114 n3_2630_9503 n3_2630_9520 3.400000e-02
R44115 n3_2630_9520 n3_2630_9536 3.200000e-02
R44116 n3_4880_9424 n3_4880_9471 9.400000e-02
R44117 n3_4880_9471 n3_4880_9503 6.400000e-02
R44118 n3_4880_9503 n3_4880_9520 3.400000e-02
R44119 n3_4880_9520 n3_4880_9536 3.200000e-02
R44120 n3_7130_9424 n3_7130_9471 9.400000e-02
R44121 n3_7130_9471 n3_7130_9503 6.400000e-02
R44122 n3_7130_9503 n3_7130_9520 3.400000e-02
R44123 n3_7130_9520 n3_7130_9536 3.200000e-02
R44124 n3_380_7160 n3_380_7174 2.800000e-02
R44125 n3_380_7174 n3_380_7221 9.400000e-02
R44126 n3_380_7221 n3_380_7270 9.800000e-02
R44127 n3_2630_7160 n3_2630_7174 2.800000e-02
R44128 n3_2630_7174 n3_2630_7221 9.400000e-02
R44129 n3_2630_7221 n3_2630_7270 9.800000e-02
R44130 n3_4880_7160 n3_4880_7174 2.800000e-02
R44131 n3_4880_7174 n3_4880_7221 9.400000e-02
R44132 n3_4880_7221 n3_4880_7270 9.800000e-02
R44133 n3_380_4924 n3_380_4967 8.600000e-02
R44134 n3_380_4967 n3_380_4971 8.000000e-03
R44135 n3_380_4971 n3_380_5000 5.800000e-02
R44136 n3_380_5000 n3_380_5020 4.000000e-02
R44137 n3_2630_4924 n3_2630_4967 8.600000e-02
R44138 n3_2630_4967 n3_2630_4971 8.000000e-03
R44139 n3_2630_4971 n3_2630_5000 5.800000e-02
R44140 n3_2630_5000 n3_2630_5020 4.000000e-02
R44141 n3_380_2674 n3_380_2721 9.400000e-02
R44142 n3_380_2721 n3_380_2770 9.800000e-02
R44143 n3_11630_424 n3_11630_431 1.400000e-02
R44144 n3_11630_431 n3_11630_464 6.600000e-02
R44145 n3_11630_464 n3_11630_471 1.400000e-02
R44146 n3_11630_471 n3_11630_520 9.800000e-02
R44147 n3_11630_2674 n3_11630_2721 9.400000e-02
R44148 n3_11630_2721 n3_11630_2760 7.800000e-02
R44149 n3_11630_2760 n3_11630_2770 2.000000e-02
R44150 n3_11630_4924 n3_11630_4967 8.600000e-02
R44151 n3_11630_4967 n3_11630_4971 8.000000e-03
R44152 n3_11630_4971 n3_11630_5000 5.800000e-02
R44153 n3_11630_5000 n3_11630_5020 4.000000e-02
R44154 n3_11630_7160 n3_11630_7174 2.800000e-02
R44155 n3_11630_7174 n3_11630_7221 9.400000e-02
R44156 n3_11630_7221 n3_11630_7270 9.800000e-02
R44157 n3_11630_7270 n3_11630_7294 4.800000e-02
R44158 n3_13880_424 n3_13880_431 1.400000e-02
R44159 n3_13880_431 n3_13880_464 6.600000e-02
R44160 n3_13880_464 n3_13880_471 1.400000e-02
R44161 n3_13880_471 n3_13880_520 9.800000e-02
R44162 n3_13880_2674 n3_13880_2721 9.400000e-02
R44163 n3_13880_2721 n3_13880_2770 9.800000e-02
R44164 n3_13880_4924 n3_13880_4967 8.600000e-02
R44165 n3_13880_4967 n3_13880_4971 8.000000e-03
R44166 n3_13880_4971 n3_13880_5000 5.800000e-02
R44167 n3_13880_5000 n3_13880_5020 4.000000e-02
R44168 n3_16130_424 n3_16130_431 1.400000e-02
R44169 n3_16130_431 n3_16130_464 6.600000e-02
R44170 n3_16130_464 n3_16130_471 1.400000e-02
R44171 n3_16130_471 n3_16130_520 9.800000e-02
R44172 n3_16130_2674 n3_16130_2721 9.400000e-02
R44173 n3_16130_2721 n3_16130_2770 9.800000e-02
R44174 n3_18380_424 n3_18380_431 1.400000e-02
R44175 n3_18380_431 n3_18380_464 6.600000e-02
R44176 n3_18380_464 n3_18380_471 1.400000e-02
R44177 n3_18380_471 n3_18380_520 9.800000e-02
R44178 n3_20630_424 n3_20630_431 1.400000e-02
R44179 n3_20630_431 n3_20630_464 6.600000e-02
R44180 n3_20630_464 n3_20630_471 1.400000e-02
R44181 n3_20630_471 n3_20630_520 9.800000e-02
R44182 n3_20630_2674 n3_20630_2721 9.400000e-02
R44183 n3_20630_2721 n3_20630_2770 9.800000e-02
R44184 n3_18380_2674 n3_18380_2721 9.400000e-02
R44185 n3_18380_2721 n3_18380_2770 9.800000e-02
R44186 n3_20630_4924 n3_20630_4967 8.600000e-02
R44187 n3_20630_4967 n3_20630_4971 8.000000e-03
R44188 n3_20630_4971 n3_20630_5000 5.800000e-02
R44189 n3_20630_5000 n3_20630_5020 4.000000e-02
R44190 n3_18380_4920 n3_18380_4924 8.000000e-03
R44191 n3_18380_4924 n3_18380_4967 8.600000e-02
R44192 n3_18380_4967 n3_18380_4971 8.000000e-03
R44193 n3_18380_4971 n3_18380_5000 5.800000e-02
R44194 n3_18380_5000 n3_18380_5020 4.000000e-02
R44195 n3_16130_4919 n3_16130_4924 1.000000e-02
R44196 n3_16130_4924 n3_16130_4967 8.600000e-02
R44197 n3_16130_4967 n3_16130_4971 8.000000e-03
R44198 n3_16130_4971 n3_16130_5000 5.800000e-02
R44199 n3_16130_5000 n3_16130_5020 4.000000e-02
R44200 n3_20630_7160 n3_20630_7174 2.800000e-02
R44201 n3_20630_7174 n3_20630_7221 9.400000e-02
R44202 n3_20630_7221 n3_20630_7270 9.800000e-02
R44203 n3_18380_7160 n3_18380_7174 2.800000e-02
R44204 n3_18380_7174 n3_18380_7221 9.400000e-02
R44205 n3_18380_7221 n3_18380_7270 9.800000e-02
R44206 n3_16130_7160 n3_16130_7174 2.800000e-02
R44207 n3_16130_7174 n3_16130_7221 9.400000e-02
R44208 n3_16130_7221 n3_16130_7270 9.800000e-02
R44209 n3_13880_7160 n3_13880_7174 2.800000e-02
R44210 n3_13880_7174 n3_13880_7221 9.400000e-02
R44211 n3_13880_7221 n3_13880_7270 9.800000e-02
R44212 n3_20630_9424 n3_20630_9471 9.400000e-02
R44213 n3_20630_9471 n3_20630_9503 6.400000e-02
R44214 n3_20630_9503 n3_20630_9520 3.400000e-02
R44215 n3_20630_9520 n3_20630_9536 3.200000e-02
R44216 n3_18380_9424 n3_18380_9471 9.400000e-02
R44217 n3_18380_9471 n3_18380_9503 6.400000e-02
R44218 n3_18380_9503 n3_18380_9520 3.400000e-02
R44219 n3_18380_9520 n3_18380_9536 3.200000e-02
R44220 n3_16130_9424 n3_16130_9471 9.400000e-02
R44221 n3_16130_9471 n3_16130_9503 6.400000e-02
R44222 n3_16130_9503 n3_16130_9520 3.400000e-02
R44223 n3_16130_9520 n3_16130_9536 3.200000e-02
R44224 n3_13880_9424 n3_13880_9471 9.400000e-02
R44225 n3_13880_9471 n3_13880_9503 6.400000e-02
R44226 n3_13880_9503 n3_13880_9520 3.400000e-02
R44227 n3_13880_9520 n3_13880_9536 3.200000e-02
R44228 n3_11630_9424 n3_11630_9471 9.400000e-02
R44229 n3_11630_9471 n3_11630_9503 6.400000e-02
R44230 n3_11630_9503 n3_11630_9520 3.400000e-02
R44231 n3_11630_9520 n3_11630_9536 3.200000e-02
R44232 n3_20630_11663 n3_20630_11674 2.200000e-02
R44233 n3_20630_11674 n3_20630_11696 4.400000e-02
R44234 n3_20630_11696 n3_20630_11721 5.000000e-02
R44235 n3_20630_11721 n3_20630_11770 9.800000e-02
R44236 n3_18380_11663 n3_18380_11674 2.200000e-02
R44237 n3_18380_11674 n3_18380_11696 4.400000e-02
R44238 n3_18380_11696 n3_18380_11721 5.000000e-02
R44239 n3_18380_11721 n3_18380_11770 9.800000e-02
R44240 n3_16130_11663 n3_16130_11674 2.200000e-02
R44241 n3_16130_11674 n3_16130_11696 4.400000e-02
R44242 n3_16130_11696 n3_16130_11721 5.000000e-02
R44243 n3_16130_11721 n3_16130_11770 9.800000e-02
R44244 n3_13880_11663 n3_13880_11674 2.200000e-02
R44245 n3_13880_11674 n3_13880_11696 4.400000e-02
R44246 n3_13880_11696 n3_13880_11721 5.000000e-02
R44247 n3_13880_11721 n3_13880_11770 9.800000e-02
R44248 n3_20630_13924 n3_20630_13971 9.400000e-02
R44249 n3_20630_13971 n3_20630_14020 9.800000e-02
R44250 n3_20630_14020 n3_20630_14039 3.800000e-02
R44251 n3_18380_13924 n3_18380_13971 9.400000e-02
R44252 n3_18380_13971 n3_18380_14020 9.800000e-02
R44253 n3_18380_14020 n3_18380_14039 3.800000e-02
R44254 n3_16130_13924 n3_16130_13971 9.400000e-02
R44255 n3_16130_13971 n3_16130_14020 9.800000e-02
R44256 n3_16130_14020 n3_16130_14039 3.800000e-02
R44257 n3_20630_16174 n3_20630_16199 5.000000e-02
R44258 n3_20630_16199 n3_20630_16221 4.400000e-02
R44259 n3_20630_16221 n3_20630_16232 2.200000e-02
R44260 n3_20630_16232 n3_20630_16270 7.600000e-02
R44261 n3_18380_16174 n3_18380_16199 5.000000e-02
R44262 n3_18380_16199 n3_18380_16221 4.400000e-02
R44263 n3_18380_16221 n3_18380_16232 2.200000e-02
R44264 n3_18380_16232 n3_18380_16270 7.600000e-02
R44265 n3_20630_18392 n3_20630_18424 6.400000e-02
R44266 n3_20630_18424 n3_20630_18471 9.400000e-02
R44267 n3_20630_18471 n3_20630_18520 9.800000e-02
R44268 n3_20630_18520 n3_20630_18527 1.400000e-02
R44269 n3_20630_20674 n3_20630_20687 2.600000e-02
R44270 n3_20630_20687 n3_20630_20721 6.800000e-02
R44271 n3_20630_20721 n3_20630_20735 2.800000e-02
R44272 n3_20630_20735 n3_20630_20768 6.600000e-02
R44273 n3_20630_20768 n3_20630_20770 4.000000e-03
R44274 n3_18380_20674 n3_18380_20687 2.600000e-02
R44275 n3_18380_20687 n3_18380_20721 6.800000e-02
R44276 n3_18380_20721 n3_18380_20735 2.800000e-02
R44277 n3_18380_20735 n3_18380_20768 6.600000e-02
R44278 n3_18380_20768 n3_18380_20770 4.000000e-03
R44279 n3_18380_18392 n3_18380_18424 6.400000e-02
R44280 n3_18380_18424 n3_18380_18471 9.400000e-02
R44281 n3_18380_18471 n3_18380_18520 9.800000e-02
R44282 n3_18380_18520 n3_18380_18527 1.400000e-02
R44283 n3_16130_20674 n3_16130_20687 2.600000e-02
R44284 n3_16130_20687 n3_16130_20721 6.800000e-02
R44285 n3_16130_20721 n3_16130_20735 2.800000e-02
R44286 n3_16130_20735 n3_16130_20768 6.600000e-02
R44287 n3_16130_20768 n3_16130_20770 4.000000e-03
R44288 n3_16130_18392 n3_16130_18424 6.400000e-02
R44289 n3_16130_18424 n3_16130_18471 9.400000e-02
R44290 n3_16130_18471 n3_16130_18520 9.800000e-02
R44291 n3_16130_18520 n3_16130_18527 1.400000e-02
R44292 n3_16130_16174 n3_16130_16199 5.000000e-02
R44293 n3_16130_16199 n3_16130_16221 4.400000e-02
R44294 n3_16130_16221 n3_16130_16232 2.200000e-02
R44295 n3_16130_16232 n3_16130_16270 7.600000e-02
R44296 n3_13880_20674 n3_13880_20687 2.600000e-02
R44297 n3_13880_20687 n3_13880_20721 6.800000e-02
R44298 n3_13880_20721 n3_13880_20735 2.800000e-02
R44299 n3_13880_20735 n3_13880_20768 6.600000e-02
R44300 n3_13880_20768 n3_13880_20770 4.000000e-03
R44301 n3_13880_18392 n3_13880_18424 6.400000e-02
R44302 n3_13880_18424 n3_13880_18471 9.400000e-02
R44303 n3_13880_18471 n3_13880_18520 9.800000e-02
R44304 n3_13880_18520 n3_13880_18527 1.400000e-02
R44305 n3_13880_16174 n3_13880_16199 5.000000e-02
R44306 n3_13880_16199 n3_13880_16221 4.400000e-02
R44307 n3_13880_16221 n3_13880_16232 2.200000e-02
R44308 n3_13880_16232 n3_13880_16270 7.600000e-02
R44309 n3_13880_13924 n3_13880_13971 9.400000e-02
R44310 n3_13880_13971 n3_13880_14020 9.800000e-02
R44311 n3_13880_14020 n3_13880_14039 3.800000e-02
R44312 n3_11630_20674 n3_11630_20687 2.600000e-02
R44313 n3_11630_20687 n3_11630_20721 6.800000e-02
R44314 n3_11630_20721 n3_11630_20735 2.800000e-02
R44315 n3_11630_20735 n3_11630_20768 6.600000e-02
R44316 n3_11630_20768 n3_11630_20770 4.000000e-03
R44317 n3_11630_18392 n3_11630_18424 6.400000e-02
R44318 n3_11630_18424 n3_11630_18471 9.400000e-02
R44319 n3_11630_18471 n3_11630_18520 9.800000e-02
R44320 n3_11630_18520 n3_11630_18527 1.400000e-02
R44321 n3_11630_18527 n3_11630_18548 4.200000e-02
R44322 n3_11630_16172 n3_11630_16174 4.000000e-03
R44323 n3_11630_16174 n3_11630_16199 5.000000e-02
R44324 n3_11630_16199 n3_11630_16221 4.400000e-02
R44325 n3_11630_16221 n3_11630_16232 2.200000e-02
R44326 n3_11630_16232 n3_11630_16270 7.600000e-02
R44327 n3_11630_13924 n3_11630_13971 9.400000e-02
R44328 n3_11630_13971 n3_11630_14012 8.200000e-02
R44329 n3_11630_14012 n3_11630_14020 1.600000e-02
R44330 n3_11630_14020 n3_11630_14039 3.800000e-02
R44331 n3_11630_11663 n3_11630_11674 2.200000e-02
R44332 n3_11630_11674 n3_11630_11696 4.400000e-02
R44333 n3_11630_11696 n3_11630_11721 5.000000e-02
R44334 n3_11630_11721 n3_11630_11770 9.800000e-02
rr1ba n3_380_7221 _X_n3_380_7221 2.500000e-01
va7 _X_n2_4880_10596 0 0
v21f _X_n3_13880_13971 0 1.8
rrda n2_20630_6096 _X_n2_20630_6096 2.500000e-01
rr1bc n3_2630_7221 _X_n3_2630_7221 2.500000e-01
va9 _X_n2_6005_10596 0 0
rrdc n2_19505_6096 _X_n2_19505_6096 2.500000e-01
vb1 _X_n2_12755_471 0 0
rr1be n3_4880_7221 _X_n3_4880_7221 2.500000e-01
rrde n2_18380_6096 _X_n2_18380_6096 2.500000e-01
rr10 n2_19505_15096 _X_n2_19505_15096 2.500000e-01
vb3 _X_n2_12755_1596 0 0
rr12 n2_18380_15096 _X_n2_18380_15096 2.500000e-01
vb5 _X_n2_12755_2721 0 0
rr1ca n3_11630_4971 _X_n3_11630_4971 2.500000e-01
rr14 n2_17255_15096 _X_n2_17255_15096 2.500000e-01
vb7 _X_n2_12755_3846 0 0
.op
.end
